`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Q2RY0NzAYOX4aZtvuSBdQ57+Q5x40zgszLcnDO2AyDzN54BMlgN1mW+QzrRlO2z6t7eyNW1ayvrG
M/GfPsY+oA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
n965+Tb4giNN9ZtzdOl0Pw3cJcxAQnzjWP8Rx6wewpaC7Z6Ir4YJHxlSxyNER6xdPaHzdrReuiOv
HYxv7BdKOFBRj3+EfVJttlKH83/T8TXZKeSmvTouMMMWt34YYWlZJKS2GeviMjBdCkgNIOYq/riI
G7UURGziy+q0DfGafx4=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Cq61/r+PAF2C6tVUk7PpHQBXV0AIRpC9KUKn7BK2R93EcSb0vemDXNPBFWvftLX2+x3SET6P/iSP
stpQNkGaZcJ7afs08lY/C3xeqhAvyhflVXp+CKvUd8Dgv8YsxjHENEJNLyuG7EwEyNe6DmnSBfpA
X7XA18kXEhQrSjlQH50lCSMb+M6pszukDnc7jbyWyVG8W+DAMiXha2X8SC3qPPJ4oRqr0jgoqqdR
a+T/YTBv3t2Ifp3exv5p2NrKMlNXsk13JT7gw0AcRJzt8lN46BjMg0qLGcebcOAaBVzvXzBVdPkv
5UtCMCwoxwkuQNZGo+/FATLnTAwakETfh+eIog==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EDwWkLu1lZe7pxkx2nwH8GlbDeZfuEh9tvcGWyFtkM4B0SHZPza6zitc8Iijhp2xTCHgCKYwfplZ
Dyfi8RlC5gH6hBOgLN1BK2NGx0wyonqDWRpIalFuOzI3LbN287dyIXJ3ysR8J0oJMAkLIhjwkAO8
CbzRICgEdkwKMknJYrQ=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
1XSjEz1FXGL/HrLLAzbKduE3TnulJ4SF7uls7W6Sc1o6DVsClLu9J66ijCmApppBQrNV+LVp+Ljl
nhh8Ah8heZfx+inUTnK0hkmylFXGF8UGZ1XqfOZrfDUZe4C26rBKzooVo9Z+U7AqtBtvOO+J76Nh
b4PbT59WyL7cskTPtm5xq5qC6WkvnDlJFXJ70lq8Dxi1bdsoXhJq+9fmXSflaGoBQw4/1FbS2FpO
VaiGXiSRYyGsEM8e/6x2kSacP2o2Pacad2Zm8Os8aKFO/pycqINbtekN7YFH+W60gBZPW1KE8Fyu
SZl+P4odBkxcGj4bw34AHF8Le8J6bqCV3Kd01w==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
X4xjaYk4P/LGUHSiYGGkWvAZu5izn/cOCgBWx+JpfwXd9id71urcDHmcFSplX3g4eCV9MRO51QVs
cD/U/UgZLGm2Iz+ETgBqPXWqiKMV4hbsL+6Ork5NtEzNMt3LOGT6yRvM/tNqllpa27fwBUrRuEEy
DcgOgKcnOs3kjRYkMU/oyWWJarw/ceSuGfnv+T+fUawb85RVjV+/PahS8J8RtxwlNvBm5cHiTI7+
4wprMIUqATy/0CSl3RSZnv31POKY3rsSMAAzccnOfOR8ylj1lgvKqQ+ISSL1tgxluH3pLaxe8wmq
ojni1/3VXVg+ZtyAaC+i4b8Zmb3TvXHL9VcM0A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22080)
`protect data_block
JoBOllaM6EDZYEmxgR7825YeNIzA6qHUCWl97EpFvMZzJQq3kdczAAcNijKblTENsSX861tiYcvP
Nh5o6DnzB+/LpByTDbhr9EbvPJ2jpUfngTd16IsOoHZK2rgSAEab9C4I6Gd9RQESiKfF9mM6rRzh
2IgDb7wKz5VjSQXgorgCStwks05CGxWj7v/qlkjiLe4bvgnNXdbs4Czazt5jDCZiuc+mmZNyojjV
lr/KCJc6K5e+cuyIcEaOcBu3YVlOOGGmY7Miy52lN2W1tquYJvFH+jmcnMfdsjyYPTkL7lOHC+sO
IpYNXpg5fKyFTrc9WcZ6ygjPoQXycZtCbEL6j/bmRP0hnpQiPpxlHxNyQzWnTaBmb4Bpb2PQLBr4
xNkMlB4st8fE5tVvnfGvIlR5qB8ytC7zLyNSkGg9H5s9ckFQese2r4N3rH+TKOBW0UNmKtpL8+iB
Oa9M1MHUE6RmSpKshk7pVcTmXxLlmpCLX1OLiwD+wzRFEyMCMk5eACBWJ8WhAWgWYSgPrKpYwCpb
vrRvGtWNSoIdtX8PyJhqLuQ5aTz/WuwT+3B16WDHMo974PQ0E/2QdjCq14FRyLPOv0KAojA87dCy
I7dOxdVMh168VZEyPqNIFk2hJCrKncxwzI4ZvykpjZkNqTS5PIPZLSaVVcGwvTbAEHOvejnDfvb7
nJY2pEwYBf5bbDhgFq82U35TQa5Te/eVERbbmDkL40VadlCvg8uj0jHV6WR/1DWGLm1gE+iLvf8G
B11iqu9I03AHPRdfsC6lX52zwY+ow/QortH5J3aNu/ipXpZfg8VvCFNToORAhtCdZkaEyOSw5K/+
Zmwugb4NooL+WbqlRQt/g5TUM7ojdQbHzleW5d2VfIP/GXUMNXg2qk6E48j24vqxoDhq+AGQHfqO
ivf/Ik9dj9/9f8rW1TR7A1lieDd758z1/qieaTai/Y1Ayj+SaV+Ei44tBiWLekCjVFGD4qyB4tjO
6meABMvPxGgxZlb1Bryxe8OORKrTLYSXgR6Nc443kmNdUoMd8sUZ9Y+gHLJuBlr0DGhSipWUGXNP
Yfbqpyapd6mTkYzygVdYmIb6OrzRAXgPrmTUpfH+oCsvd+p62E5W5pusCCTh/oYOh6i4VX/lPSZX
Ymb8+92ysNHGfzAksN3Dwbp9DlPvXu9Zj9uJvPMH3E0wMiI9+ipORqDaBzN8V7PZObV5YVN0xQVh
MK5sVCFGgl1nn9DVcFwoZgiKbDoRl0at4UpF9Xvc0ZjwFDYoQWKMnUN78gvj7iBEMGQ7Umg0mLJ9
OhSEH6QhiQJBx21yK9hMvt0GDvfKMNNdpJNVD5hO8jYwwUmrtzS3GYtKpD5kIUvZ3SBW0Ao3TNQ0
aEnffvRvOhXLmjUZAbk6nk3Z5HqMStHMtcnGh7OJcZgzugQmvDB90ZMbktOyvjpOBCYH0+9JhOWC
9ZrkaD51T+qH6oESZo5b0di0diWNePsGX5xk1K3WzVZbmbKmpsJwxmYMuKuwPSLZBukij0UkA6zl
PB4um9Wb11x6uWOgA4FjgyMM+IOPbVirO5DlNEtLspjPt1dUcAf+f+Q0H9kvcr7VU1wUVlk5jg+D
yHMXAWGjsXIn0Dibf0M/pRtkVETcn1VOT84Hl0DhAg+V9lTX6wk8W5yU8EJRzsDbG10PsHn2oIk1
Jqp3wEpdorPriEhbomstl9NZVIJtbOgmukg5qtmY5SsSXYGEX4vh6CHRNrk3iq2Dc1rmCVWn8l75
7xh0Dhc5FLnPmuTl7KlqeWBn/VfNGPRYb3hRCOICLLO/qRFEFrdp5q/EEZkF+aweQSAJAcVz2Q2f
VNInT+ZrS+Cbqdh0PC5ajYWYJSfY468As2v9sKtt8ae+/cLvTd/DyXrKWEPJKkNfKk0MV1BZceIe
vMIdZP/Akol7vDur82GB2JDltHyGi5XTtECwEi+FAU6qN9szHh5fvsZKKhAANaEgyJIJeYT2S0sl
PKKAZiykG48TEIoVoEBVj9GCHVOnBqtyK8oNeWJSt8JD5VwXDvjgum1a2eF2exvXaF75bLhpqaSP
cB79nU6wrE0x5ZOVMef9ZNhlrK355DGF4298VxKlilWiSRANH2UcHpu4nUzjUcHM2swCQcbIFWuo
8AcpuawH712grPj8BCdj3HYSoZskcnh36xw71hBVNgTZg2Rs+fykevfqffKgtkKcSFHkfYFGhi4S
K+GsrqfkCNZYv1kCAncVL4SX50JLLurUrw+PpubhDwtV3txo5dz3ADLXoc1tbXwPizRmSj8fSBEs
k+GRmuW+7LojJIPhAlC/W2awOtrCH6VJQ+1NVcmvmp1OB4SReNfV5g2UDzuamnLGb/IMbBLA72Gy
JHx3taQQzSVHJKD8U9Xi/1JD6KXJGwolAh6/9/BaPF6s9tsDjIx9bOFuHY6bTMmVN4W0Qp2ZFbU7
UoQkszEq4om4x12GCX1YDzExUI7uVM22HENF23henHE0aediSIYNWvY4r0ZwcNrzPAFYXUpv7/sQ
RwO4tmQjyZ0lk0BgPMV+8gaTU47+N1dmCDgEMT+tYp986fRmNj4Br7S5mVdGv1OqOOEDZk8q5aSc
3r8ktkAySthhOa//i52wPme0X2bTYtNqvIZYjL2lNH0ipuZasydqJ6ZZUciJexV43tbQMGDBxgdt
qvkIdyZnNk37u60qf8L7A2H8S15rm9M86ncUONT4dg5RWmEhQlcQmgK0mGyETnbEj4S/nIVcXk6C
kIF+/ltF14JILQE+yIzWdJssMNfL8P8dQGza5wsK8EicQ8Nr6NrZqgJhGoRV8Er49pmQaqZSaeyD
TSCOQdAM3c6GD6JUBvXWjRXN/eMU3O+2ZREE720V8LwU5bTWc5lU8juxIkXn70KwJGOmJLLoRMgm
ILyeYd1Pm2O+66Jn4NXQoIt8/L56crh/r0M+l7RageocfC4TWXkyUoFGB5OZkWzH4fhUTBeTsFmS
vYtNTj2dGtfb88gWNt/oGLHpiHj83iw0TA2UH7xtRyV1tnuUWdttfDYxKpiFgoPqQITkBTPJgmz5
lwtphVg6N9/v74R9nZzAK7DjY64gIRHheBJXyLNlmc//NnXm35YhOl9zr51+st8cZmuBAx6cTxqj
Sa3lRFXi/RgewjvoihEkvGMpF3vPdZvoU7Ee9WUwhvFMA2SvRq7GefY/W649DjL1rmPt9zEwcgks
+GqRDaY9xE2EO8UZYtu13kS68MltkHRlV0x508gsTm7ZBvmDyxEKlw6yQ+cBMDRqoOETNd1LiODa
a26oMe7JgmurqmABNS3w9UrCvoKPXams+3wVnDRxw3NAj2BpKqPWh8gR5QHJ1pbriiyqByxhXmgT
4fPTuFsVH/UNjz+Aa/70pjCkx/EGCRfWZEt4PaDWspEVWnAIEsU66LgyfIJ7dDvO/0bf6Es8R2pi
Y8dzEZSEAK6kMOuAUdZjdTzM44Gm8FGYpMZ7BvsgBoiFoK19NP7gpy6Yt2UKZagrtWvQK+e9ijHQ
MBk2ifpAHk83Y5nUgBDws3bHcW/bK6fmCoHmGJrc+FtyI2yIDAnJ0YLA+6nyU6tQOAL4RjHhv2DS
2DNoXPWjVghXT3cQHXIcYNiOD9h9YHQHNO6G3Rdi9U3//qf3A4LCaJT5fBNJbXARreybh8MbTI6m
87JjOexHEtoh8lq5Io40tNN3cvtaE6dJMebIHrqtnrWZmCg+/qNA2CXXaS9VRu/7kU+UHZQQbLz8
61WZ1lPNFgEyujFNd4LKWJG7OMMvB7Hai3Jw557YwU6+KJHEHWrFcHHSb71nJYazm5gslTS6C30V
o3eAbe3F33QlRBWoQkmOQm57A/WPBwryDUXJurTSjwhm6IdW8SfF3W3tq3wGXr6E9d8wiQ4hYbhI
KQwHK88ZoIVkljp/fv8lNWWbAvdsr5xxSJ2htvKLTkFyAfGx4YV+kEndb93r9WkImDMBZmMdnK//
iutZIiO7an0pQ5poIgC598GbwvW1dhEVrjEkdS916KHbm5qY3EryxpKLicKNdNYFvmAMy3yDmoPZ
1xYl8gPewVq4sCXv2Zyp5upnc+7nPlVB4RqjmD+JUB4615y+sZPKZ0nnyXpEPR6goO8YIix6Z2LW
PmkK31eokO09FQL081qb+TY2Xens5TjG738YEg3WNzytBVBdlnsNvWrFjd8xNZ5GHF8eDgR4K/zB
SNrO1r2AOsW5al+++DIKp4UwCTnssh/8SY95lqfzfDIqIGmY6fv6G5NFKsseCRTmwaQiujz4l9cX
2pfzhG+MLfhkzprqu9QgUV8nh5K55YZVCoVDSv05e43cEkdsAaVcckejk/REMya2VDKGcU+mVZb2
GsGNrxRxTDcYBP5nr9T4364xYA2Rzo6wMpJJ886NkX5PysQKv+YDq+gzNW9a0FB2svCFkqsotV+n
XaEZmARgtWoYYD5yim98z4RLxwS91Su3Y177lclDTI+OUdqeplK13wzHpxXucP3M5OherRbHKs7d
4nX/KFO/XJ/exBbzk64tfFML2u0lykz1+fBGCeFZv93E8CR0XlGRWi3/cIHBkudkUpzH0rvGxieD
sp88qJBWDiKMJXP7SyDTc2I+bgXAVKWIg9q0WL2Jbo7QhhdGBnABz7JCNdOzaO1N4+la1v/PAxiW
c7rbWGA34AItgz2nGmbTMb833QV3pOgfLWImwiH+9ajWrJXpfBk3zYALFowoSlBvvXqN0bnhuNOT
BPxmCFfYCUTnCjTQCjxKmq5E5Cfc+Sy2QRt/jXyr7rSkkNuD/tpPvYbUunX7d5taIo8zP2gNO0/Y
Y72q/HDGFvdCqMU2A35OQiIQPnGJgPaJ+byqR+MuZcWqR3pGfilVNHWfOnfPx6t3cTOmj91ts9bS
K3o9P4pCJbJQe+A1I4OqVG7iWroguruEZH7Egfw68kcGVpIR/ZT5ci54gJkfZpCIqmV8QTnLaVlV
6tGIIinWopMSG6bJqTe9OxS9898XF8iDOxtl+aOicRCLZe/PPzjIC0avN13uHrT0Rj7+DySRG1Jl
TNqayl+I91b/85JpcrXhQ4TqC2kMxOegZOGU6qV3B/tVWWPf1mqQ1nZ7H6BRfvHNJLeKFHTlJbwj
lKvUBlufmZFb1a0iDQy8uuAIDDEWL6HV+L9xxeVvANDqF9xbVS8zTpnVxLX+V8o1llHQcXYbGdc8
rvNU64HuNDXSyCzJli1u7vKyvG9r5k4ec9DsBMd7KUJ3toj4jKmbeE5fhWT0NAmf41AWP4iCpKu1
mv21RHMUCeho/6N0MEhWgFmfOi78z2D/28IaCLe+O48lnNjkdAHLnzUHu2HMWprzRnPxc94LHlyZ
syFh28en1pA2QnG5swg4MEZlyVsNin0HFTmJ6qBjP+MHHFyRJfBxZ2zIUe9rpsm1tGnekUg7Epud
ecP4FlxkWuHznIwxi1TTyG6GIrQD5k6Lkjwty7+lRD+h8RbLTt8KYC+dlf9ebHHarjZPQYUlrZR9
vyBrwRhksC1qUs+kYOSCQZ1F1hIIsUttLHp/KnjdSXaH3Bvx2yg9bzTfPdkl89vPPoWN4XLABARB
RolkxaWV2g4NJmtzgjz0mUuXWQcXlJukq9ImVWIE2BV4/3/Jr90q3nIvuCQUm11YyctowYGbR9rQ
IN3Iy36hAMPG9sLHvClv0KdVe2JxVbXyUe3YFeDWRNF3RgfChNhaD+MR5JnLMQm1/XoJuN6dOPUk
JwAvsWKdODGcqIXsb9SLoYO4t41cuimBo41855vsZSO7ysnQYxwUgIe2N5ZX1fPJjRVsfvF32HsP
9jDet/cvemzyqBXyYq6T05x4yfEY4zKlOBHNP/0aqcMf3dVq6Rty21LHpj5O+J07ZCZhqj9xOIVb
iJs23QDV6gU7QI7Hf2l+JJQP9+AyCwL5peqaKBUBst3eRvZZ/8dC3Lw8CsCoA0hAyKrYQzAezfUB
6TsEzoYyNik3MM9tU0az72btHHSIgvnWamXPiF9+ncW6ovuDfDpHHA5GTJJGHuWo3oQalKBeG13a
JIERepEAJbXGcSypmf9uHF3nmr2UZawIL0ksgLOj5RczCcxGXcH21thMa4Wdl+uDotFyyxXpFzNy
/6o1rHnuGDhh9OHF4LcId/DJK2LURbmQGoYmDYqYi9VIRSmMUitX7fPBTzGekSoSSw0qm1eJFtj3
Rir3R352/P4EAU/yBr40jd++s8hHbTsS8LjTAHP5EAERGjMyxAGhJr4f0XIAVDvGsy94aFWA+vxw
i3mTDu5qaHUbhhwbnbDlxypd10HpSVTyeRUNx+nIkMPDrWgC9DXXjEohF2c7U/X4oVU2N248LenS
FCR/iSz449+ld39cGYOBYzde+hODclLJW4eQ0LIra8TBzZtvCMTUQvfiGcCT6lmT3yHLG4UI7KgE
BNaV0v41pmfi04bF4pcf7+7/XNRiE/ZGeoMsFD/LR6BDJ1YJLQPiEbGrei6lNCR3gTtqbYS6BV/T
5R+fuVT/gIzU0/k//Rp3ChJE4+J87AfMiJfk2NgR25LsE/75KjTQd8HErlzERQAxcbVu2T0KGrM5
wroAFJfywJpWGQTZfenbcVwt7UaZEqiEVMwZXb93ayUw+vOO3AeU7Z5LIzVOti0/SAdU2OjfcOqf
3bBk5uXcnR80jwuASOUtOTtyUFMuwf5liT9BY8mhe+OjLRkDW7/wR4nDOiWuykXBVsHNXpeb4UQf
A+oNzkfTx4hB3W3JLa5cbIpZnC8Gu1aQrhyEupg/3J0T2mEX5YArmgrO8335pOEj+m4tsCog41YF
c26e3FUogu3LgdcxW9VF1Ng+bGpP0PAQGexcyatCfCgqK+N0h0v7ZXSfKWyxdpjlxWI0jIv68vVE
6NYZWWm9RyR3qZe0ZJC8xTQ5xrSUDtVvdWnKZ7a3xdK2Oubhx/bmfD+joIXv9IToE/Dg1SP8nEAw
opmGiHoe29fduEGuyDYX94AqTpQCVhKSRSpkxeNSMZlFTfvO0PaoZG92AEkUxRJFOeT0OXVHb5+R
85C2uFobUmO7Viu0qPta/BzLP4siT8bng/IpRzDRjQ1N+saDo/e8i/Z3gfIqaOFIY88pqoXCNuWh
tHhJ6DM/4+W7ONRZd5iym1eBjVrCMFktexQ9mn5YJVVvnK+39DiAkncG4VjvVQl0WqrRZCRL9yUd
mYqXzt4h0aWTQul64g+3EvJMw/u0lRNFrFSPXEd9J0UAHtdTfWZhJBDkUfeByAo/8qs8zBFSSKRl
PGJcLMmLgStK8OrXdqeAKK+yPZ2bGQSMVIRRNoY0rZzKNuDWyy+UOwy2aR1RvLMOGPu4j5+9VfgZ
UfIXWe1foyqkkvU3Fqttp6kE4g/l+AiQVjee1Ifo0YgHjRROmb7DF/9HQip8IZIRbQgVahneByfV
FKIWPYw/gi/RkRAaO11RCmG2E7btu+dzAhVot27dlAEsylBdXaxzDKiGHS0fmL4iS8jTMyOpWTaY
SpLHWGJlK/cjZrioU+zFooDgy/GI+rGsDzbdlwX1DBWtSE75k9PEVqO7zXY1xau4+tfB1TP6A7cl
2du/bU+1h/N+U4ekfC+EZbTSPw9h+zRiYUhYf0KxPcn1L8LhSh1HgFawrxmalGSH9XhKErUIdm4h
30wQbB71JAGVeF2KeKLm+WmPQw3rwfM7a+K7liRbceb22WBIQWbBN7tCvn5Nx9vjxnqhf5Ib5Kua
96dOs0ubHAMIlAinaULSYFy36pEOYLh1EMnEgbEsAYBGBYa4pJPn7E9kiiE80U4SaoTQG110aUZJ
9XWS7IHA+JimXWqw8nfqoqzbvPECofqwtSF3c636QdOFKmmIE6xd82VbI2hfZpqEnO5wSfqo0FNN
2lclamtURDL0bXP01CRr/AIpye51fME7Wc9RjhSkl8etmRIBFig21GtTL/irXQVyuM4qbCi8c/yM
oyrTnujasEoUlgrS6C4i+UEKoVqbUWCZ/eM3o9AFPulA/z7lAcR/kVOhr0i+6bMVeWIIv+CuBDEL
4aF2RaRSB3pWHdSUsq4DfoQKuZ/+JROZzhHo/DjUYbv9O6pvtyECg/Xf/TpnEMiOUtH3huBIhwNJ
Jpef0nNflXZ3uKKTnf0IllTuRC9B1ksy13u2dViUxMgZwc2IcbRD0m8/ljzQIIdmK0Z0hPONpJEH
itqnDWFgQ2/7mcZ21B9mZ8G4RSpHl4Nax4NpFW8RyQPYZ7cYJsXsH7Udd7KoG/LzmM28pTKdJJUF
NCJx/foAUC0wg34RRGpn82cH59EJAzjfLkdn1EaPmPPyOqcw5LW++DnEPCVmJRtczQd/Rd7LjEkO
TkTtxU1mm7g0/fGe9GguIv+ifkNnZzGhDsqurH0UthSYfkSE9IxbM/0Vt739qG0R/E0oLvn7LY0g
zAeGo5b+MFUoeeYmi2fw9GdH9rdeK4Zt+/p5sxJsd+1JP6O7yyNeALQ5RdUdg57oahacpW4Lp4rC
cRma1GqnIkfHwmmScQ8wgqghly4NXgobE7gzbcMBGsiZ6XjJvZWK7O5CYmlIWh/e75Z7VK5ChkHU
w9RFjcu9IwaI+8g3F4NIaMdz/P47yLffmOxFQgEDg7GhOCjzEVGqnAkLpfRSLbEl9BMZouSf2fGF
dhW5e1/QakGmfwtaHN5tjEmpdkKR/dja/zxlSHpgr+Z+hQaCx/Lt6RBEbNp5dj7NBwppCdt6on1i
/pJOepsmoxHLERl2gFDKsmfNLsbCPlJUm+q/E4yi1O7Antc9orxw01qGTXfKrG+WvA1eqsH+4nLe
W5u1uanZ9WB08QhxALm4BL4RQZqQbQt6BUFXqpBuRBHKgBTqurWVeIYhFSJAN4oK9SakldEB3R9y
b+4TVkdQRhHRutW0i9hpkcpXJpJm209CMAda0juj9N8urwHCM3cqQawncvk2HJygmtMkglz4BOz5
q4iV4PaiqMyjrgVmqItlPhMJBgdFULsPNB/k6BSj2mEAung+GYD9VvlvTt3Gq7bErnogZYly0W0U
MvsYaQzTHeDq6kM0IN2G6/1crP7q0LNpLpJgU1lnYzNDdaXljW4Hi0P32Q9/d51qcp65HQ1LwAud
bfm4kkIzWRLKOwdVeAurOlXGPA3+Q7xOnh8WHtmDoGc7gKupFfNI1lHkWE2cKOdPgCJKUaX5zXTN
d9F8dKhpYwueWx50jppb9c/QnhNIjsh2oHaYAXCeplY1iMEFzmca+2V1V7MCMKE7OsSITHyeHwUG
hgioSnRjGAefflZtHsav667blsA21HlSWFM7fTFs+qebb+k1tfMxr1dj6qmiFruONVXzF8mCaoID
bdqMX78QwP5yUCgXdgi7dh5xR2p1Bx8ND1wTp5Iu5aG18NB1rX/WvGGX/b0iBxGZcx/4cMwuqtJ0
7C0MI3hgU9hEaEjpi4JRDo0g6CBdkPpVSmvsn5dEbaoR4Z6nh/i/bSHlPbeGS/wSo1krIll2l8wY
xGi3m9GDrZtp/nLR04Qbu32fTlMDUDCWr0AeX/WOHTLnP95b1zdjepyQa1JBt+hqbsQ/ZT41qi2C
M+J7Ip5xkEeZ1C5LCgiTHM5PbNxF9Rz8C2sm++mYtsUo2xQSDht59y/bwJILHXJtwLZRwYdpjdCM
AoHhDkNLn0RP5So7KZsXy/AbCbZigHfA8gkQZEQwCo+9Ba5n9XBzSdW2gHoOQTeZrj2kadq7hLL4
sOY8nTY60aeK75DEhGD3a9rwN0oMpQZyeM2frNq+9EvyRdMMioMs5HJk7+8lTxschIy/4FlsUEpU
j4fcwm4GJzaiwGr033sdjxs76ar/3JLWn7vaESI/AssHpnWps//qGRRYznwTnDsbb09283goOsTd
wtF+830FfBusk9EbVmpvqmrh6tyoRK6RGobtGMs+FL/sd0/37Mma7j61YBBtRuoVv4j2cQyEZqRR
EoJszfh80rMtMdDAIeT9uWqWds1cqlxWtjFPG5eOvR08n5DIvVWjKCpGmFoqaSLUkfQc4IsTpN7q
oCncKF8S9W2pjN0DO7hKxCgnQl3qEfIkCYDaMdfOxoqNmy9p/EmnY56GE0HT0/LTmXaPvTq0mlGO
0c6ntY3LWT1qKrgWnSeRfcwNdWU9uUiqFqtQmDg6XCxky+DBoh43ZTQVTcXx+6dccixKGeIdeBW+
08x8P+BsJUYnjhzNT1f23GWp+8g6XiX7HhQQLgCGNMY19WAGcgMzC1CgW+156qGi8yAKaSpMMrMC
pqwYxaF3qnxo6asvv6IFI/Xge++JIBjWCjQ+gDQxRyK9A2pIjMJmgdzG+yuuhHs6WkH+t1V07T9o
sdgLpQb5FW+VZTEKscOw6icHJL9dCJl8TtzwQolAYDWHaDWszL2EJX9VO3o2q+z8Qzsy1/kJRfWU
asHOykK/gKiv3FBXuEWsBZ3aJ4pn3QG0bR3Fhzc+p8xZk3U2Zzea7CrTA4qqgFVo3Gt2B97d0LjB
8gy2JbttFFIarj9SMWdRI47aBBy+yBaLy2hc01y/BtJ3g0a23m/YHhRbxR0QTLhwE60GjUWkFt7W
kksNgFR7NBe3s3lnyjMWGQzkLUEKnKpcq1KYI+d2bD2+aTv6Am06tR8F7HmK9uLxW/LFjVUQMeJK
CUvGDPznnUL5aTPYGS7wfFLy4wEY3gGq+Amxxnul/zYRnCGiBGg+plyEqrkD5/Vaw8ccPbXDANN9
B0FoK5KdJq4H/QnAdBxooAqt4U/vBlQMeFlwczNGAibB6wSL0W9ynjWZ5L9q/KPiVboqPPcigDtH
aaIVcG1xi2kd38e4wScPK5L8GvytJzXYqjeAR7OhQv0wEF5oJ1ML160ssIV9g67ckDA6+AMwoF6F
NILQVPFGWNntGqmr+NCfGEQXSnzwZe07S3rpuh0b6kLo0GwSbfLdqgxq7BH1PktGi7L9eEy8UvNw
ZZZQBdElmrZJxtjdKD2OHvqgN8x7K5nD+/sveuijxB6ht80A86sjr9rDgwcXPHZH0OCPeCKJcf0y
UVNOZU+WVs1nF/XsXPaSOzKkDKhYJsbE50gE4jnfTPMeO+fuyKWQhtS1O3HDdIBgRn/+bLtdHiIU
XjrJlQnlbHlGo+EbCXEYqa9I25snNXp+e+dXEcHwvUQGmUCF6EUPL0WenRwNnLE6w8vBvmzLUloy
XJpkSoTZQ5CVX08FAr3qbbmr+QDEKEuqTNf8bxCXmFNVl+3tJ8+HvVkZ2Akgi1QkqboEaMGhjKun
wgF+zsfzQpWcb2wu5LE9BgpnwRSaLq+mKi5vxSvzuT6z/E5QqkugJkDRsxZsXvuWK61jtfUvUmRZ
9xVKIuDQ2B0n8Gi5N32hbTHZkq9+xhbX/vrQkzKqAxmS2PxBKDEtrSoj0iFTYRZ29l/huNJyqcHD
JGcCSq2CkxQOKSp3p8FfETpTze3OV2Sb22Blan6Y5GntRikNNONd6VKWUlwZAmdmIDdBl6hJP6Ol
Z5iN21oUQXZ8cUTH3b0IPfBIEDQOxuRPCBNNtz87li95+KPX47n/7NF56ef10x7s0Qzh6B4gthfh
t03W/URmS9r9nD7iFYbLgU+SIASD3+XP2lnLsTYxm37pbAZTMUqtqVJWHQ50RSwzS6aXpqoilUL8
nlZRlYFAoC2HhTNOjIRCtJAyGeQ0mu2Q/77oy2jAHeqvyFMd6WTkXIANHRtC91cb1r5FMEvRS7LX
+35AoCg+4IAy8cGqtz9DwhcQ4Y4OiyCi3sdn9wxi+tqisAOe7Tga93Nh1KlWlpQqVlRk+4QHlXgf
jMHOKARgg31sazv2PL+/J9Uxxjp/bUXpgpcGCEXaYa3m+xAHlxM9Xx6Rfdl/imRIJ4XKt0JO+fAF
by9vE2gapMTdAL/6ZN1FWcQuGmX3hlMT7zb3KAzwOZbKFWT1rx15HDCms/op7EmimgZrchAyM8NS
Yxtk/z9WmDQtSTRChaRV45RdA0S5dOFmR5r1ZztbkSfSztHx5KerEKkgRlxd4V1ONuVTLDjJjrwQ
TQFmN9FhmCWDagoIIIlNkiVM2ZqnWcve8tutoswO2+DJSqTPM4Im3Q9r/VKu6IxR0vhja/stVx90
BZ7en8yvhNAqf8lyrCwZdh24wGzDCJZDUk+eynBqlq7jeHB8h/XJC2s6ofdDQkjYg6tyZVEQ7/bz
Nzai/+97HdSpr+s70EwRayqQ2N0ebIJqfgiY7J+ePuGPyOu/vc0sYROhzb1z9xpDIZZJyM+XSNUs
YZEOEAk7Gq7W1Rxigwk/zghks/DP+GAw79hFuZgXuXc0mluqOt4Pg8qtjqwcxztJ3PB1kR0THnDj
o/YuUDxGdTFDuh70gnZ/2/heb9GAbx5zkXRDbQepvrzaSW1kc/IWt0Z8MfYufVUmR01KjXvqY++Q
rfiRbyZs7HVxxrcgUIMJhrJSvCohqcitHQ+IiQNX/8RlDHRUd0Tq9NDaUHbV7GpPOs0ERxt4eMYl
UE0Vl1Ko4z1CtEzt1BV2eUibvzQIC0qK834YhEyTGXploHv/C89peLnwwUOEzDYLYvSK9n3kHYKk
nE5Er62WWVrRKvkeHKNRq47vSSZIkcMIFGDeT5IKm6r0k3U4CnuIk7ynCEtA+81c9nrSPyucuPPo
LIR0P1Of5ruKZX9Nhq1X3GRZCAEp5kt+aqvCl90fs5aMxgShvw2Yl8oG999olPjZ6/szGaNHC4l5
FkbbMMz0pJnz+Dg9bYYd9bjAdBoEN04uI8e1NW7vB9Bpx8agg53iIXQSy+GBDUtVi9EsUKVukxPD
eWx+6aedtPm3vzx/ffowRXrk3e+S91OWUKN/XR3xPJ7o+qrrHQ2qPIRuy2xqtPhZbspk7DMbEzAk
tCZE0QViueBBf6iFwsPF60jqUhZ6wtyHhwmbye55B8gJU8BeYDH0RIGXuB3L9W+5+8hl2LSWbgRg
BCSpdyKHaox07HuUTO9vV2TqexElw1BJbt97HksnwGTePouWtOhAsotB0vjYRg7ugCubgj4+LugH
Z5zINYmwsndsK7X6rdnD48+pcGZDcSVEqjwAWD20nodnPg4nPdlpDVLttlJuG9n9WwdN2PngOEiM
jIHAO98juneVo2aUdTaeKoDpCfVNfqsKa9sHLcvR1nstAdlVscjG281P2QSjRiRPIIccamScD88F
BZr3ZyD/8d6Pk5ARvovqLXKZtsSvsA9Ij40HHD3kbQuJEu38F56MsXy7NzQKcVRxofPm6oF5OQ/N
S/CfOuADzDjAF1Hs2VRi3YJAZ82w3O0+mK+P48UczCw0r773WHZPurjCNgEGMH7XAWvLcIPEzT7Y
M84CdmtHXyX3tE8u6NIJgnL+grZifvsQlvDh8/8fqyz3YkV1tjjeOp0UmtjfRFTlyRMg7n5RgU9F
jKgUmLQxsj7NFO/q/WKTAITetYsG5fKpRgZorRrV8ZXebaz9c7tSArc1qeyzCf61bxtP7HsGJsaK
lTP/HQ9kI0C6xuy3yxTNucdIDRohzNrusrYdsm22a7B2+OY3GfhYpQO4S5daxWv1G5stjZIl4AN5
NFvYpDHbyV/eg7akTWDQQHxt+mjuHrb8/+R2MgwXKOEsopzZYzqA9zBkSVaCoxarMrfk7bWb1YTu
iksf4JFVmL0/UOjPmwVbJcoXEXa+lB9TbWJHGaTeQpUEunbCDcV32dqF74MCmVVvWpk17vv2w4LE
njGQXertQDygZYnziIIcx66J9lqiAy9MiHt4YB2M6SY5p/Ev4x1n+17eAFTWZlXCLNMPf7g1bwVW
xclnJnjrie1pyKS2p0SzUKx8i9nyCt5mioHG4pL4KNTs07iCYxvL5Fd0dgKaGn7TIVLY2ZLqE1u8
QzrxMd5lIP0ZY2ronBaHh7bOVxJvv0J8Vu1Txw3w644PlLC8u34800TVBWk7oFluOsjHzVYXoV1v
ZJCnHFcVXFUzKCxGOCrZtNmFFjexDOBuoNLozu1rWSdGyZ45XHJ32Kth1maiJgPLbskaTid23Slg
AWsStmg4Yspdd4MDOz0nkHl02BvKdaJzLfTC58eggpMKQmA78ePtcBy4fTV8GIY4LZKGy/WQnZXP
FHeC8AkNgSvCn1zZ6AHP91KducNGk+D/F939a5ehwOS4h9ewXTa8Kqh3b7wQCm10hgvXpsOH3PWZ
A0oXg+vpf7XtKR9lctLtS/XMeHcYlRvMzmrCygdSb7NavXJAn5kLlH+fn4+2zoJyaRwJBoyL0Xqo
vM5pS/RxfI4hkPY6AFbtec4wUm9i1swxMMFNdQIg+iHwLMbMmabw/p648Ekd6L2tH6kO867RiuUW
nxVZEEGoveYvx32Mowbbg39rMjXn1XF7+7NYv89yXfDT8DD4xHqF5wVJkp/C0LyMklEP/WhHYX8j
kFTs0Ds/chNvH7Jy5zVdnGcJPXXG8IQkYBbJ5bQVQFzvEhXgjgVASkf9/cbOC3Ui0LQBwHVYpAAb
20xVcJeplzXZtvtfIF0MRiQv0ygvasPQudG0aUC3WKpIma525eKEPnfA2wg3GugeN+YIM8UHcijQ
FAazsU0jvPslFEEH2Sfcgbn+Pp8WLaAlSQrjHKmN9GJltxaGMf1EKH5fBOB3dfuyyMSA5V0g1ocM
GCQQg0bj8G5ze9KD1aX58DDi6yGcD7ZAIbT0zwDDWNRRHNF3eDGtlaYQO0ZhHT0hoJJOp/rnUgB6
52eZtVvzklBoAPb4o/IFPibqTvAAMKWLMmusde/0fBv2vvBV38kJIcVihTQr8YKYJFSIFj83XEPm
TULCvyeid1UQb5kTq65gTMk4WTUr+TpKt2la6Gevl/VYhXvSvBUPz/xDabj7KEQSJHm6tIsj+QoX
8eCtBQesSNea4fvvXcnfbZ/dQm7YC2XNCzx+pY+HX29JH4zD9317f51JdiiPBmYFLRlxh75kL0uI
GKlawK1Di5mXr/mtEC02Fl/jePSWeOgxS5dZbYkwqH+o1S+NSadGqXbGXM4Uw9PiK4cV8u7cdgXy
SKsgj13K2x4oDSGvm45FX9UrIpAq8v9yShEDqnGeayFM8hXh/tC6cM/k1L2kTZvyqysJdUIfAH00
13rGI9pwtMX3t5L0iX8hpL1MGj9N+90UipKQejo3eekDbJBuuaRQ6U8951BoePi+yVhtQ2LmGNcr
yzSJeiSRG2rhllQiZB5R+jhG2abBmm9yZT5mxEcXnPs4lYClYYypYpjkP5PoTO0Zqu22NxF/cauu
ILBM/A/eU7gtUFTE9OjdsLU3Fq61ckEfxqoZFZ5SQQi/ZhupangaOJRxOVR3Gt6T/TTxDWN3uvXn
lSsF0GVrGfTNS2yePsPv9qD+zwUJZiXXT2cOKW4D0Wftvj0aJnPW40cuI66TwiWnBZsFSB2AaLRa
SB4tHFjUtfo4u5O5/DXS/EgFIsUUO/uSQPX05Qd6qLqitaS+lLOTaUJr1bdnPglkDfDgIHWMa5CK
pPv5+kKa7LLjN/7wqXx9rtdcgxFDqdVc6pndt0duWgQ592dsev/9gkMlnDz0PPI2ZekUV59ECxbz
/IjT0gvboXYqcGJlbpxDL5i7P1Dodd9OXncKhTgArlGWL8G1Qry/t4UBj10TotO9Vhgz9eGgzYrX
26JxeqyAZhHumSTJNt6pEb2E7ERDCmzgA9PCIkQT4Fu3YBqYZiDJUYjYCS7DfzECfePejpg71giy
3DnZipnj7/JwQBnWjRzHql9iHBpm1ypY3WY6Syt2vohUaJ6R9OwsFwW/UqCkwiSJNMK95ttE/zMh
VMUh/BBeTMmRwfKa+ClOZXaVaTreVzM2i9ccnpA+yfi2y4feMpznnx/ECviAPo3641hPvdsPXTTU
CghtnrbHFELO0f9bR/N8wxoILovbOrJgwvu2nfpNdTT7s26zMPjM7yQxvZE/fuCj+oarujMlpBc7
kW2foWb3lEz3K/XAt9p2tsPjQpmBb3vXZ3FjAPRTc0TVpb5UyC64gDcZaphXefLqPnm8nREC388a
eTb0WLtEwrzRbAt1L8XiIGEvHFB5qbpkACoNddnCpA8VPyUQe5fUFRszUVgXdyoSPyHK8XCYybBp
WoTWs/JwWei/Vt8DAyz+4zh61aEsVjrRAvg8OE9lw2yRrWtIU1zbvAGl6otXv4V8vrrCy5zKkhPq
0z7R6ASLkU4VBiNU7KbdEqoK9oouPXM+XiQ+RwX++B0vG7FJ+tJ0cWH2b4H7JUB2X2oUo/pgVhiG
8N6PBmq9tU85elUvw+L5umCe26gE6bekDX1LtnPClSpK7ZyY0+IWZWE3c5QWKPC2ffez8ZIh6wKn
VQKuHWyxzdODfHcyxoSTYvknhDxumYjW50VpXqGAKLy8Ep84Q4B7G/Ucegi6zM82Ihjn0B4rc48Z
DJ/htbAYDVbZi3zG2zVp2RxInlBdb3ThHYMjNu2B0vG/U5vRgUqbM9ZOU3CVcMtCRfYmpbeduiEk
J3xfQJ0Zfo3YZ+YwlenDMR1/E7MrurS+XbfYl1pwDkyg07h8CHCoNsyj/lZyTd+5X7Eaqy2UyBq/
4HlAepsiuNfbZ4X1K6L7znBCKltGXTvtF9xBFy3IeY/IDDjzHZBRIjQAOIg/qFJ0y5po6R0oKSNv
H8OouHLWN+y7EeMo5MQdPLxSlZa4ws9cUYntlajHxr622+RWUa5qi5n/SJ87WsMMUKyGszh1O9Az
nMSt6+TYQz7O+nm2RZ530vibdYN/ungwMHFEh66TZhx7esWgPvZNCCkVOVbCCc3OGafu9FI008iL
2ZXXMcHpJHV5O/oqN++URR2RKwJozyysoar1r623Jz8K7gk35zAf+ulw/dqNHIdj5fm9honpweTM
Fk9gBzCRzX7EpboVmwgcekZCYmDBiCJ0Nr4lBzw/uMF/6H5RExcHg26ziN8d7gVlpBg54FQXJezg
B9T6T4PaPc0SVXD4vyLq4aL4pDh0Qdv1sUAD07vQR45x19jRzwjajIw3Ba6Fug7a2ZqEYK1CoExW
vWOsoiA3AAbdt29UFUFRfk3IJjr1Gs1A60PkiDjo1D2pMNLpuK+pv6ai4C1QOGnM5J0Q4HpeyRR2
voE9Q6Q2VV4euuwOWFhiUW2iGQaegiPLFwe1NJza7wNuKIpm722ogECtbIWCX8bvzCZHzut6l2lA
6xM2pWganYywSSyFDDJ5IpG9YdrOmIxZYKkchXN0OlwDU1rFcfvoZjA00Df3i736NyHvE2NHZ3i3
8qtPlxYDBpetdEh2OwbvR43mNmF9rTKQca+YnZ82LwlLqnH62HtAl38fYFQYyqKHxnrkZxH5WnTk
gskr7i3cFeahT6OvSHtx+S+7vVOE4QyVnwjLcqSGrCYFvwEOm1eG78z4aV7c9A5guvmJjLwILfxP
IOPOYVAOvcIlwchcsfCVe7ntiazM+T9Bv4zny1m19sP9Z+5Y4VEBHzWjPUlY5PfoxBBWFbI/wYWm
7Pm3smTfWWDa+LJAxZScjTtCG0KACfIC1AX8AMKqAjSp2TsQHyUqTV0H2GH44/zUWYRNF9qiJUo/
bbQAs5QfdlWD4PhLB38aBOErmpz73yalG6Yy3TDrjLjwWS3UBehZ5bL7AWrCTeq3HVr702Iavwge
UJQiwUGrOCxcdUtZZiEBImYmeaBcfAG9ag4StkMMXGCDE8Mzm3vGaRE9Jdjl5ntlDhPdPAxU1SaS
vUSy+F2gT5QZ2I3jLhgkOChH+O7M49SIW30lBCN85kkRYqdGSoOC2DZAPRJU/z/SzSABMwImw225
xHxC2u8hBB2Mc5Mq8+oCd2jJTEKrcwEMygYJHkEMKSUjubuWuuIUzTUwLn8NgVdm6gx2bLoX7I5a
8gI5x68mZjnUjowZorWo0st93Hk/CKb29B87UU5SYi8RzdIj8tqsnRn+FrvMJ9atT6Zgg0cbslK8
smKmQd9jbnFdgHRQhPGwfr14ax5uC6tcMIZW8e82D2LsF4rKPFq4PlRCydk3IpLsq6I93lYb1zX3
nmOBRzRkACov/UbgG15fydgXJ7jQPcPTc8WtyXFC2ukWbXb0PDTnvzUhMCDU69SG1pTMLBmAJ6qy
t5xERRGm7a7ygmrmLP3j86KBY2etamC7qRbEq2sLTEqbpw6CMGQeQ0C4njnIFsrzaa59+j89JGwM
+WuWY+SDmyl7DMiScCH/qsiA16v1VF8q4NRiTWUAKnrb4zwoHyFH15OqcZ477Dk6w1SqOQoNgVOT
8Y3SI9ysHoqei2u50YjF1V22u34mSb7Goq05L5+TpOBFwVlOu82sF3Z8ymbzEW5wvsWFFqBKkC+5
FngGSAjcuDiosozTHjlaCz7KI+IStjP8vS1HBmdJ/LKKS5QYWB/cszAGgNgztPsYnhRt4YBoPJCZ
JAzaQdnotu6FFJri6Cu+M+vrz5GYsuGa3VYOyja8ltRf5T0zxBG61Eifp1v6YmyAHLqwtbITqeGM
LWhDE6u3DyDjlV1t7An0WymB8xfaB7Pb1DpfE33ingwk/I7UyZDM80LX3ElbqnhP05/5HhiXNihA
IFLuwzwVeSCAgty7DfPSZctIN+yAr+eShukUAfhYRGuEWAmmgwBcSHUN/nBd5DgTa9R7hPCG4eaC
QECzBg6aWosskNs/0BA9Gz64SDfr4HjuARjikEAfwYhr4LpUVrLhzMTfSQEGr75ZX+UVMEc1Pz6l
3SGxvOCQAjsQ9IiGkGTtjUCvTGB0497l2dnV8gA87NAg38qwZoitIzIYBvHqu1qfopy2aU9tOjR3
8C72sSQ1oA7JvgditXDHvTmtMoCKHlGC3YzIKpNDCOJ38C1KzyJ6goadih/zViae+t218dX3vJ8l
wDEO6pa5DD2+24AwCNQHZQT6AAbpuVPX2UcCLRNH/pnUj2DzG+HFE1lRo04P/WPBsM37UiafPPyx
XoSGa0N43V9Pzat+nQCbqOJK8Vlh2vujzNNMLJ2e2pUOwFxt8LOlW9tsYCHNxeHwUHiGqL85gRr2
d3FvASpNKrdbW9N7FaeJ1tVYGwDjuxdZZ7rFfBZmysvo3gnLTWWx326+eFpNMFSdVCn1+GMA/rHa
MXqveDeGUx0YhyOZPpKLPLbblLDiPzRl/NT8EQ9Or3lbxs9snUf1OpzoMeJWAZvkVr7IZFqseWpT
W3nSWBmReU/N8bBW1UQvXgM4dru7Pboy/lQrnW3dXkOjIH6rB70Q9ePrKglkpHn19+k4WKjgW0E9
1K8F1QNyt8shV215c8ag6jtp63Ld/aKjLurRkm0xKatMILxt430D0cWIOzrxjlQMF30cmMQ4d1o5
GXJgNtQBR0Pjhyrzy9RJVxOrWqB2nmOve0IeYT/Xd0AMBiju8fbs1IcyHK0apA/aR8Q8rvdIo/G9
tARqiG+1ZDXXeIyIUyy6pCz2tnpnrELdocud9n1M2j4sgVo3FvYTPluMzjV/Cat540ZRdUQfeDh6
TImh9beZFvnYP5VZsaA3KQYKDsYuGv6XqqrMqmlZJlI2xq5RLqJhZCpAiHeH/zEoYF4AvqrjSSG0
uE7xHiG5+3QiYWfwTfyKr8XlVeH8iR6HvaSS5ww2EwV22DXNcoCHdDWler87roAE5me+q66Yn+El
Sai52CC3iT/qrh5QSDIGmanOzD+z1mSKVRhVo22zh3148ZJ2wZEaA9NOmzFUwLeia2nASmeUdPI1
YlBOT1w6FyQFkTHa59iTA4ZlAuKCJC8dPT8mhgPZUdUryyNcDtVFomq7vNFsL4Aii8b1GH8mshy1
MzO/QIK1dlFAm+zOyJN4cX0xBzJo4VzbmR9yVf0+2zCHVxFV2IxiVYbpb1Guz5w3XXipJQ3C/sPg
ne32CCzCQE79S1GwKDplWsxEqNOifGVSrnXIo2AN0ZGhK25K4Lkp2UN0MYx1/aTkY62ZmZxz9Htz
JlLT09/B/ofnCgZ6qEIFhqxHaf31YeKUH1Jny0NPfdK7IxnHpqsl0ZvsM9bBEKBaQiau1zcbOhzH
uOpkgUvNXo0KjnJHvREPdC7nAf+K5ivlljzlwzp94Nmtw1SclmMfgyGb3mou0SUaNi1s2w2EK6nZ
HGZgTh/HAffa4NY/b55K4sBGaj38R+vzFmVNVUhS/cYDqJHMyYK0ZJhuauYFWCjhkPf8agQaB2Zf
Yg1PzKNW7aSXyCeYm5hChT+K2RUYLre5hCNnDHm62Rp4YopEnPtFqiYZqetnTO5YX0j/Q6Er+/Wi
y4F0muqqQvbu0TrMkGWjGjkzjB65zRtGQfVLVmogGUk7CdyIf4K5IVckRHea1ZBQ0wk/wXR7E2he
+7z+KJBPYAhVCfeVnynrEX5ixUCTJ+ziNb0PtZCYtxLeYhscR/MsYb5OWBihsFrZVL9s//zq0lXS
j68hg6xwxjCiVScmQ51bmUPZUPk6v00dbivxzIb9Zj3m4vgZ2HWid6h3gDjQG3hfCDTeUsWGV//K
tX1IJosA36rumCziF+GIFaQTa9g55J+hro544rYuvsxuQ6EpNFS2ouXKic6UzLdokQ+QYoQ9t+Xk
oDhUyiJBj2Jjsdi6jiLCyBSdC8nqXsYLXn+Mdc2CppHzuut/WvIbh7bQyIoMNtuo5QXKav6mxCck
etGP9DusZLyMYwvcSEfrADEme73J2kLBD825RtI4HK8FEg85nyenot/kmCrRZN6qi7GjfQVuwggg
wcKVFD16s+aFoBXWNIyO6UrZRAeZdjdguMq8rsEC0mAAF5FWKRPjbHOPDi3m76En7Zq1AVLlyIgB
cb9kFt0u/FvgqgzWLGh2HeSuF33sV8T3PQiI4i4rMOkeUlhs+v/6Vzo9OFaxefJ5V2FDNbReV+HP
34ngiyJM8XaofHzCThMrq04rjxgEQ3s7EId7Ou4BGCinxqDP7A1E3eeYlG9l1oxN2c0swDwMK35v
1Q+fjRJ/SpYyxZcVSxwUUc+CtKEDkhAynWQrVTX9IaaYDryaRGZAnSlWad+c5ZIImoGbxj0t1E03
ngHpQYVNqQrK3QDsUvA6jW3jgC2i3/ep4KHciBB+4mfbtLi1xpRTl/TBZMCacciVH8GPG6BCBr1J
tID8KD2r0iTYoSBwEBWnU/++opXrKGjtq+b3+sEXaDt1D7XSDJlWiIo6mjCxK3m2elPJenL81+xr
k/CQvCU8+kskgOnU9UnC63DcB12Z0lwdF47nyqHM2tWD3LHXq7WgNXN8KcH2Eh7bDYbvie9ckWms
WoCubTSX1cctmJdltkJerzjTVTGH2TbEgn6KERNN5Z93uexqWkclFCImwAU7ue7Phq6oGdxO1pUi
TjMvF7011KvT3d8etm9LTF4C7xUr6B3sd0tbSUjayb7G5TW9UyISTvXTRx1ebXWFjxDPMjG20p8i
xpVHaF5XQpyS4m2mTh6tssLedV/l2zBreHbNSlb+6pnwGEaHxPOvYmv2RxF6HqNZZdMvWN7WaY1p
IdCyniisP/tBB9LFzBL37z9pDaJx0s5OlNAZMU5DnHWFtuAKNPIOUjCbOyHKwsvQonC8oykhTuHs
5HYz0NwuVFHOvC9iV0BjRttXtaGm9qEM32ndUE0ycLK49YH67Pe4gzQtv9iiYnLyCwHkdmnY+Is/
iXGiuMWjfG0R/TYG2Kp2vNvkVNt2AhZzeYzqh9U3kZifNp0BWE8QlMfU5Vg2kmsG8jA3UgddRRG7
TtfLSSdKynxiA+FBoIp5Wv/67q6xDcBvF0YyhaKabtorzEw8m+IiuCLH5XxQBJFldCAjJJvvtVt0
FKOAH/abFjfoPZ4etLGewzz/oFqM/CwP1WllXjvYNGVoEpNI54zETXwevPeHClsQ9yW/TvAEhcx/
65mXWZWVPRmkOP84qwFG+W8t9/IHfu4/2L0zuVEHH7VXjiSoT/Is3XaXwN8SvdeciyqdOInJUiyN
gA69o2IKv5XmfEzntcaWnwF7so5NFKk4gfntmEKZ1Kov8FVG2Owr64pXsEPrbTG3jJ3EzdUvO4Vd
RbJHthPY6sDiN5nGFDvpu/xB2g8ylav9xjOe+nM3BL2Ykz64DzRRBMrDV+KcGJ926ZR6B0XMpC3D
Rh6lFlEhCEZcRUx3YPVYxsomdP14Tlt13iJ7D5NzgY9T6bFqRwnX/Wyx3Lc1upseVAtZfpRuxNtS
t+hRi+xJ+DuaZtpahX7eto+4vNGnkg/demjUNXZE3tWvfYyVfgNk2ow1LUp5tDjePJGlyXUJT1B8
NoUiCq6yuGIT6Blr6cQ7kbJP8pT8h62fDutq+l10xNMcM/Uh9SZDBg+8VPz659bwZE81BVSYwz67
HslpspFRQul/YvaVQlBisMBn5sWF0estZAEVHu6oX0iGcAAoRv6UKFhq6ZuYUC3FW7LNqPUlvCbA
gIzeg9QHVVu7A2fFgEQLwpgc6FFapUsvYk51C1UhvX/1lEIVZD7EK/Mz5RE71pPiChu+vG+ioNzq
iHA4hHkI/IyuqITtltzxkBpqDI04zNakQ0+gtipINw02oEzY6nbos7WM6Bojky2d41YKeldPSw+y
lC3kiCvEORlcjXfAgkCvKZXUiawSFdePRxY+q7wuvYcQNXAsReIrURg4aKheTgLJkPPP54YWoyBW
25pnrGQDkNsEhyZK3CitPolgZdWlKvvGQHqCJSAmUK8ibJRi9Gp7Klg0RlQbIoDUg6IyFwc1ZJdh
pnzYYqtv+Lv3Ejq8YiJwg5TFPVqoivs5pO1KwOysryhlyc/BwuVA/USiD/Xqm5Q+y049/NAFusHK
h61hRk+Zhkp4TPqbxP37GMObTpy0NCfZ571VjAYMkl4LQnoAC/vS028BGZ+kVCol9vbf3XORO8nS
Xuxy/BC/xX3M411tXeYB+ZWfdJmwVITCgIHSVrgV0i5qK5pjM1rZZvc+mOAUSKek/vv8+WlmLPEc
MtCuDftZCyB4fywFA7ExlmR5tJbo27r7SaW7k7n0Wu3hdj2BVq09SVkfOZVmk/vPCN5DLzN66fAf
LlE00hnL09LRbgzuPhbxl3wOLwpgCPPXwCPMqfThcFn7Zi2O+XizZC6sccsSjx7lgYzuao/gppeI
tW1uAin7wENX3gZrlVGUaRrEcuPOGHHDWwGEEIXAKtuNIxb5ncMqsAwhZC/Bg30hp/gtqt7fI1ta
qnAKojHSZ07uQxD0SIxTVZqFIuI8oPahiNEF1jMT4QhGc9gpRoMcZKxCQYQPuWuAVlYrf3how4al
r5NhwtetSMB2vhYo0yNc0iQECrYV5lyiRDKChaUVYNlA163vxYr4kajPxfYIbPZ0rXKWEzgsOZmt
UVFNxN42e5hxOl9c/cRFaqfrlHuwu1meWfD4vn5aSyC90dqMsXmlmH6AFeVkD2yL8TkqhvkQw+M4
I6x/cwmq0VjKUYBUxvB6rhrImK8mqlvz/MEskTld8BO0qzm/TD/ngZ9OS7RiXivTdSpRYOM0BZXv
C5ZWFlFtu7OdaLXk0DVIrYOdiMJQrs4rgIipFKk4a6E2sMX7v4LKVpbwkAcduQv9G+nbe2tEmjec
vwxlJCkNTrJQtx0Uc9kphnGlpay27In1Rnj96x9dpFik1CkAMZNXQH88dsKyXHJnJEV04higPYJw
fMjSolxupvoioh/F0WgeILA9BGsG8Gudqskf0QpdURhKOFbxdMXuhTkiX6m+VUb54yYZ8I/sGLF7
7k5rWoiAiel4Qs44mT0ilxgfbbLkkWBvDjJBvfqHYl6Mjcc+tqxn7AE9hoD4PF4mFRSdYQvAB/xp
QX1qjh7aK+1uD/OBNi3EMAwnCnFCRhW/mUF6BelDiOT5zKkzGJBe0mUEisTccsYVj1R12bcgCph3
k2/6JzN2Y5StkuI4FxTr+6uZ+/+sLyNQZh6bdHnyW680CaLOxKiT3TeVDOEQZwkHt9S5+9ua4AQ5
F/PMF2grt5wNclzYsKbm+ZtmtD/T9JipRq9W3pX8un6q2ZvAaXQHKCTfrJMV3V6cxxIaJmg7GIXJ
Ix+u6BCbikcJ/goAwJSqPup78XRF20hXWx8X/8FEvtI1HUfX0NgCSsp/Z6q9YTZd1458m3IpYCAO
t22D6I33yuaa6F8stXa1vo+KzpJ6by4kuB0oIjdQFaapJtLVQwP+07yi9PJLJK3sR/xdx63G8FL9
4jZhVJnCFoel9jLHEA0DD1irSdh929vkQV1SJAlWuZENnz0KXsUWUnOMdNQdmMdeglrcNBxj9LuC
xajB+BU2hGd3+QqJUVhtif7GSky0L7uF8dXVfbwwFLOvnGxNZlxAg3Si9gcuYU1RPZwS63Ae/qq9
DKG5B6KCT/HgzM2JwVUhX+Xc/RclofrXNFqi6XD6iqe0BeGDjEoHwGJkG/ZVq0LeScv3sKksD6m0
HrYAhlDDYixdVx4LanxmDWWUSougkCZm8Ye9/s117Asph0UgZx818N/cwC2umMFR8DQb8KnHmYaY
ZPTp2QpVzu22DWr7zOOg5PBnFxyqrtSCUKNhPHP/Vw2raxiEPJhMqP2MNuPk5ybBrWZ1Rtc9VVmb
a7guu9U13p8BRImdFyoc2BY4esIOC6YGXizN7WEIvKQAxv630QYrz2+SEwfKqjaBbIjfXvLaLTS0
3YKnEYf55Jm+bfHNYMtuXa+Kvx7Zw/+daMTjav7QHv4D7hFtSEZdfZ42/5qx1uIqzXQgCI5lGutj
RYIEBjNq1k9tqsnYEvEq3gfgA5h0FRZVtxdFTZiNeNN5v6bWeGKvp20ON4UbuaSIETTTTcSJiZQo
UF+4rFlogL5ijEzz0Tm0f+oAafYrvjBbMMVeYOBBJYKgVObSPeUaXdgEUXOGLNotU33VfTmOTL2v
9CEBIJy0EZLiCg3EQJ1w5PI3h2FnI4TtN2aK6zMVxQVLDqizJWglL41qQ1WGt+L06SN73sFvCQ9z
CCSe/RgC6ylPKW7GeskGmE8s4grkIq/QZcOtBR2NjFDpI5AJ4UOTE3G6ymGg5Jgo3gm653EOcqyS
1kdMjpThgVTPDYSSOSgOuhfb1W91y525t6L98yjbBaPH/f/3ovmHNkxRWPYTQzojAEsJ7KZsVvCb
gnEVkRKSrfGNccDg/TFe2GywaBxyHGx/6TXwOZ4dSJYuYXkFpNyy6ustJHM42Pe6DYjGxn3NXUda
cn/ylL3vzn3jeEM+0XG+s/SByRzq6H6X+Df6XCoDad9Q3JP4yDBuG7MN+jRmy1i8r0EJvuDU60gQ
6BiMo4xjicAKsGV0zfDgCqR7M3/vqFkJwmOZGbIofwZ+PWldPCWpniuYUmrSn9snwQbkqBpRNLE/
wf7BXQEC9E+gPTvrPwG/m4sh2iuICn+Feu2xzOOvGOA5opwOkO1FKk3GAEaHjZe5KfQhUR0olMLY
979ATHZFvP9bH/EKtbwziKL4bMP+ZvCAt8qF4b4PHQ7o1SEE8LXYs+TONBBg+3emNBIV+o5LQP2X
mtGx9YhAYA8YdtRqfO124KYnlnBvfpHsCSqjXy9k9j0CIOoscdpop8bYu0tqZs3WHuqgOMfr8svS
qZRMgcjh1+/iFuGuIRolAE9LdDK1A1wQ5Je0N+o2EBvE9yZvrr4Zcjmka7heEJiE3xC6s6gOOd/k
ZX72wB04HIhe4dtH+tphML2h6qcZ3iFhGFJJMlMHq/GiMiGBpb/suRjvHGzbACs/7WgC/eG2/Y8k
F8/nkFr8Xf4+wm/JfQOOpETHxC49TP6vgXMChne/xBPWHBtjwuU2C6o01zFeAqNOfU5TstFAebGm
SvCi9xkyNXbbJdg5OoHpHVoe2Kq6el0W7B240LnZqA87LKiiNXpd/BEtKP+Nby5KMf50cTHvPQ7d
ARwGWk8WMBrPjakgyxriFsY59zE6lpu2kzaymG416QmQ6+6XBjCSob4Gn/quTvu6zvruaEd4fWVT
PFWRDRSoBFOmB1a+N5wyVOiphW+q9xN8TI8RgZUj8sLItBjJeXB631F5wvsWBLZnhzzNFfVw3IvX
2dwEZwZb8SNHZq5ITzW8hhLGyJbMEKKUPbRUhsUn3W7OFCACEEQ06L3utibNjCaURbzHf1a4TMdH
yN0IpBDIObfMcNMw2yDx5EEYyPYV3EAmTrUna/Rn2sLcykl8rurs3WLDLHtVicKGV1yivdz8YgHD
Y1Yo7tapmIwMHTYLaDl1UdEH8P/CWIqHk3kpQSm3JEkUFWxngq+gLO+pKE0HY9SD3Gn7dpC8kYfV
xntt/ZAOg3Qhv0mrhilPxNdDvJ0f9SvnTfuYw8V5WfzOEIPYyApPiKsYEA00GXpnfXDWCSX7nus9
n93B/9ql3UVnr2IbcmsVol/JevHBW1DhFhjT1by2YU50rcb0g1MMMskxJpP6njcI4D2d6nn8x4E+
C0hC7myDKLCrIYdSaBDbFM3ADt3SHWYiLGPusvYq0pCvMOnU7DO+GhKftRamY54f8azUx1/3mHsL
7anpa8/sWmneqcWRtvbTFsW32vrjuFdLhSYnHfjd2mgLyHhSLclh6+PAZiRWFThoKblMc6R+hy49
2GSs/q5CXifysaCVtz+t8NvZw6MxH928RXONGyzae8cofXLe/dtdVgLYw95yISQ/k2wuYBFEMAY5
FoQhtGFtJi5l0TgczfjxNTLmJuEt6phl8GiXEekv2HDtPaaLQOJ0t4oZ91AYd+wA3Zl40kp4WnPw
hX8CsD+1MCsMNNfKvg37dVeCmHTPUXdloS7iPyP+qvw6lt1ATVkCfWxcBbsy+pBwv8iQid+kxU7J
t/F5Ny/nUmzMusHlZos8ZFV1MfcNJw9XmA+dsUtLsJ2fRw6oIrqwXP0IJ8j3duVhf08z05FcTNpI
dzvwUIZNc7Gqxjgoxl3UvEV3RomqqwUGc/OvOqPISeEuLgQIH/Mbu1S/aak/Au8oCfNHF1MjTKu7
8p0GitE9J/ATiWgyb8coN/1GLWcON+5ENxWH5hAdswRxpU0zCKMK/G8AqihQXYMS2evfONn+dts+
JOhURsa42r/c9yu6kqnDm5HxMolh2x3KoyLBF9HdZ1za3nBeEwq80Ogwh6VAwme+ztREsMtvRSHv
sspzghu0xdEnzvkLjT28Ea//EgRLPpgoMjS31ECxgdXjuJYaYxh6hBGFtqQQdNdZHjulLM3I5HwP
UgZJC/pBIsO9nqiUOll/OR34T8YQ2jsSHiRfD35zqMjYtalpCmwy/XfxEmyZlBT12M4q9Hma8XdW
TpcUBCfvd5hx9ITUZ2B3dIdXFHzlOM1Smkcb55rDUx1LM0my46p9sNWmvGh3DfWy9Rc3/pKj/Xih
o9LemuLAV8p/C8rshxKA3ODmJPrqCBvvdyGdOF2/S9jBf7ohKGaca/POI4GiVv+chwhB4I1Qfxt5
XsM/qw8CqRqeDNp9O8cK/zJsczxnbqFzftUq98H89W6b6373Oy6coHihkRlmsKYtkhYBwYxTXSgg
kw5lPrRvGuIdxQ+oXyvtd1HYHZW6f4qsHhcCSuOnixnLXhyjCOepiPyUQyaRV5BPiFtdZQ/BHVIh
lMQLkSZubnhNEJVzfWNTovz4wM2z1puSTpjvpMDM8ckkWSX1oGU0cbzb+YYabb0TL8mYjNgo/zgO
UyYw6+6Rz8gIdERZGaIbGnhKYl/O7w5/hk8dO2grbV5n8hXLW01qZNKnfDZ/PpQQVrnSh3KRZOXM
OdSn0Is5NO68QYNtPqIPE2wbIr8rzlfkDSYJdmRL+J2Lr7WTPR8Xwsuk7sH/juK8pU56TLZZ1zIK
iVeAtd5Pi30i7dcSwQM4G1MANZ0E6qrPp0aNS1RhtxmxCve75DidTYiip9w4ofebsbGjYMmolGW7
HXQrSt0mc8jhKjzgBA5F3TP1irEMjCO6Cm7SlaEob+2OyE4bWxsmc5eo9jU7A5tQQ2kTwv72wsNT
8oxGnsexAy8Ro4bq2qFZrhMn4HKxRnP0Uk1IT/VY5uYwsscCjQkdKORd3E0RLnq7/KdmeJAADls7
cdvzGwBo6csV7JYz/TlC1C7sLbmtPvI2J2V6EXNlCASkVKh3hOKVfVk3ZbrIdUNVg70Q5NSMfqdF
KTMJ9m/sIlikG4jYZO9gwSNrWnfJx3CblmHE5h3SrcXGAHq8o1GQ53Pt8UFOiloFHSZ0yNShIxk7
ggjenysFhA3DlrsXwr+S71KwZo04qebzaX3LTDz2orgQCNWx+ZTeM3DK6i4vhlQ2nNKIZhv0cfLA
Qw/ioIqRvfBEx0FEyFhNsXR14kzNbM6aWK60Cxiyn8yacbinYVasN+R3k6er7NLkMewlDAGOuiXX
y4v/zZt7Qr8bmNp7v29GL85wUu4HGQP2M+aTeMLS11T4fIAC482Ej3Pti0gjDNL9cRPIV65WXvn1
pcgsR7y/k5nNQtBHcn4oN5vDITugI9Mh647IdFMW7fEgrKdYNKxjFGsCOu8pfyfNp5Rhn+SmE1qq
5sWApe+xg5UzeaLGe1weNnXddKdipeYNeNepwMGhv0ReymA45dqBEuQxPtB8irMsugyqPW9P97sz
fgKhKVrMtwaq9tWdHdAXBNTNLQtCYg/0Dp5e6CW+LcxPNd6fNlYiVwdTG/h6VPjWicMj3Z4k3Cu7
V46YyK6U/GgHk+tIeTTt3o1AyvC7SdKiABzzQIb7gKiVj+m0uMAqp+ycu3bK+PgvBEGRrfzWJA9V
F5ei7UXOvws5v6xFJXtbYHGQpyqhFf+YkFb5aP1pxnXSXMxgCPK79SpzYOQjw1JyhioedxIgpgre
DxyzJ8it9cX+FPpWujIU9xfCUSORgNHNLNOSOqSx+9nAvC+rxwUxo8lU+MlkeM49xb7d8/mSj3ao
Zuw147DCd4lAPwbcs19+W0/YxOJpcOi8cYxAIQnjfJ3LV5dtI5S8ZG1V+eWwuGpCZjyT9NYEvuf/
G9e8g0bwWAEoXLoLoPylVz8q2W3T8TVis4mj7eN1kBguadFVH0anMLzYCFuJw72jDdx+XxmsFM9s
OiXYNfeqmxcSDPGdjK49UQc2uPckxopyN1NrQGgGsN/BI/t5L6un8TazH1iSqQO9+ZG9cJR98z3H
FVt5imoopImKeLtCR0qummhR9B58NyWyG8GaCImEToPUspfKcV1DcxwHWylreoBEH9dVnVIpd9k9
mgwseA3Nad93K1ak4XJEnbeqk2TCzIAnxPX3L6/8M2NmWAQBD2I1nVWRP0C9lYJMIpfdTMhZATV0
5nQEKH5+4JPBWW6/7LmrYjfMYY8TZOF1KmJgOngDR7jpaaEHbNxmwMZPyO9ob469xvm/4R0zLRSG
3b6Qpnbd4/OGW3E/KATYB8oeWSx1NbGJxxnIkv5uFThMf2ljiPjOz3xNh2d9u7FJpeukIQYI8rY1
GaNCiPcIR0Z4xs5+ETN6k5QN+eAFJac4xc7WH0eKOg66pt434XAMgf0zpXMi1w5QE4Zc2kJ9BGSV
1USIsK/4wKq1p5EagREfVB/j8xikJXKxj1wzY3l/aLbbgaHtIf0MPPAjAyd2NevTmlSjA0LSxCUK
rcR58cRypMU7vy285EZy3+qfU9GqcrHDMj/LnpuEsBefqcn2wrzgXLAZ3Xcuy/6q/yatciwCcNk+
Aunm99sZLMNRjwwnfsw2fcBYW7M5bvctlam3pYjZvLgZzIXN6rg/7FhVtpTgCdAA5ZINljr+H3dU
jbfsdWjA+PIIZLk0AklmJ9iiYFzO
`protect end_protected
