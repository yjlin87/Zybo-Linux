`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
jX6nBZHm/CZUQxtZltaoV45gK+VW40Fw+ETPZq7K6mCnlgNG9+yiA738Im33GaIfNL/ukQLYS6k0
jz2HE4GH/w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
LpQaId6uZu8FXkEAFRkCY37RhRPMTrJwXq+996GDjpR+DCfkl6g5wwEZmpYlCYSPKE9PyOttCRe1
LOAu+s2oVSQ56NDGpL8R6ax2m520Y3Lxkad7Sfp2Oe0san1XYq5rk4rvKxLogV2LooekUKKaXsgl
QXobyffDqz38XhJflzo=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JrqgfU4jgkjfBNPtFEepIL1EK3kcJcH1/Q8tmCFjqmScVflYmZksk02FdWt/AI4ZoEQ8r7ASF750
iFIq1dAc1M0eXLvexmqPOacXDZ/G4XQeRkSgdlren4dOL7K1zdpt3a0gLeUlricQpBtM7OzysrtH
Q7Ium2kD1Qc6RQwENjSw+4gk3KwWcyyqy0T8knqa/h2qc/NX+T9diE0/iPeWiEKkRoUWXnCdaaLe
Gu5Gp4yaHw1/Zjm4Ybo4E4hybEeZlB4kyKDRCb3MdoyyfKmoDLkPHJJW8ho2Fk4S7Kl30Zc+YRX+
UrtQHQ9otEQIPFxKiFwGHh5ktqUryR9DecGeLw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
vo6cjpzpOmfiVanKZu1I1amNNPT35nt8rvHrbkhdi4U0FOvXCo4uhOSBfk+S5ArVuDjqEPgdjhtC
mQbqmB7WYPzdsUzTcSeDHDL5S2iEcYCnGghDurLKBTTMIZyuuuxD1m63QJeNhXaYqXrTLrMkINWH
CwDU08Bjb2Z+At4dYsU=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DR25+jJlpcnSpvC6NskJwbR9pCuuQkVzu3PB9HUB6k4ZD7nyIHPyu+fzqed+OXSwDNcGDwIF27cg
GdRm8W7imRqZ9WIb2+0bNhwB4CpNpWjCqMWjGd4ZwJVrK1A9erBKQqpe6w44qBO0JwmDJuP8J6Ev
dKAOvxSZc+yTAN+Js+KlJK98Lw8hfxdZP2fbyidFVv6JqvhFjyak4tw5T0F5xXCLSauUYH0PbqA9
0rwMdlD2G4bSM6wewDfewD3RiIGnJY2wtyz7m9SUcCaDDeSMmCyMiG6UxslQgy7V5DC32LSPscJs
E1kqwPGAdbZu99dwb5oqzZGTLMIvCRxdgXR/Mw==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Noour08l0tMplA7BtaQ3seUlMk/AUEy1b0cZRxj6XLnIc/NDLA+GTRf2+PUC6bW6Ynk7j1/bUIrj
XVJmk2GGcYWPQu3EqbVRi8HXFTr1MyFx7AGxWJI1DYhiJPKWYKwHU5XaJzJ6ZPT1RHW3A8HMOul7
ArYxWDdp7W4JG/a+OL5xgkWR4avFW46R/Svm19K29d0sg6xAzFT0ODUNft9KC2A1rCib/cb2qeKH
jPhbdDowH3ze/2NGCPPYZo4agBnhan6Fh7R1B5DdkGbNFQVdNh1ODsyg3vr4912+YfeAY/+5cupT
fKup7waESy394xYD/lemURqQ+D0CvrvVH+udYg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 288720)
`protect data_block
Q9TVM0d0fLMff605TtemlrlVPTIAxARTuwhrQtP7vyU5Ujkm3joYm19XCCkJiuCLPifck+OgONOs
/05akuHA8nVVWl9aucXpHY87Go5x0jj/uNFVVikGPL7XvtmDths0t8QwaJD3gUsJtdFZcdytvcvY
uG5O5Np9udKe1nnb7hEWDJHTFqY/67TDA3uz2oAQbOakxB2m7Nn4U/7zrRi6HldtDZGsdn/nEXSv
3Vuz1k/xQoSPqAiSWlBbHWd9VPz+3JCCdsPAIi2auL9gavetk4gz6jfNTG8UEUWbB0eWtdeDKgx6
FGcyi2rDlOE8MWqjyQnor5V2OAoirTc3WGbuZcFrS4l9bHNBAgYIIp9pvyog4yncJRNyWBz8sXAm
Ge5xT6RHH1yHI0NeGE3cV78drW1jtbwDZZ0nqu/OxYNh8qm2vEHw9KiJemE1bnyQ3KF6imdZK5CD
AXyeWNZ0nIxZ3q89ingTfhCe/hbos7b82vxa4nhmWxYhrJrUOF7lTa9ihD5XPPWtuWLam301RA6f
z1wEoVH72hc0VMGbI7MkSzP7LxxTulXOE/5EVXGBfiDV+Gz5Vi2f6ik8UJtcAEQ5KS6m6fMA1Yih
iRwXWiMbsDez8fAyn4esdC5Y0d3OHpx4j3PCf6eCuEK+g2kFBE0gizlh0uYmKmorMSSs1iqRHIor
w4HywJXfAgR7DCC+nCSxM6IUl6ZEtqWlk/Is2mYYABhuQ/+cexctYLBZW/oAOlod/Ng3oWViEBWg
bi0Ro3yqMqT4tG9N9XmeeNp891muWNoYE/0k1xA3aLbzByWz8LDgxEFRqhPR+nNhtxVvMuDis626
M3EZaRUNoCSPyfX/79R7fCLf99g6fMWQQpHGng2B9kOOoby//IV5HSY+GQ08wZQnhygnkRd1CENz
SopwUcc9h8bVzYg9lv+ZjWldAr9u0+Y82nNThFUzyXiEzrAAsWUBpqGrmuxj+TUskrrSJMScSNOE
UXdAGGU6kqjY1+h6Cu+B7HzcEPTAfXZf+Pqqq9tMJr8fziOTRDG7Q4S1r6e7A9EHckOkQ4ceNZFc
OXWJuVt16f8X4yaKkQWIYxjA38gGMNR/nOyX2YJUPN6NVYmwdTN5BujaWwv06z/r0GnP43iwwZ1E
kE2spQPrL8YOgzu9g+s0uEwYWXh5TYtXnuhxilP0knk98q+83KyLpjszLLA8wY8BAYv1tJ5KOs5y
EnqMVs6X16xs09gd8KXKIAwatnTloGqjzQ03UhH3SlrzbYCY6xESJw78/ElwbU6M5YZwtgIs+1zN
pDf3DF5adjfAdgd/q2Nl0aS+vwQnPuasavYzN5vjgM1btdfQkbru+7r/lODv3VmvuCI5IXNA6thN
wGlG9xDtEm4eqn1AptEeKVddiGYeCLM30zmWVca/hY2geOAVtks7lguQfiM+e9I4gH+1vFV7r5qL
RjdF6shRGi8nJ3QPiKH2KcdsZ+5OJEjFfSaerFS3GHWDERZQKAl4ma5srkv0dqBOP88BYuo3xpOZ
CwfoOz9buhSXRAmULNF6istSPUeYjZ9fOvfXIbEIr0ourL3IDrismrM3ogx0yc9iVmUpjy5W1Gr3
Tw+rbBUJ8mwyJjs1VwyYm79nViifcqS4ZVb7lkk8SECXRH01e8aFrjH9/FjifrVX5ZvAtE2Uqkk3
imwyKtQzWOiisbV8d1J1L6iuCw82q1MVrmRTKgUqqDRxg3UOVAncyC7c2hSNmMw95HIjxkDNAgai
rkOIWUXQOAwWauO/yJjbYnpYe1mcSXKI0P3ehkLg0OIMZ2p9bRIaAHeGpQUN+twFmES8RUIr9CbT
0D4A1qflWWs1xSA9ChYoS7DFoWfV4udk4uiAECRuWPp/lhh5hP9YLvEkWCPXSpZK3iQFKpWf8YRT
BBw9dyyYGefBRVrA7wPG+YigeWQjVlJJyH9OZmAesWQMOA8x1bUDouKw6Uw2gt7sjJ662CzHIfgV
4yNe8C/TjMDoNfZ0XORGleyjQnsktRpbMo77hp00BH3TuSExVILoQvhuSqCFpt7saBewK1/dnYIM
3ULd87je0G5Qo9kJJADz/vfx3Y4StLmd+2GfrGaeXG4Pym2j9xRTokoiRXyM4GMGw8bcm/mioOPl
ZAHjTf/+GIuHmcdb5btReoIBXX9skoHrmZaaoQm2BxQ0EFfUXM9W6ZvEr+0uzP8JS9CTmjBy60R0
NQq3Wu20q0/bX1HP7Fwn45Q4GCTAnxgs1qN/VbB0YRj4/0867jRdMoq1X9tNCkZaRjKi/UZrqqiE
Eis8+6ci9coyCJFmEc3aMAXsWLuCPWU7JkU7GMqtFsf6837tMadBVNDTmSBYY7/5p38zwI6ty2J3
fviX6YCY1wsp/BChmF7DJ2BQaBEzoftYiIKbWSf6T+rOseL8BZhtpJk2kytHyUiffiXA1ZFe3Wjk
lj0pjbXzDOgEKQM9FTPTA6Npi1TlTdRyn2kC4PFEzIP1N4ppILZNzmRVaXGfSUVEmX8scpp2BPuK
4E8bqufMjSSGI0d+0YaVvqfbwyJ8/O8Kn0EDr8Oy3wEmQEqA24u0O2nqOx1EAF93bbr9O5hMZ88R
odcYUAFyZ09aNK/N0zVNNkFL6wgc2ex+KnkxscsgtOXTtftLd+dNFL0ALzhwDx9dpK0aMlCCrrzo
0A15CuqT6/QF9Id4O3vKJAq6nlxGhv+oXTJh1VfqlhPt6J4/ruHa9niJrR2J65PcMX9avD9j5qJT
p4E/EIr4Oq3O5BU5gyRDZAtOQFN9xscRa1zK4XYG8skMhwwjHwzyfJrSxhDBYWsMuj6ExabUbE9y
zTbuzj+qvexhRXtNS9X0A+gLqS/b3TRP0GRecr2rydufehyT7nPgwMhJDeuHHTf6UTLu7/dmPkQ9
wOP0+AYIt/MtoEoIUspUB9+HHQ+6gz8GygWlsu6htg2+lkCHWngZ4LGmtuFmhDMyGdgChbzi5R0c
/MQd7k/VgqUB2FR5/YCqaUc6nL2waWZzVDQPxqXM+QvEA87cUeK/cim5MsxhGORWMjos4E2837rX
OvTb6R0EJVZk5zXS1Iu7X13dsCEfru7BnoxRPY1q+KeGVrA1AJHykPEUTetb68FhQxCEceiWZ2fR
m01q4e4ThrO3VxrGK16FKGYruraPcbJcV8eD5hmhBGwRHc4Sf7PEaKcZAfeAtIGNlS394SdOwFl5
SnCGy0YaGBDxwK9g0nhEiYg+JfZNl9BLwcWHvWp9befecUJDgZNT6VALPVWo5Tob2apWnF96QL04
rEvFWZnTZ88HZYX6JE2gz1btNrS5rjDgBizeRzPR8vhwZA0FstUQHf93h0ngnzN8keu1rQGzgj9I
dOKTu8TWIlVySCcabTpizFz9SWLA6GOGWcGlJzfkTQMCYgvhU0cgx0R4z/hexmWvlAXOF7HCtC7p
mqTKRjkbtzMp90fkIDsywK3+R40bVExYUwsGhvpUMK371VzZXPgGdL4sib0NpKhY2B0KomsdQD1y
sn1HWBRsOXLAYu4mKAAbv5V8HL1n4kaWsu4bof05TMFqd7kMnsgTSw8jQmT99jzcMDTi/8YjerwY
6wPj6vpxFCc/17Tno7IoIV3p5lOSJQK8dcas73W1QFCuv2EJVXLM9O3mncna+XMG06powZkoIwtA
1kAYWM/WEHqStokAcOtQQQ/gGOeFM2qSoy3weJUAf4u1LWWDhxi77RbHhfe6ti5Doc5+jMAbknqw
F51b8a4TYgxbSx8iDvrUmFE8QLMJLgXmfi08UlmVBo4pZaiVwsqDQjk1zcT+8CeMUoHCDgFkvnp+
a+ntwvCc3gvu8vDO7rcxyp413fMAgmD3j+ZpTH7cCNMAHSbUAkuZ9V338cXKZwfE8ulU6StjeK9E
BndHrKdjFq7inPaigJ/k1MHSODDvu24BovHFnCSax4ZAx/ij5wGDRYWPrPlM0TqZqaTRtk4a+UMg
tXfloBgR0z1dKvQmjEW5dA2EtGy0/u41ZH+KJ+Gw7ifFdeKElsCiW1MeY3lbRPROlXDMyNnoZbkC
f4emMLoOF2EhTiyViUgnqeFLJEMiIIvXp6+kGdSzi9wfOeom9KWnNSruE3BqYiK/YlPL1q/rDJ3o
BNPYLIIEKWkRm3WY3dWO90Wi+QF21ZSLSpoywXRmQuzRWDhDli5tkodbh1V95rPV9xOs7326l1Hj
SS8/QVM7eqIm+XPa9EFbhGK5Cw5QstKkMGefzvfw24hFw1qmzABd74MPkzwp8GlT7B+2soCDo28S
P4ilnIzZj5v3YpihdNkazfNib763rVluDIloD6RiESa0Vxo6/stngdytXp322gtv/Bv7cScsxuEg
krm/5xRU9crQ5DARv+R8+ylDNhRCvwzz6XuuLNpF7zyS5o+Sog8L+JS9CLO9bLrknZE1ZFdB2xvq
fmlfNcRJOEgW4HLzWirkLEopXMwEsoh5yCfSXcdN6QaIdFiEs06DrLcQXVKufhbGLHHhNrbp/3Om
69RrM4/Gk0ASNQ0ypYdB3xKYY+AoOOeW8E10E2eoRy9QCgkWsSiIY47CpiEprUk9lTZ73sVVJ0L1
xlgzP7Tvso1c1oQmjJKRMN9xb83O7bTwCq5dnpmrNv13MhY8wlGWaozE44yESF417BPBMVebai1v
RJed50E3b+1VzL5t0dlFK8s/V+KAP5AmicFRnQrNedGypaTgWkNvvBYut7L44qlhq4G3pzcHeW/R
YO6iKdhMICULL4t3TwgS6Es4ZmLFzN3szZGO2d5l+AKz8i6Cmohv2eUBV8MKDADZYOauvaI0YOYs
ORw6o5BhHK17nLWCMO9BVD6LeHHec+ybDDeapheULN1xQigoCX83hUm2sVd+t7yw8tBGhLNSR+9U
+vgKSgMeQKEO/rhQmRX02A8qHBgju+yZZvs9lXs99hRfoL3yBWO8cMHcRy7p482aBEiB+UcQiyQs
F5shd68gKzahr8x+pPIAJJqE5kTUf2xHo2CqBj01nwvWHuw/n+iBj9v0r+vnKT2MitBJ0CYsILDe
3W747ozkBd0oDKxR6LG0+9SGT8gE3e2ArSvvXykZka08ceQqOYTSATPi7N0FF+G50B4ESHJVKGUg
T2M6vyJajbYuyOOI20ltbkWF2OAkRfy2kRbHNuNv7r/yT6urQrkFAtvv8P+6Np/sVnng+7gbK7K0
0LHd672qIENzrD53QBRcOQCR9OxIoEoi7mnMdbfUoQrRLmIjFsnjrOo7i4zb4PJt5AjTluod7wsB
zdsFX9Zs0RfXm08rJ7n+VCe9WpslMt8kHusX4BtpBuGG86Kv5vcTpjsy8fHVjzAoQCuZtJirTwWO
zZDpJzsvEQQgp1sGSHYLi0qmmIbgs+DiEWC8lIqa+AKWJSDC38wamaQZ/jDKjvcNKyqO2k5d3sEn
3zwVgciOkavujSTjVjw++UTrfgAizj9YlgOdwgVw84FPT0dCEq2GKKF+y3XP7PIK2Eyjmdb63Xpe
WbccXyXROdE+tW0fsbRyQq8WOy8WkNgi7ESF3DqYRvRFeD8UwvoZP1pJltpf9oKdbKN7wxpdwsfB
Wfal4mHNuxS4q+JawC26G75Xm9TUQ5h1tnXdChkPKGeo5yql5kwo1aW8DljKD35a8Mitw3gREXzc
kTkHKQJXTdzi9FPJccAG5fAVx5BukJFDdKZ5FSjf6z48z327XPvuMMyRjxJxCc6jtXoTojx7KcrJ
wMgyHuvscJDEZaOa4K7U8vvmtqxwjAwz+JJhbkou5G6958gY804uGPxHvI4Fwr02CMI3tPHPYm8o
G3rCvF/VwQKKZynbpYRz4ksmEQ/DieP1zWRCNOgHxlfy8Gs8XxKGKabJxmL7xutw74+qqM/bxV0k
EEPbOvkcsFaHEfYuPXnwHKLuwUDH8KCWj42Pa8Qgxj0kO/g0AvGstpVIcaAmPwFzYAkeAdvL4K44
Zo9H71T5ED7PCmpi++AmycjyZvsSu+SZf/5oMNs3jS3eNQmcCT4ZCEvZ0rToLhdoFfUptNpbBE+J
6IvKVYFKtuRn3yQfxwBbTgzHn2uFGGNtNIqCqx+uB+mf4lieSeRPEXenSBb3gxiEZJ9r55fNkzxC
2g7+LUD/R6miMPX+u+vMNYt472a6e+Yj+/7UmMBBWLrEa5SOKLy8d1MYQYC31FqzUz2fBiQ8m7Y2
9J/0VzUa3cxVo0NfB1oreeE4u6gHF6+4OYxYCBbn+ancC8w4wGzuv6+YlYGzfufy/8TbDC1AzQFp
GGZO7vCWvHQi853MJE9YicehTZ6+7jOgb9s2ZwLleDz+nSMyGxMBpiys1vamENmZdyMsVZGMG0JN
kdHsBs4yyc9D+Dv56Q98dTjwcGRx+08mMMV+S9NU3o72prw9btPgFcJ2MZW5zDydqzda7BqfhPp5
n+nrqS1cTo4yFqPplgB0Z+4IXQdsoMamSj+2ZMVMYdbvXpcTMULryqKX9UXtFFQoc2kwEkVwNA5Y
5YPAHCM6VV4wP/KLA0HupU+2XIwy8s6h4XFTXU6UoA70uZBCaAzVnz2RzuTh/td9Om19FUbpkP51
KGxFWUX2Wrdz3HRMEVbmubz/g7IT7YETGgDjWZZl+PtmcD1ZiEpwjxS4CTRkFd96L/QeP6RZob+Q
FNrvXSUHg9VtCcc/agkb6oUhA+etuON3iin2WlCM8KMigeoat2L3YTbTFMrKGWcvGUntNbzPMeVu
XC3j7cde2ANVrXs63mz+LBIdqyZqKwBp6obzo05B/o+VgLFdP8veFeaKcsXiRzlD8s0jZjRezUxx
HWdR0fhFPZO4EHYq3CvVEsvAYPR9yA0uSdgjNc3zQfGoFezui1cDxG5asJrUCuftLSYiHk98+9Xf
V2n/qVCF+nbuEWeK1zJmtLYg8yEeCuxTIJ8ruS3Rh5puaYt4eULm8aef1K8IcgIaS1yXDsg3CmBh
YIAAO7ICkE2mV7q0VUW9fsKcHrBtkTpEeEAAbfYPmRUdmmmQl5x2r0dffrHBkE61eQdSBNDzzYUw
aRA6OE1zjxsCLZs+xijAnYhqGG5/mitkESkd0ojRBdAyuAbE/aPvTtotJoTaB8m66xHjP/cq6XNz
Wj6R5KwpA+z8pnVMsf2ux068LS1RqWPw6qzTGknG2EIUrfyL/QoeCGQo6+mu2G5UGmYrXV26YPVW
+fnlW6yGc0JxfH/B+CJsX6OIKBQqwq9ZhvJFFTurMA3ygUHbONZ2q8nDG+wds3YLZLLCImu7DxVL
ZBNrcEdT+4M30pyUAmi4KNm1LbXu42kq6Sd96R9xtaVuyE9uHV7DNb4UrLFppni+JnpthIy3VY+i
1G2LkBHGyeNVdm+OnPR4hWcpHNcvmg30kRY0Dl1iQxef7xE8cDdJF5GPvMPeuuliBTh7jfK3Ti/4
AUUOAafLAghJthylfRLlM3nQF+x6YPz5FiXGIOICusDipq43s1ERZO+nwA3jgXT5jmESMn4X/fXP
nyQUJaQ9kbUb7OyqzLgO9sPA5bkH6ticG4cboyKlRHjo4nAKqAeo4VncC/i4G1ilL+KxKl/m+2+K
0HSENBlIsglJXVWbB6RnhDPffawbk6IRR4d2bJpiuTJivz0trSgNKxQkEZW8YbZb+s2xMt4cdYgS
MM9Ar53KkZqdqTzMevs6epO8UgQ3gwmIg7dfKmAvr0SGeMEKOsfVcIOq+kTD6xxTcfqdxXCbh3hk
OmMrOv0ievh/Hn3EBGNhiHUs1ur39+QupYZ+2x48sc1ZmSwZVHbKDbx7zVl94EVRQGUzwQ52qTFu
TRKKO105uLMBQK/SBGjCz9SP/+rKrjLeHMFkNvwIOaJ9G7jR4g/4Gqhwa7y1xiQsN+oqfESliXn3
hdljKpyZ+Bi1vgq+3FktLmyflm824+b03zERmYipBwFxFaISCPnypKX2/qrZ5wpbhIgO0npMJpJk
e7NtZ0sJEMtQX5w2gsYyEyx8oo+f3xNvXiOfG4HE9pkLHmTLV1j2pifAgHK2vK5x1TxxKe7gvFfw
/TJgVcftZY1EaAFz08Wr3raFGD+V/dd1pDloVYT07p6yvLRUzeChxg69OB2mMfHfT1llmewBfas1
wSI1f24dNt5ntfcUtwgCBvks2DdVZ5ern+0XM38g6k1lm5YcN4bAZ45VjX7O71c7YU6FEUVELPND
jj5SIFNunMbbRCOJlzGVHhjl+Tht6vbEkY6ZLCvs207Dlrk2nyk8q9P+L7hCpjllHEanGmuUtjG4
m6s382z6hCJN8Z0RkEQdxuqhgjMZmUye1UHOD9aHJUTvbeVxslG61kAsM3+yrZiY0g564Cc2OFxB
TRCMQxpIWWQptjpxkrjkGZrVKlGs0Nrdq02WpZRbfT4CTXc2HCb2sOky4lpxOiiVY298cFdsqpgu
o6yaqH7V/gnFYnQlokQOMbuil9aiy8BTxuU8r/pki4uHErrYb8Uvh1D26+ke+TcsgZc7GwJgP9l+
5QO8x1yCt4xYpmEJVpXGl9x7cBUNClByhP5993yYnp1K143ZoAcXVN56oa/NX55840a00u/R9mFk
KBi9IMiCJ8HxHlFjP74JOAF4A7hMSDSZ6yYMSZMTSm2iFZSbVdj8TWj0LbdciuA6IOR/IIqaFJkR
FZdlkrVBwXxOxQSr/kTLaTOWQA1KU45bofXNsyXBFm+i+/kb8/3bjW7nuC2ctLdRxFJg2L+Dgocp
9g8YsTV5UZuVXJnswWI7478zXiDjfHSev4CGpJqvar0ZPMNVwMY2miuiFbxy46AxYlexm5PwnFrk
5/Fl7eI/bHioSTQbUdEnjCMOUvLQz9DmhSWUbZ+DJ4Q76pevpNPlXZIRpwv9fCEXpcHpU5iFptYr
Ky7i/IIwfbmpOPd+VKu4e8oAk6HPJ7NU19KFtBl3PPqs2icXUWiroauXQ7lswwJ29/9L+k62sUO1
JzPsfFCZtAXKUpTEZFY9O0WpUOuvBF0GsQL7B6ELwlV+Ov94DJawNvezO03grMa769dX7TJp8w4t
WHb2km0KWIJjCar5HnYhtnq5gnK1DUhh5APgeYPww9k7EOJdnG4mfMw7oM8RD6ZuL7QytX8eaBmW
E1n/qDz9nUX8aoPnGDrXV+kv3wq8EBpEh7hVH+C+JFyGhj3X0gUO1YWkFR1TETiu8NR22AH6rK4m
Sf3ZjD6x+oAwWqSEPmX+3VlEvWIxO7uGwDIiBbs6Uci3xryNkAsmVYj/CueZ4Y/4LxkQFQMofxwK
z9agEA1Ud+b2q/CttUGE3OTjtkDRE70DFCP34cQK110OJvwEdg7GNVPswTNo8j+yoepaHSdx3vFe
RC6oNBDQDXAB3ZyHEEws04jX/fS9IcvIr4TVUtitpyejX7ETwK71qbqaP+HMKC+c0YyezcSAjKHQ
VMFrZ+uuQVOuHNeMum/bq+OspSsuAm2gNJ5HSCstfH6S75TZ9sguIrl1vyAes9W98ahdGhbaF4i4
C6taMS5FFt7Nk/FKMEwk64JQ00hUiyPh5etAKmx+XSdTcPGeu+nOJsvijz97OAmur+2IQTvEbrxa
Y+ocVuxaOyTaCPqxjAsrt67tGLKbEMs7aKprkxmG8SXS1Jr8nflPccVWy8lb5KoCYHA9cfYiAPrz
n7k2SCJ7lUyDpZGqUAORyeY5UjwzRjmtVleuj/6AdBmRfeTCANqw0rlEjkNkrwbqBa7fR+u/Df5q
aS5UGL3tUuujwZwyJSyGnS6PYZPsk6yfJjGZPn9SulX3/8XuTqhn8Tn5AwTqjqMVihLIRk+CVa0m
Vzc9PfF/t9jgBIDjGbt/F4366zRiPTfSkCzmnqLdGXzFI3pk5LBwufCEs+1hmnSnfPa1shkt64cs
bomWtLwzFM9Vq09ICwygx6MvvKEARNoseKJxnmGwLHmhAG+f6gD66NZwaHb67hcIpJwMYXJuzB8q
g5Rnr10pKlAqvFKO8y2VFA2YXZHHZQClVJNZN+nenIDMkWq5FVAQz4EcCDInjE04vNrbKNT79HYW
Jqu+5XFmGo+Da4CXVzCoEKniucDT/tlJQCpHAxlx7AJ1s1M1r+j4cBN0dxR4npcmQhzsUKhEmQc2
Wp6HNYP7mScig4mmbvig5lvEEEkwcgRe8oNTd3yccj4YmMoNiJHoJ5ZncQkQUEegQyqXVriqBf+n
4M7/7WmS5CZJPcRdJIl5O4CIbCZK8QuJ/Y8k/OAo6nt1xnS4nkE5ERZZAJASDrTYkZAO+0AFjAHL
/Mb3rmzfBVVgzgnBvAXKeUJLpobg8nKwh4pb7qUxaU41le6gFwNZRUEfR1hEoE7z4mE39mzT+hL6
pQmv9zK2gmgFJmfiwqxmfRK8ZbZiHq4ygBFHkVV4AIJTUIK3IPylpfMN6rEBn7vBwRuGAyHQyUQK
7Hm3m+FECVq3/w/weA2Q5Op8MDfXBQ65l3SiCLxvQkOoARzSlMsheVLZpxPMzn8gIaY1s8MVr143
sSWp4IXDMIRnT0MjqPbmG72PCXwu0MquYruZA2ddSoqyqoJ51aQYu2wrZN7Dbs0z/Kp7GDmJd2A2
/72GA1/UYJGKQ45pbjcTQG8EX3j1LI6RRfbWZYFogyCwYw51kPwZxAlES/aIsIPk3lsnwk2YWve1
MeFkIM1IHUIazKIISWtaOWH8JvEygpIKgNm3eUsqeh4wVXAn1VpsXKlZbjnzUA70FZbcRt892FEV
FPX9RRIyZzKOe1woYizaDHQSZ+HIfcBQ4fGDWSF8M3rDMZcLeWrP2WvFhnPEOqq4tKPFgITeRZc+
/L4NlGfTO7J5zZd3TrQtntRqCTg4gkVYdanZrhpvNWujopahnJ7uARXXrXFkProabr8chtpiwvSz
amJHkHP0McxJZI4nZ8ADLbhHVQ04efWlruZi0GlEBOgiyF8XQtQIPuDwqD/Uq84tN8gSW5uPk1O9
Nr/eZmBdvgqudKaQKn4JsOugD7KE5FtmHLUj6Lub1Id5vn/kUCTUSr74P/D+N44vMGjiKfZgEWZs
BwPAeKJp5lqZ3NsZKo7oHYFZUkd7k/813O9bkb+t4sKVzp8RnwtAvQP8KkOnJFzg9gQoQL0ePVEU
qanHl9/dAlyx7YhYS0N/pHpyuBxa8hMhoLU4aMsVMiNZxx8u0JFye4dJovA3ndT25OlVIsPSIWpG
to7UesnRaHz9jGClgxONN4fvMfzwqRojmFUQAZ7D8+kXj9yrZhi0iI9ScFFD/It5o0XGLvsaJCkp
+Yrr3xtXGZGSUqUDQhTSXdM58dando0DqLH35tbNoBxWSuhleh14zxoBHJBNos2Ns0voD8rU5+Rt
ahAo6GP3xIo9MHmty29LiLSzHt3MDhs9mN9R1OTcJcH+Wxj4+wghFj2wjsOQFgtQx0SxK/5tS9At
cEhK6XPuYxhNHEkZDbT7NhO4hwBZWK+3WoTrPxriE1uNboLABVGv59ftyKdnkYF6jefNbWvNzY9Z
ZqrD2LEblDmA0pqXzK2Uada3cPDQqpwQ9q1finoydGp/kazfSUyHX2XstjEZ9XLrlOLK/zmDaUpZ
AGpxm/ejR5Me39vSZzGgMaaxjatFOQZiGa2uYyCeOgXllPKWOV2pxav32iQFR8oIXFiWTddCfkDx
K8OvjH/2xnkM+FD5DSYM8ekIxZCAl8/AO8lj0nL+n3wz9R+7eKyyxXdj8FEveYlZeYr0cyBRgsmG
yeoYhGA3bGxtTqX8JoA+lraOf4hJoEhaZYrBCoXIzcHAaaxjPhEENTymMVFZDNH1cDKrWuxU7NA9
A5/rpnaKoKjEF1yJGYIWFTQ1B94IgHY2gePHY4xQ8uKwby+6AQSE+JXFLLAHPgagDYmogkBXm1RN
hP4xu03AZj2Oudi7KuWjRbo3Jqpbb5YOrxixXW2rvMSLNNTL17LDe0m/oRbF+28w1OCf3pqq4d29
MPr+Ylr/ZXZZkPBPrNvJ5UZ939uLJCZztEg6D75PYWVX3adQAlqu9uP8hPE+hVrM3bAUtzTiLUos
PPY5Vz3dZcYMNp3Yl7I+YoF9cwDF6bTM37pJVfbnnQA/r/uQavn2J+aec7ZqvwuOrb3HySEvi3Yn
s+jmhwhLTR4zbt3NIScWoQvLtr1Mb1RcKWwA5tWEr+3fRXgxzqQZ3ompqKKEKKodTd6Cuwdh9+JB
XOTQwDFfSYnArUKcZgNljyNsQFSOjlJsSqPO0gOcYF/OrtVpmSn56QoKGmnAiSpKtkOtjzrHyqo8
qWCXUuSgvZuDfR/0ei8DAlTAITphWTAztOImKqV4XjpYa6l26Ljn/numtElY+eAH+6rL09oU2OOC
J19u4sP5II0uFYbC/C3jpEarUzp0SY56dc2fESsRqhnNIIvG44pmH/DrJZ6kY8RlNrbd3HQLUp2B
Nf1m0pBgdOliIzwk0Z8XMmlEFrjYTAb0GYaBR/qUfnWWglJFdNNGj7/Xy7KW+VzkvPi2/yPBAIyd
YK/yKR4TlDLmurdG5lYYRj0ok5QJdjgTT9J/8K+//jhMtjokYfoyG/jjsBe/XJTm9op+FLpu58mj
JvutpanHZ5pdEVELsZz3FG1JCay1hjRhz1h2mKClqdg6jh5bbe3JwFzbPgPy6ShOjcbSv5IHzMS3
YKROZu9A9tKos4KfaBZTl/5A4NEvH2E4Shu0u9xLCkaZOt0GB9pE85uZPNRIhr5TSEWCLxWg/GOM
AwG3AgIYxe2R23S2paE2MjT4YaBNx9KJzMdcmEec2zJdg9Itd1gqAkEpVru93BisSWxJqGvrApdx
EmbLoFYAgjZgsjPNsBfEvUniZca3nKB1GJ8yhlgAoU8UQg4KCgRWsG0zDAwj0LIS+ja8aLzn2Ton
0LdmGRdWDQsGGzE3bda/v/jsCpYECLoXwgYbQi3shX+0h/rdJHDy4OFTvMmoVCcq+CMZsc8oXyhr
IXi9u2O2pFnXmPAJsTCJ/2mIEQHVxL8QiXpbgeYpxqn+Ce5IO1vutAwMowIhI3mU6yvSDIEp6CPo
kPzmd+/k8vGWUoQa8C2cxH/ywcDU+XI21Ivvd8Qk3arcJTZVdkeOdmiiauY+BxuHrkL2Q674J2Ia
xV8IjOEy+6XmOEt7hNBXrwD8vzjUTsFrb14v00GnXTurQba++l+Yza5bQz7Z/KnfugliZYk99wQb
tBCcK6i02oVSVzyJiUl7RocTbWymxWaPDXrCxm996KakbpTpbHqk2vRzttg9IkoQEeDJKiO9XC09
Tg4DY+BtpkZz5Aja3+yvqKYtfiPqNfOixTNFTSfL1SeqfEIq1fUUv+/2yns7IktKptmqm6dDveCe
15nL4oZx7twZ+4iGbcEvmHDeIZ3Cp7+/qigsjMeAP+vGzq5MPYF3CiphQ9toOmWEg+giySIWxmV/
Zz1z3DpSHOPXvBhqoUEAVbr50MSrqh6fCao7xPd1szoE/fDygkEM7jciPj91auwCCYAK+R2OnLHx
iN0v3ShE55Dam05eRgg5ZVQEw5VvPA1KWWVIf8/kbu6HSJ6h5VuML34NfaGDT91USdB8+6/OEE9p
tHDlO1CsI0+9ahprYU64rQ/AlqQvP3BkSygfRTOuBp2+7d1CRn7CxiFZiay7NTvzGQJ4dJSB4juJ
LpFP/C1bSq72PkBxLR23l0tdznOM9XemVWXzHPwAt9za3k+48SLvoZKQeCS2kkm1sNoStsSL/ivG
zsY4L3MV6s0lAibcURF1dcHvmFO5pcFScsf7VRL9Plc04+Gz6qMMBxXRloFkqkp3arlb7X+SUxl3
wrg8oLc4KGZ+RThSHSkwE0I8HckLt+6VRSbR4EknW59eV83FphHdvmosj3bbfUQ8zMHvpWapaguV
mKZOiOByVUZnn4EoD+LEQCXiKHBkcrg69sLh67j5FHmkwD9Jxw7k8SlGQKFzlqlclARlxlZXFS1m
lM3JNT39IEFhyKIZPRbhDbTl98QwJCCPCcVAZ/GNoAV7L0UxsxL0UNruLwONnQPZLA0C46DVKt3A
HeZYgkzIiAS/HFrs3vF4rNoIDlxy46bXnhDItVCOdzCTOCKJOcIdGxmcZYKgXmR6oE/2o5h5fZ5j
waWo37zbmLUwBTPmnLyfgI/x0f2iJHpmVF7AlWHQCQzvyWR0yfZKIYZNr5/Opr++OmtUqmTOS1V2
TNXP11z0E8T6NO04h7ICEf6jFDndnGrMjYA0UTm5Njm5PkSBKeHIsRHJOGyABmmmjXCJNN4leb7z
SPyIZelC632AlNaW4EJ+embuFJ5YxIShwbnNvP7hjDHF2/BvYOAobF1MKakIISeq2vHdmtwIwQ9B
T3xoqM4aVgRHa72oXFBESsT61JHlUhfX1Buczom2K+SriUg6guTdBw2Sq96oD3i9LB/+Q29WpRYe
mfFaHE7AcWoi7eryDvtcIL1b+TfsDQiy8VCS0Qx/LHAyEO4YdzeatJqREOJE4yDqv3DtqGyz4Ua+
7F1pBd34xDboRHusnXxlDE7hdnZudm+FZNwg+23eMh3A8Sm/ZXgIJVe6nvJXdEDe31R0AMy/HW5G
Ba5NQOXQO9fd+4SHZoQT0YJGuSAeoZH2Snl6ujwte1y8mGMbX62gJhh+XMmTOh3kljd61l2SNj4U
ObV0C8FGVSicNaisRBuw69TzhSbr110rhy2EJMtE2sfKTamcaj/+GZgjJVwdZpVaoEtTAzHfyOUT
SZRQJze+EZszNoZjgwsGpoaIeqSWkEK773KLYqwc1XjCUo9pt0NAp5H64KUMl+b44tni/Hbc0z1S
6Qr5CQqJ+dVB9NKp7t/PqQrx0z0LTHPHZU8cIA7UpO3WfCaAgliIAxNiWU/ir/t/orWvQm4Sp7H3
ihkwohxu/nwdQlRqEGSPqo4SLezAQnUPtSMHI+s5+oECNbL9F+L56s7+Q+BQES1GfLmwMfYNTLyg
tYpHI7NVVX6hFkxVhfKuhsbA8nI3QdKm/dxoZP4EJ98yYDWdbEWI/Swofu4W9WKOM538d3UmVmW3
9+zsk+w8LlKtJaaj4NPm7DFzAgOrN++28Pe+HgnG/QnZrPghp/5KrwTvOZvNnHmfzr1mBYw3AVjU
O0Qr2Gsgz9AtXT6r8Nsyl0epoe3zM9JFBhbZ+0KMjx0/Bf1P5cKsekUHFK/XojSP43PqjT66TTN8
F2W2lsd9488MLgbhA/eNDo2NtFez+cdnG68drbKKnLi1o28eN8ShQg8aZszoQy1HWno58ezUcZ4U
E1laW+RgU3ALBYort5bQyN3ouhE/fnDZ06V9NZEObIXiQPwZ9HmlHMUe0bjbc5TV7MA9F/LP3x9x
Eqmr1F0uQJlXgLS3tOKDd7jC9Q7+qiui7I2GCLmG8ats/I4D+myNCWPg3HhZ2SPDsrZXRCusFfAY
wh4fQEhFZH+uzVBNJ8Bm0MViG3XxVRMsq9ul7V0WdmOBsJ4Xk04XsY2JI/LhVuOnfslMlxPp3+X2
ggPs0HlLmyUnyelmIihZVQjHRBni2EE1Gs7qmcfqRPahBtawXTmoU8bGQXs7PGoesZdFdYT7cIsh
U2Dng1DdS1czFtZGDikHMCnvJxRMKcYp0cJyiNf9oFwB/rJsg8L2FarZnHSSy/h9gs3TowrqgYd0
fCT/CPv2/ELQ4AxnUrR5aPcyc3F5w9tiyzPzH98h4f0RQVPldOwZ7oh3/GKHVoAQXHfIqohNullX
/1Hy5kqwZ4uUIOGpJbROJAYQEK8m7WUIQlv+2SesAsK4ecpiiub5EEc+4NDJ9rAyRGZQRcQNQJ6H
1k1Md5wAQQt2xym2RNKhR5F4x0ST1zP3p3zU2GogVmUehAVQczv4gSj6wOUNxEcG1A4rm4hpT/3H
x7nhdNLhXSHjxOyp6NzXjtXetjpdMXETHIh5zra9/poIm9/BSzCDJF0c6hpc8CSG8GVgo8+7/f0e
2MIvrnyCKvmz/FD5B4MWZ7cGuvtcvgI54h9xrTVVvWq80hEA7a1wD2GwsVNwhUYeCwPkb7EeF6XK
t4+mEpmsFypCVKHkaDGTJ6Dezv3wrYehmmFvAp9UAszMxXY1ZQ2a0M7BUF9MC10ZxPaHVCMZQKxZ
eUP1fcJ++WKAkEMbwd0QnNGw2m0A3RhU1/G1hmeK3gyCmT2BauTuv4QaWEM75e0wX2YNr6CKOV9p
WolQ0OrlFzqnyj1q1Asxzn4iBTDPWqqQosXRTch0/CKWN+Aea03aT8ek0IgW3+Mc8AEJQx+78Ecu
IDqXOJRi2M7Qvs5QM4iHr7XDFW3l+Gi8foekJ+0lHaOmZnyJvKu4NlLv/cTOgnFbi8x+dwH0DKcW
sQSgKfpiXSemP+Ca8saS2gNZ/PXksMt97YD3CNS/V1KTtZHu/YmxMKl3YyS2Qx1uy66KSnlQgaGZ
r8j4yBQKdrgSPeVhPura3HaN9XBj/2m35V1K69QtkatZN83GLOw6uihLnejXJBRuENQ62bxhdlc3
7zbZAautbqXMa4UoTgi8sVozdcAKHtPxy9aXR+79/6HyB4WJFvEVnUf6a9lmpwPIxzt5/Q8+S83y
suOuJsyKJeWG3woh9hi+NTVkIF8R8V6/YA4k0OYj7cSuLOgcguTEku03Cj3jUB/r8oYL9A/6nmKa
sUILj3AcXX5dxkpMWfHKHnGGIg9ICTj0kEAb2rgyTLwKq8ADwvrsMweqMIE6Pitt7RmWz51aEZW+
4s9vicpPtJA3NjcoKpOYgcFN11ULDE5Z3fErZvQ51cfDj03F9gDPbRw5c+ZrHG7TkZkLphG1QAFP
2Feb4bOT5jaLAnoqf9VZHCVSMHNcx1zy5ME0xZO/P+RY4uCgU+WIPB4P/Cdh2vFNdSirEyYvl3OT
QlzA64h0qITpbFPBNygGc9Acy98w2smJpmjuIy94AMsQ2ky8AAjpAeYI9R0E7ogaqPGTs+P8LHsk
IgJYDZefZJo1mq5gf0CngYVnoWV52a6JX8JoFa+V3RqeduXnp4ZYKCog2a5/xRW0N6Dw2hM9VMr9
ZXiFizrfMJ2Yqgtaxet2imX0gWbSRVL0uRNrVQqJT5f1B6izylCfaxTBxlqhEP6lcNhvbbIL7ZMH
HYZuB8xScM7ifgacab/VcfKGNzkjQKU56oiInCu4pCjp3JxUmRIF4b77CYNEXGL4EmcNFSt3UVOT
VCeGd0YgFecxcFIQJRXYkDLgvxIBu8mpZy5sOBUysZH0BPBakjCU+RN2Rhe4EwL9/mQzVtjF+oN2
GqRqvxCPNer8h9osnrsn9AyZUH6RWS8adnv6RT+I6gaaDfesw5sspreZV5Dk252mrZDN2ggaZYlg
NfTxYqW2jZAbMw0N44fx85pY/mIoUZaAC3EsgXXH4mfTrJaNPfSWCM78TQ/vxqdPhtn07+jApULw
wS7ql2faag+FTwGh38jGCag38DYmDDyf6eyoslDDKQ76Q5uTdvLjepqBn/M/8ZmNQHOxhBHOa0bP
/FGFZls6W/iQNjGvfpCJiKgTzIKt21hEu0bD66+At8F17tE3Xv1PjYs+kXQSgACpTfgspb9lv1qD
vMaI5XDGpPPD6vPySG8iRWFHSGNNTulwDFVXAktbYQrTzt7cwuRZObSqQmVdMKeWoYH4Gecc01CX
FpdCzW4+sQ4jofW/skky/P5T9RRTBx+H7x/I1AhGvcgiji3Edf23uTY56/B0Zm9tlS9Jl2GmbdzY
fF1r8SQ0vL/rH9A983tCKJxJuZ4qXC99WmkMMuWhN3Y3xOdQdFkH4eZDLDURIzAKVhKQipyZ8DAp
G2BNZg0qW+0fJuHjd/d7Ub/oAgDoFCIlK3F7CJkNhJ9Okoh9GYL4C86RPBpF/s1boI7JuQhPUxDx
f27jrYDEqffBL8ABaevzy3cGcoiAwK/uqV4MA/+GqWrAoCYG8QCbIsds3Ow56YjwgYQPHHe6RRb+
Kt/CdWbGFY0XUINTKmARG2gnECRpizXCyj6JZcDjaMrKpg8qsomGQqJACsyyyy/QKlO7nxL6omoU
iopLV05i101AMEqvQ8LqFeoOUsTktZTzoAzGxZ8cEPI7HKZM0OV2rTsVgEni6Ira9EdlJP7g4W2X
Tk5/UjpTGOPxpAUghk9DZGBC/7KWsLfsXgo5hl1T2fEeHlOJgIAZKR5t+jpnljl86MPwCp3gz159
TihQe0XG+cPUfeyFbIdSHI1C/+ROkxgnfHGeEf8j/t181ltxu5bHty/IFevNeIr34sZe0adtopp8
KQz9Km6dWnS5CHc/WmjcBBM03eqlOGJC3wo49RWYJlqm+Wt9+deXAORXMq/HB0iRHOVO8Oqaz+31
uTpZsz1BYkk0QdyOdF8BCSYtq2brHkPvdkGFIsjDfHrBlScS/R8yFJnJH5abSA/pxXNMpzKxRl3l
iUrKCDD3XKLbU+Fvuhy07oXDxP7dYbk+BwbPllYVj4X/+OBEvvUa34Wm+edzXYY7Id+mlzYwU2tu
n6zOmWru0/mAZzapvCg7o1jHb8v6ksBDHOIwa8fnMW0NsSNpBorxFEppvgl8I0swkd8U/AMaolDb
kJiH71eNW3hg+rGQa1vi9gGYVeqL+/Hug3Ptw5INM67tJvmeYyycqbgfAA44B/qW6Ic2rtfur5qL
d4PUZ4bGC72XfA6egXetqKXyigSP8kfoOTGiTQ+6Ht7duDHZq/UArfFXrw/QM9xek5fhIy0YImxG
vkPCAn28/FsZXui/Izy+mAgPjWgr3gD10PasUI8MUWtYkoODE13rOVDTW4ec4FTjz5oloBWPFiEY
VYFWLhm9qW9PddDLXurCAqGdSw+JB4YHb9MJ9+M6Ck+jLcK9sEvPSsNJ4m0xOigQ/4l4QNsZODMG
KmaTXtf4xWrMQifF4xo7Xyzxqjfk6+JGzE7a4/oI0/CzhTAzXj45bXjXvWhzGDLAJBSh9iqZsnk5
nWa5vDOHMVrB3m4hujUf3a/FqvTl84ZN5mayH+wXUuNBlssqtCkZlnHFW83LbHZJCD8CG2hVM1oC
oWV2pPEzVSEZgSLKfOq99cB9kGnsFPaAARWlQRPReS4mvlZ4Vl2dz5ch5IPNHxo7p4NkMZRz66Lq
iqNDJYg02Zl2pLgl/BCU8OEvTELj6wNJw1hRQNE639L1it5Ur8ju1G4H1vfMFhJGRi5t4vYtludF
BnrEzRbvhdfVWr+Kh02HsHZbMAxHa1QEsQNeLVu2yhdX4y4Ds7FBeDGmDzcce/stuO/APeMPuNmg
R1H8Gi39UfMPWyyBLeCUkXSu43siFq0v6docvu2jVc02gdCWyTrnJmp+g8G1hKcrfXczFYyySccm
VFx60qxtR7t5iK5o27CvcvxWJ5gzjTApqoq7215yE2xBevpfY3ptwMkMIoFKXD7UAnsVuv7Kujpl
1nIKZmmXDuJgfyO7eG5z+qWj3a2Qg54H/iiD4wzRv+e7XcvkFr7lwx0YXR/oXUDtBOmdj3b1Ht7R
PxFgQC8N7gL3jNfaieP8KYY6JmE4/qTfLaFGHhcUZLKU5nPmaJP+/Is7Dv4ZNLbjxu+BDtezeJoN
mRH6saOUE6F+xzsDedL2Gf2xFvjVpJ6znY8OLwRwnhF/VhuQre9ZDTJ0tkFVSkVgbyeJFvUTEaZK
bPugUUQFSjgwoHpRfJLuVGChOwTvHncgOUpYqeBJJ5Tk4tsKZ+T99LkW/mo8BU1LfJ25E+rC4uxj
HVH9fu8ba/QheBW5hz2XuVDjsI60G7XFaAy0skFe5cxl5gl3EdaUQOtbSGSiRdTgWXXhlyyR2nUZ
6C4y9CSKVyOcAIcIYn5qNJPgQkRkthExjrIOqoc0xDtLH8WvwbUDfDaj35PCr8gZhufdtG6Pdn+q
FczNmN4mzhyQX4ifHiU/kAwrUcRElcu+QIHKJXS8/roGwGV9HORySvjxPowZG3Ov5bV40tZGQrxS
uV1A5e374jibx1Lg6dRFxRJ7oqAR1GJS1cjA/OUqoumIQKCbLobX9lW3Jh9/GlBQgAdYVXZRkSjc
pjYVgk0nWcns6YdCHAm680TgV9HUMTVV8kvKqYqEigq5Ih50M2zugKOWx4KGeniQzedxkYa+U1k3
6cHKfjnSCyel+UV7W1hLKvh+Q7qEyRqLrrYqq5UMpro1Lj+CMjUTajt1BljZWH+TnpYSUhI8qYSa
W08Ab25N6A4ZBvOA581VjKFh4UXHy2kdldJxVbvBxhiJM5LXceXhjx0w1QVb2aaK81ReALfhJHrM
Na4ztuC1DitVZc6a/tfotmzIMYOzm1VX65YlcdZuV4E8rYLxmqR7a7v7JgJ2QMHPFlSK0qVu0bCg
CCIKD1WxfKcDu2b97dKsSsz2Yyme5z+JnjjXNBsVnKe9Q40WNG6zoyuKGKydJbo5C+Zi7GZtgabQ
uNJjFJY8EqCl05F4FyL7GuNjvAWcSYUEoBFOYAashZdwlt9/TbCI1wE1HT8XyJSgVWXCFS6SzN30
JrWe5sxmWIiR3TpL8at0TDpibUIzAJPmcPmxPB/aLH9Lg5YqClfhXetpoNEHR3ipDwCbECbLCnbD
8mFmCjTRutdDXHn7iPlvjYiDllVPlY/tI8+EeJoV05DtjmU1LXIyRMskRLY3UjTAtTiBtoCup+8N
nvG9L1e8N/MGewcRKl5Go6Z8KW68XqpryO1xpZ8bai7xlJBH2NpzdJn33zYo52wh4+LXJGDL9JyV
GVDk6WNPO+zeZlCqs++9hjjGIGSJBwcAyE5EyofLttK7K6/Akquhq49fcDdnz5zoR08KIhgBbzXk
TRo64oXs911EZs2ymgzb2DHc0B35/uLqsTvBnrMcaZMrrLmUamv6SUoZnyL/+zgGkx8qLC9AHDaB
bRriZjMdNunU70NLbpIp2TXVP4ZP1QxJBnxRvCNOUNuDRYXC1C8qCGPtb1QvBJrMxKPjLisqE0Q6
klUQi8aNvm0tu6kJxMfdHWq+8gDlJe/Zx8v91pDgpEUjxl9uG22p8+P2nDUBLGKaZ6i1MCCjBI4v
NKRHYlL+qRHjLYAyT1+JoYVMchzK2G2+4/S5eVCxJD8Ja98LxPd3nw7plYX+CH07KG+txS1Mho0E
sSW30u2rCvQaMVhgXvCL9GYG0a9WxGFBXrui9Pf6cvJ56ESz9ZA+s6dD4C78+noJrLDTZ4Fxgzsl
1+zT4v/Tsd8DO/n89/+2IAsLP5PMnHaRhZ0oRCtvsngRoIgGkzEq1KEFFDaxhXK4JLJkSlSJlbU+
Uq1aHsIa2Ik1w2jlM+BOlQOQTvO0YXtNrUgQrJSdlV7gLDMYW3RJoCfXj9hNs0BoAkxlmMUarxHm
W+/US4HIW1UVF81yBMyntjo2RrwQr+Bp94SXDvwoqn0s87px5W/i8EFgwtctaESIMftcBQIDEh6B
h7MlhG35Xe1DYmB1qw9Sc0gvdVHt7v1qhgjlVVR9/pkEgvQPXCVT6gnMDoxBD7w95KDC7h7T2Owp
nUYTvUVA0m9KPsi3XvqB/ToASTQ6m2MW55EPKcTMGgG8jU6EPrQ+GwiuB7BWLlDaMBW5FkzU6+vF
m/4dX6HZ++HZSi03UeJTb9VU4RyEK/KEUf5xmIUrZcnQKtRrJw71C9uUdhHDytbsWyDBown3Mq+X
bNgYRs+DBS86z/rYXCJjlNmcqigRKegbMTQFL8Eyti6GYZztyClS0KIIs7NKPpAIQaV0EoVlAZoa
S0zE4NXk6REh+6XIqqxWvDRwGbA2K/Js3rwz8UnNVkQoL6MqmTYVqF0IEFGiHot95A+6U8Ut2Fqx
xZGukUkt5TCwMliOKIkTOQg+PwZM5ynxF1YKY36FElasT7q0xFTjq7li+zq8ZRXD/rgJfyBeQijm
zMOwOiD1pf7ipwJH0hP5Z43uA8Emd+tflepqvzPdNzpYDFDHLhuGT2IpTpSE4m3ZnL2rhaSrTdFp
SJidkwMPw6BNh+KPIvxpyqvanunfCnv8FDGtu1cfgHVr+NCEGzQkxppfuIrxVLl2I5hM7EYHgrXW
mhViOduSO0HilNhEdO20zvZm2fYcxzJtroPzCXEDHPR/TtSLXpF9nWfwvbfsrsMwo8FFo5gwhhT8
dlYTMRnuaXfYiYhJiHQpDS3XMZd7uTtM4Z9udvREI/ClLaw+p5SWq9q3I4C4FF7DiEmJBQs+g/H5
qvuYrUXCOBQzMDlhVR63xOraN11qrkc+eo94pOyRJfPMvm6R/Kw9+S5snGvMrodA1cL2AysmFdqL
uSxUcMhcrZccQB6lo9Jojg9D8nPYgU+jovL4dJTkqHO1x1QnOgdCMmdikhdYAMhVDN4ZQazt5/Yo
OqTB7L7VlRyfz2qj/SWyq9DC34LnORDkK8+BslVXURRRszrJaK3TDBMJ85uSCBuEzjilx+REPaeB
Zt5UmOWMHN4ruQn3V+Hc7eKptgk7aaUnKvFKDigxxXZ6+UbhmtrFWmT2NF6mzflVofJ7dgY5FJ4r
zCJ/0v216jypkKSmmQTC/oLTOY5CdKZx8Fo2KDUyb/N8Eu1mvdMxOXq5ZLmlSGELR13tjtBez7L0
u1zuIXjnWb+83Mb9NSV65HWOhYMZyaHSQgVca2+X0mQjfr+h8kIideqwawU1Tihr6+NyMPe01KdZ
CqvmW0SmcELA6MZeE6wQ2IsR23oDcCBYhtJ0hQSgaNvGqlKIvQBvRwWWG1RrJA7dgZbBRKCGe504
1D8UOeZ9IKp1DWrhXqKu6roy3o5OY94jRBRuiBQt8TjxSDJxhuj61tx+1BTvQ1oegCQHoDvUZjCU
RjKgeITrgZOVlh2elCedHJ0DmV2Li3gNULM7kFoG4gXEg+IgfuLxrNRXz4tZw2m+hItCFaEPuWH6
VWCgVth0Y0uyd/BV1wcsljA3E/8we7P1KZIvW8owXRCMCl5ZV3FabrkUf3GfYJRVUtdd1Mv8Gotm
9MhIhmAteiKPPxtrcUIV+IAjnxdd8PMFATj+p0wvkj2lyoivigi/NTvKa7I2viqiapmSwCuJb5pw
868I1myJExGoauvYp0umhT2hFV/3EKIg1Ea0AP27GL5IXxZIhgGe1iPGlpZkhIdFAk/BIAByAHnJ
kIJoteqyue1UeSrrsXlJ0mkrWCGzb45jwN+lzrIUdXRqZjihndTFRAiKogXsiFxbhDibtqhnHWbT
Kl/ySuY2zKJvtD0ilwbJOCgeDrQWDfqQZyhbEYMG9ddiv38v6aP80B4h7tU5Xqkp9s6Hh1ofkJeb
hJki9sSChJZVSItz5H1lgyLvY+NebipGeY4pIFAEp8TSJuJ+uyI68Etf8FcC/NjdHUYaqi7KtEPF
5RfguAvJoMqxTulN/jSg3RzveYMCAPb3MdP3EcBTDEOgWsVq4LjSUST4IQa3T2MCLyJXMyhpkL1p
Is5fIolqdQo4pmn0YLNhQdcfPx18eK59Xio3EtUwYR9CJELnNHXjkSemADuJDBKTex8jqVqCpQmJ
pXxbGLyZhcCSvXjnN5prKuQlOsDn5l59v1hbkfqVS3OOp7fR1dMFAM1aM2G88e5DaEVHispdbk2m
9VOp83sRnGbQvMDABmxTDajakHfSsoxh6yk+IWVJrewv1tQL/Uo8qEK4SGy5bIVp55pxbisEhBCe
inXeU/GrJOjKysJ2xsVGjsVhRwjRi2JzXa+tWd2P/iwXHOpllU7aEa5njk6QxZTKXUsYJ/yP96gZ
0ZFVYc5cL2wTqiOhrpYr2AqCWuhYvn7B2iC3C+2yy13sLCcf3CpTCcodPEi70WPBw5Xm8n0c8Aru
n8uQPEZF0i/TQ0M6SR/Blvlskq3edfP8NLqP+1H35l0y2FuqGe7nQP3+WzDLJsSas0bZ9CEzaj4z
7YG+uEamcMGAM+dBriRy7C5gbfF2Z+9ZyLbQdeeibBEaPb/4xdXn6xwCm2cII4BB6kCvJBaFtzWq
PMk+xSmDEpslGI79cSvMEOWfpi2ivgDSbdYXxGeiu4AKDyBYWKoHklgcJ8yH4Ihz1Tof5yjHMjs+
k1jPJkx2Nhaq53lW30o7MJZLYoyQqM88XN3lFlc0wjWDoKJZlgK13cQ/tYKLE7e0zVUhJ/OoJjB9
2X7UoSZvztEUtGYzvfQF36aOpw9QVJKhj8a84KFDAT+VnqPTeYBYGYWizRu2rSauxncEeaP2qiDi
HnU6E30cPMKCS9aVpgxzD5KF5wQGXVmiebc323UG2eXTZSS8j+gP8/SQECUsyHS2iueANpE9fKVO
k9TB/J1xDFXeZgpy7Ixhev3+51etkxQW9qsiOp0zuu+Fhxyg7eUJQejKYsdyspzhoJ402FJ4/ezt
V6mbF0aQ/m5ElGnC+1vls1A5D7BZP5Eugf3fZkgc9K5f+JrQ8Uz2HDGxP++xX28PQFZXcfWD75E5
qZSD/K8YyCm5EROxFxdpluaKZ2tVMCYeuAoiZ4VHbdreXOqaUUDL2s7h/xuV7G9CkNNR//OKGXr3
7J2QIBpkrGZ/rrzm+6y6PIYxgLTqDAQpajIPFmjc7jehcu/J0bV/8WrudmTVc//GKhN0R3jXHywj
NWtpotXfjKJp3JiylnESof2ljDfudCaZVGC0rD16C59vFJbFxNYfPUr1RlZaXkSNJMkHG1R1Yoe+
2Oszoa+u12R7wbnvSxcwiAIGj2JdcTO6g+XIumy/VZp/A7FLEz96B01u8+/04WSxf7SVZaVw3zhV
W66ZhXd2dOETNpsIOB05TU5fjjow/FYAPkufkJpXCTvyKTOnmzPUlK8+PZVrn/gvjcbH+TTHNlTr
LM7s21Gk0ZWjitBpnI87BLDbIaN0+O5cYvBDXzon5bI9WRDPZ++2CzMZxVmMlDfV4mzDEezr+zbp
ebjvKcsXQXpWCYeryZShm3TQbGucuFRGBwcUwSVDuWueGZiNGBgMyL+P6cnrvRdBp5cow2xd1Nuy
KY6Rk4BYa9bcY36paYhuVZeJ7D6KW5BPI/yT6ikF560W3jixrvoZXvs+VDvZeoaRd/VdZ7/vJefB
dUWC7YSAkFPyE0RxWRMrSHQQjIikrsEgT9KuMIp3HzoRTQXV187gslxyIQZnF8JrQzo6LU6og6tY
8g25MzzwqSc9HHD3Qlate737rDorq8QgE8efEzVUzYhIuFXY9AuAkCoJFwLepP9I12dyQo0LLUlQ
Yzrv/Cc04elp1So3IbTbwJpAxFU79XryEGJmHURdZ8bKjkqTpNteA4wRe0RQvYvTNVI7C0CWfIwI
XZf0XBmOlWlDc60DM2ZfcxvlahZ/IBKYRNopnnF60kkR5tQ5WkakbP2s8s4jqwh3NF6xcKNdG77O
qiOy6l0vdnrHGBDAgPyQMxGwy9pObeIc/Anslg7i/iUMDOGnifGLsRzTw3ker/+zn6ZwXZ5uIpuf
gbB8lhQGlEsL5lLXRloAylp5T3Rin1kZahQPqn+nQF+LHuOlj7Pbg0sCyESbO+49P/QpKlfdiFgP
nnfHCzsD4pk7KdnLCVyDy7Dl0ayD0xxauqKTTY/QAP2zvrKUodVJwdoyyAsIZjEGvhqwtHD3v3vn
diyXvpdvZtdBnzgdij+vcI8szGCGvfbFZdbYLZEGg4Wu1jVdsm/MirEarrq+CzLRafhPzpDQfz1C
Wx+Pe0+30PZ3UFIPjCQhC+9sSKUnUI8b4eEqZA8egcMwHYZmdZeIW4SsznhcPXuuVDhpEpR1gCwq
m3zj6lbK4SK9eWMF3xmoP3WOSeWK0S7g8DneHPsLDv+djFp2KO2BbBx1yYIxEq1vqfyJxTVKSPfc
Aq3ciKd6k8KlkVk2XzqacKzgClZbyAATLD6e4Ts8kZt0wk/BjaZxvPI4bk9MteK6UI8YhmF2WhwP
nzKziaijKS3o/qaGTEiadKh2FK0bf/WyUrSgP0K7NDd+9uQypxtnwVTpUOmX72I2rTvu7a3D/jg0
ffZIBVqKOBS4vJW/HfN866dxTrHQg57VfWRf0CQOQ17g3jg3dPYpCkKU6VbB1SSI6TYyfnBmrdWA
xXVS8JkgKJjilZvFQEC3jzSj+nBp94GiDtE13thVdhnlqxD7TaWOoP5mAF43QTyX/W+J7bJba/Rn
DAabVlnGuGIctYYaoB3wUleACFgij/LG5zW1UjYShNuKTJ8X+gdu/t3HkYy9Amd5gwFwBW7Me1XC
fjPQm+CQc3qQ0NlYAv3+Y3ULEEbVqieeAp8DHQo4tOjN8uxr4NbEKqiVGI/5OmSachsnq7NdFGUX
5Y9kfbr8nYbdRhw4fR6XRe2Zp0nKOX/9jZndYPzKimddE0Qhmir1tPtp//CRP9YFNcxhCRq8foEB
mzuSiIAHMAXi/B/qUTVY3Xtl4D3a33M87CwXPYg5B5LuE1HpJyovE7jeW6V0YVHTm5mBFbYT4zmx
3cCB7PjNK4t006mRoM0mMfOVFPezNYOj1lNPQDtN5xjz6sIvYjgnrsy0HJa/Qm3bOM5+QhWA6nuR
58YTDFcUpfzxzWQm322jblmiuXhItqOL15N+SuhxpNEvxxZRj/nl86T0y8jZkARQonXOiiO6U1RZ
wm2FQ3Dp7vSLku+4XUcANcX3gsaDjQdU0qqf3oJHpncQ8/vac9oAi0rljIJaYpnPvxZmukOHP6cE
bmk9mnrIU1/3AZNUpjQDXXzgMSuvDFEVSJ47TzmzxDdHQCul4XCbu6VKwwDVCIZf5VplP6pDXduA
Y2QZYRCUy4e4q1EJ9J72LRL1RRjRA+Rf028CRDNVeJWyn39PNxvKfEj108ZpEJK0UIfjwo4swNB/
u6nmLj3urH8SJ9jjqXqkvdou13of3exgRBabaSDqg4Bjf9ItChkRW0iwz0cR/HPT0ZYxd8K7VWD3
3AwCecjiLa71VVcBDyBKRM+E9I8RrQ4t1CubP9F0MtqkwKNtT4BEov4szQSp5H4kublA4m//niaM
+l/rIBtqk4vyyA8jnwXecVUMvopGRB/jdPNwdOQTf9WaHzZ1r5uRwbkJq6AXnrQ46VUxFJU/eYI6
1atczxK9AMdcvn+Bm7MVXVE1wm3AoT6P2lWC7TtRWqI4JPqYGkarNsgIqHixIUiozxWKxglDWuJ/
DnjzftvqF/M/xiWc/BEOY3MXF8a47xVFwGBSVACTXuinMqT9yCPUBm0jvwgTEErrRo10wn7XlPt+
L3Pq+LabDI7kYMxJci0wkESs2pwdOC6/56us5pxKxhqDKDkqmhQA/FI2pe5qGQ1KzLKoiOvlXWyK
MMknh6EeDbHxoqo5b1LXCsy+Mu5Cy4wu6jRA9KlBbj/rXY5fIIPsdBA2II/xAHyxQp8oZ5OFcQfg
m8l5enkzvAQ/oXUKdryekyybnhOIVnujQXxJ+lvaHQUG/bUOu8PTxmUv+VMdGigtJ2VrOwSNy2Uc
/q+RgDnsI3UsGltJuOjqErwVf+T1rMdPLyTnZ3gNbq6e7yA/je49y+uSPe0O9EDT6oRm6gS2dtmv
n8+m6Uo8gJy7hB4nEjjD2cqRP2N6Nni6oHAgSJ+htps8erlY1F4oKLYSUD2Me18rt3tyGqBkeSCR
T8TE5eniePUzdYTOdm+7g5jMLYCOnb5J1Y6rIDBKEcyjomhUKmiUnXWELwQiM/eeyjrnpYdWrM82
OFT/lUzbdAxbHWUUPDu22AD3D4F2r85YbnKVuIgCtmBKgmzP+INb6Q372IOdNxoo/PIqZxfMsm+h
GZ/1b4944wzG++F9kB7JxV3A/xK7QlAkHV5p/1egpMorVsYHfQM7IAHGeTWyKRrAS4iWRPD8dOcD
egSj0WlPLBCibzqO9jRSaxOowRJ1tXP0+enkBWbfoZwoCEyZdUmFdrA4YNCziLrbsVBz9FeNBJia
6HP8QcGtXxr0V7tqxhnGwoQfSp15O9MxQfqF4lbX26vj+yWQ6tFHNLzyzsSX+1vmN0ZD7W29xhIH
9gyGE9ernpwW5vnVMtGMuLCd97Dt9tB34dg55YAvzy4Ntpg9dmvBUsE9Ogu/6b4TJaaVRuNqrNtg
cKflHwqZoGZcqKVsnusWFgc50qi2Pbv0fkELyo2/Z/FXiykkSBO+oqtkVjDy8SM14ItPwBUscAIQ
crW8NjeUi7DU1gKrBqSmBlNpABXbJI92Q8hnZiAu1SMEHZxpwFRfJ/MYDs600TmGrIZqqfs0dP7v
iByd9C8MHocr0mBwBYlHEbEOJErJZJpal63OTnLwV76JwKAS94jR6+ICX32QvcZ937NuGTk3X49s
KlvbHVI49fomGa7/kNv8JS4K5nPq+Po6s7PgHMRcdR2K/XkdpHtBDv8SYD0epCdz281OyRs4noHD
qPJYnQ3cNHKMs5NcGtQjeIAKvLU4g7BUgcDxR8y/rQWsU6t17TPERxlYlMsdsJfQ2twapLXNXcbx
TvoOICqOMKeAJuhAgxHpvzMdLBd8/DjEWTQOg0OXMbHXTgQMjzootY2VLiZqJ5ain3Vl31Xi+4tU
prE9fAnlKExXEcqqRmWo+qM0N1JbTvU3D7raVASRJ95uAL06e5Z0g8nK2raeNn7vQqQYJqtFRdxs
VOYHc8lkcRTjQFz+GduLXPyGtEDtABXvDebALdoI2AID/whgm0EfyZ/tP1PcwoAbGr+SDtP/l56h
YN0IkHRZ0voLwT4ASa7+YilcstQn/3GZZ7aTcH+Ni7kaYQz8fwY7Ztcu5vEtW6+0YtasSKM1+19/
hn7mBQQ3WmBtV1CRzJMo396TYmRNRiGf3dxepOVydXfgOF3Nz0POeAn/yUcW5Tk0IqOcuPMBdn2M
OcKvIH6bY8MydR+/qFT2+mJdzk1zhLkcB+JMQRx3F5F6bRVFmu+aoQ9sh5oXjjXHgQQeMXDySfpu
nWBsvfhdgBua4Uz3GxsBwEUBYjVyrIJeUBnLzf5fEhr1oFRwzAxpq9cmmUJnryM3UYbuMh+K8BoT
Sniutyf3aR0VkovkENhvrcwoBKhwUp/5N0jESlM3Zs5Dd8BLM3w/pIN3nvOZt+Po3JMm76unSo1E
EaCRJU+UiuO91xlx1W2dyPD2x8jg22oi0f7DasWELu56AGkUpyXEgzzisUKIiwX4BqbSiVO4GjX2
jvetK6nhYbF23DXrVneU1m29vLptd76wq9Hj6mMGh0L5UkLQcZH48O6WB/f/urtw2WJClzjDLJFS
u6e6gXtjKVZ/vKFMAtO54xkCZjhMDHZPpN3FN9a8tVr+XoISN5r7DzizsHIkmWtUh6C3T4qfUjpY
/nFMFqAMz/PSbm7a0qxNl6pSxiMBlJfTJ5tDD0/OY3hnywRbUR28FZwPcCbwnMBMYeYh+jgislON
8teQZ1fwR8IBP5VfN/3xsXjO+5bNU999GDfib+njaotuSOnBI3HN5FkwfJNdEX4qFDobbNqefqHf
ZEVMhhf75QT5Vyt8FL4Y94/jaNW2I6A/PewJMFNBCiuLP6jacGRe3TCEw+mVFpmk59O7GXwVmMqH
G8GgPb57gaIhgZJYZfVVE87Xh5gra8o/FGSGTWBj5dUiBEjotzJivTq+WdZWP5w4ttBkO9zys4xo
7dwJNwqp5xafqL6tjnUp6oKuPRyi+iBur/vDUk6FvaSaWeEulZwAYZxrFF5O6aOnS98qOcrauaeO
UfCRB8rZlECi4GDK9PDjGhF0Uz5F83BjcImte7XGWbMLrn5hVs+79im14yj9TorXdVwkTxQVxT9F
uJLkr3bX9TUVNZIxr6TtCgKK4pORDfcQ8f5bAXuXO+uWhb+cWzVFVqfpt2EEmZZUFAd0Hj6mu3am
LvAJvzjV1IXteCYQ1OpVtQUQt03xRrGxyYDdiyTFLz14W0foI/eAm+akXZgK0bWcd0MHlYpjEZrT
AM1a27QSb4I7X8prAPdAwShcZ+ZgeUtZWqPH051/tyECjyoG9WnZoJ0OuDwl3eNuf28bL//72in1
iVsidEX4jCeJvNVqx2TI+ntLLvANr/aGuUuk30WJmXlpp/6OFRjtzDG5FU96tK7PtG+ISKXwUKs0
fh+ZDeL7VToDaUCn23EVyVWClYOhlAlUJFcvE62XTBnlP4ZnWuqUXnCfzNBZmKf4J5IFFMpwPpRG
zS/DMGHUFilRW1QgLKocqExz9wjVNO/UufBm6OHfeZss+S9D4VQERUX9ZNrMqMnAYbF0DfiwevUq
whYTyRKufPc64fqJpwsWdl+y8CrKEoUjWosn0Miaosc7VD5+OCYJ5QoRCueYriRyvqvbMSzqjulP
l9yhood0gAVb6UKSm/2GGIeWhooQZONRaqbozsA4hO7BgIcyvM+fl3UfitMCYzFOyS6ntFpkhj4r
uBQ7AANtcPQeeQYsN2mmHzTqIFuvk22J3WmnAQjzxdu6JjqlHfY/P19hZg3W2VHo3ow3e9edUZZf
hHnmFNh4jUDapDcIXnbYeeXkn16xRJoGWTzE98CbssHmvxJJWZ2m+qsNJIt2a5FVPApfRd5tG7MZ
C4g0WzeAjFoDYdh3tctzvKQYAOZhE3S045XA4wv+OMGrMRzCpO7FtcE1iIdPgMRZ6sT3fY/oVpPZ
WEUgInQ8t01eJjYWnp11lQx+YdWTTpqomkrrxsWW9zAsukvv+1amURLT1PBJ35jfvG6vo2rZb+q6
v5eQBHe2eWv6OpVezEAf/ngLSzYZk/euFwLLhcqsT/GhdSKykbJnEa1LMqnFaR4nGPSqpYvoCkQ9
LIURNPuXqdvDmOorVEG08uM/rIFZ0JmSckztL3rR1DY2fSXLEBOabUw39SMd5jKvs+DE1FUBCZS2
p8ci/WSyth/Pv6jr9dhFjxkrBaFBM/38qoyiQCpijsS9rrH/73xX/xhCClZcb5rHBuBHfSsiVXbI
dZ0cjSNNNFjoVFpJKaFVtUDLM1UMx3CXWotiHky/xx4F8+ZX5RMkXTQGJ2dWjqwzesBLxiBcVhvG
gqziuEAon1dFxKv6PjEgGEDLeS1MRr2ci90YVbo9h5pp47jaiIvckul9QjH6TwwrO/QMe02L7UcE
YxfV9MS3DUxi6fcKjvPgUIwo3/ow6sx7UGNNe/EI4T4CWYwSvrR/EHDjB1g3QzCljvzWVQKJs/ZD
OloFScXj0+GN0DqQmiJ9EMh5xnf3b4TthszVOBUaUbSTnBz14gKqgS4V5LNhGOk6vDyY6fjdC4up
pN5seZYC0UZ3YgJHtFsipq0ViG0aIS8fYvmrQ5Lp0IY43FiFlkhj4GOs7CYjnNSIVvtoBa4D0sPh
v3+uBnM1Gt9BU2Bq75sekTbshpwwMy6nL5JQi/+iFWo4hwjUwGczhED0Vxt3l6zXwWB3N3uUhv/P
kSMZYTbPMfILO+GbZmiSIXy9RdMVL8L79/2tafNGf/Wh5E8e736Z5+H3OLAogxD3xGt73yBO2k+h
9vHHk6DcrTsrsudGnmHg5p8BRydAREqK1dU5mYOr77G2scbK0Zy1uEi3WXZiGER2eQ+0rtYE3p7j
6RRk2dnGYXzwiTXVmrgdU0Y+EC6oU3/uc4J6UYK/ARisHdTIQEV+QukhipI7D3DAsn4drI+9Lm7v
73TKHy4rC80USw/dBOMK/n3cz7VAnem5nMZ/7R81GuEOeRjaScHMEq4oaroBduEvg/1bbdEIE4wv
SEbF85fIsbbtf/a2or3SeFy6VLo6h0bXoRgNIrX8BspI5nuo93u1UNwToRHTG3saBJdf6d5ncUeb
SYxDgaWXepTYPiX50MrN92+mon+AGkcOHDZXRhYfZfsBup8tZnsNqp9WG4Z/hyJ+MoeI62pnQbUu
SV/2kbjWdxNY8xKYRJScsAWNF4jDtkR5qTSs8aQLXJS8pfi1R69hLCsI2fMSCuL3gr2owjRsMMOA
lL26NaG9FMR7FgcoZij5V+9jL74fs4UQTPrFBnXl+9MdNO/hCcpaPRfnm32qi7eivCnNZhB5oC6W
FDhBHRnBI2FHATbbJXgyKehO78ZD6X7DiFmqt4zra+EmjgMEThezSiAf+3f4woP4Uvki29Xq4HYN
GMdQ7MQXNJ1Oq/NTzHjdVF/NQnupgN8FulvQ/PkRHUVPUO7hn2MgHLgQnp58M/5g4rZNHkivGhrA
aY4sHV5+21P7mS41SiC4hGidTjGpRnfEPoQShBOyniiTNog9SaLCeTVFvXvpfIu2nTAfbP5wvsOe
2OXx8q16FrQNSBSN66+OIqW1doXmFTh2KnTrMs6aAe7RXfk8vH/ULqJx9r+jV1+YiQvSBz37AWcU
AuYQ7OqPiU9BVngz8ZSbS8TVSQW3q9v6xqyp5jwjtPSCKho5VuZS05IH+hBebnC9l+454hNnVF5w
bNAc00wQp0ywPRI6qu7GN+p86PWuXiXdD96oazj+rAACxdqYoXJl5GWxuQ9Jlsb7g+nzPVTzpqgf
TCV2BpTYt62CYoaIESxRxNfGk3ip+xAInUyT3az1mDg00568806Dxv7s32kC1EelpIh53wtULnCJ
51w9+JvXuoh3hCqisY18+4QxilrqBACkGahT0PziDh4aPZkmiILup997SkaRzQ3d9L5ikktPUoTA
hgPBcbjZKdyuMvoahTzG6Ui2e/bLGf87IceYSPfS9eBwEzW5f2Hz79DA0vYHox5dOxRWQDBVk6HW
gFLRIgtCwam0PLlFlPqFtt1frLzN9OyQMPuJQ2He/DeTSJltbhLtAge4in3Ggh64Bxu0KrYvM6I1
8pT4Wu6ojNMABBxfUR8K+1d1sb/7tz0ZGcVPUTqfGVkbSKlPEawh59rXOYEiMDttJn0z2QzPp44X
7rOcWqGwKnsB3pDN1ZGzUO9H0CB68cIEqVKTJMGoYZzgdsCPS5NvdVE1CNx/ZlutATASxIvaBDYN
3112A0EZsEYT3Q0inLwnWLq63TSAnEdRS5jtnWGaygDyzxsxNGdUOZx50pU/uQK7JeSfaAggK9RB
x5n1ZVCohkcOndvxrUfF4baboKhxDtC1d/7sZC7zwFUFBI4QckhcOrG86axlXSL2YPQsm/5/9Tda
iApvW9oKytiHkXbVtjyBV/TQeL9bENiQ4KnfbntvggLc0c5dVm0n2PBtozkoV8UiGLc/TivpCJUY
AriMjS48Xb6p1md37e0ZLMOSqDEVm5Q3GlYLZ8j1Kq0cjhTFrUUPCyW644sl7pO1OSC0afcqMH7x
kFMKljL2HkhlgNijLkSmdCV0LaoIk0QPGg5GrStQuV12AZYf0RYey92JS0jGpI5hxE9gyU1A+huJ
6zkyVItbhK6gwW6joGgCKe4mOuLooMN6EnM5U9rvTtUYxxlrroFRU4FBWr0wYVy5EOIRS/nmeLuj
cm7q1S1q4h5qgudipBcF6afYbgng3WnThN/UTe0528eVoplt7enXhBiPLUNrbBlC/VX8TipwL0e4
/YCa0eihI5xBLhMhfiVE/X8HZtV2pVnAk1wf1YkT5Ls16PAr32KgxBY86RcVzjMdfPZklfKoJXRm
QkWFfseqOYnvuRUOsmr9rYBdJOQvl7I3QQFxscOfdknUmq1Tm7j2HVwqfIbTsyo4kBaNQcF9wICA
JzyXCc5TIxP7b8IOXBidqtzABu3SNPREe270jwtQJzyAm1e6RzEhPELifh0p+v43tF5EdqzQLn7l
pE/r9Y+nWFSb//rj9jNvdRmL/yHE5AMcqXRKd+YAOLbw2gJZMtF5dSQ3G5CJJPMhMSqUdzWoqSjh
nKjs1FSbF+AsKONJBqUhh1kF98ss0BytmvqvPkM+KjJ+if9vM6MnCa+HRKfzwcTMNnd5MMlcnFTy
2qRwsrul5yCQgIsu1+xYfr2D/PSCjY37mNRYSAYz54w4eu4ExbROfZR4o1htWlnfUqE3OQSqPkkS
gsSUQdGKgY0Kfq3N0tsFTBdxi1IoGESNws6+fdN1XXzpwevUmKbmBZkNChE1ED64hi6o/utECtjc
VWgBcl7PivDSHkRArNws90gGkbAnof2rThUslwl3vWTqp2W7Oh062MacQr0hD3x2k4u20/daYIGy
+vxjZzgCmS4MOQdWzQ5M+7nYJWoVHYu/4sOl6wJrayvUjBDdVlrXBtmDttf9Mf4pAXFXJ+DKGRN9
PUQm0Dio/JkXEQpbwzok9SIGO/dO/sYmmXbZ8+zmrUtjuIth/bVTCPDWye2wzgsiE7TPuG7h6HgQ
RLFoi3GkAMnL1rajCvEFKRyjppaPxUr0nFPzYboVmVz+Fw92Bm3twqsFFCk4GpzlTNd8Zk52+19V
BfytMu7h8YUQs2Tv0lUuUu38KbE8GOUoR68yfwceeA59N5B1rGB+2QS2tO2CkCf/7bTYf4vElY2Q
Y9cc8XqAdpjB07WlG8e9MV6CG1uFoHchbBhnq4JE8HIE2YT+0C/giVPxxnlf9Dydlcz3H72LTUZu
HVxhzjQHdW6gFe6dOG0+QGObYMXrQtQSPgRidO0Az+kdx5zzjgIJwJoPvS/fOlcvkmLkS065Iv2r
D3Q6fnRdnB/AZMVvjFUgSvj63QXr19BAI8KjaeARfflyanTYRPfSouiVywOMZSy37rIwoNXsHUlW
4+RfyoCooWRW3Vi9coFFG1pqbU99kymp+iemh2akVT0ikAuFrEdpeYhwWYg8Chh8K5iRAuBR9Rxt
BGgYryfmFDNNheOJufdLHpjmPofsdptxBvAv/noY5XI7ujpdbj+hmRj1xHadXKv9pJ/SOSiYbD7z
gCB2HbtSNACNOtxeawF+lbe8fWt8WQrnT9xAqR82DXm4VgnHs/PBB9uXA4350kEXGzXf3zKZMM9/
jSHchzQupUBECSub97FAeCcgeKB4cirr5LBXbY7KFVnq32q7ZlT7677AGy+CXfN58VwDY8RaODDf
ieWRfe+a50gmeHUf/J1bzEmOoDQrh5Nko3SZ9d10ys6Mw9fmf1pA8b4FDQcQMowleXwn/aOMe01u
bbo8C7A85FOa4+9fV+oZhKJiUkKzx3qXVQi10W8vappzfXVD+28+HtLaqrDt7eL4Jr3omwNEtUz6
KwB7jKyaln3XJsW/SPK6rK6duuk1Mc/cmLpTKcR8DumZ+HWKMo28q/PUMaF6/DNZtky6n+Da8SuY
333GTyAVJj0Cfo++b0dxtbm+1hRcprTtRTTtNfAUUHFpLnoHoiIkZN4A8XnHFin/V+wWIKuHPbiS
7gJrP7WddgKufQZR0mo3VLENvCYoDbduR4+Nwh6ZIZrVPnm7XmqGV3GWNu26UQHt8evQmLR0OJe2
/Ki25cxnHoKj5NggfVrlfgxvrI5WHSAg6IFD5elIOLMc2n+Ttvcf8WYW5lazTe/yJGnYtpUx/2zP
uX6rwSO0xz9/3sL7fVhJ7ubNh6n8SXaNlAsWWD57kq9S27Wb/L8MQSvagCNUj1FFvB0q2ZsHSB6u
sonIWD6aRbJ0zDEKYj5Z6gL2Ns46fcx/Cv3H22GLTx5zQU6Xx3dj11x3AnA64fBeHcsTfL070moL
3RPBN3psWmtiNc1cLUV6oebZ7Nxhhka0q7WOxFX+fQWXdijoFdR3AKj8hXs24xTIkHYErmyuCbBn
tdy/2dLeW96RNmX7hd4g/1Wgv7DUY+ycEjtUDzgC12RFZnI1zLmxzuq/okglYkb6Y2N3NeLWzps0
YyLrp9aC8BKE3gINvOfDcfPiT49zUGAZGx4wzVWtkCbEl2EnBUMmGPbJ2KKr0AQky+qrQ8TWurWz
yoLux7VVPQYOMs0VnJeIo0VzWTvG/JauTuinGMxZkVbiBcgKHQWAHMZXCNN/FOYYHmPo/vvgZUGw
0WmO+bI+TKk4NYiR/kg3XE1/NL/XQNQ1IuFZZiaqLm+gBS/ZpMM9MF9x0x/ywypClGq4qToprxYP
dp73Kuzs0xrGPz16eXcKGkupGWIqWS1XG4Rq9cMsDAs0fKUjXT+h7PqVjxAZ+eHP75wrIuATBBvJ
SVKOuMrXNAlpo9Ht9egp3C7+qQ5W/tuSaRoge1t28D5QMe7K1v7SORlAzfs50S2mW0Z8fWZrrhx3
L5aoumeSQgrmMvtaSvv0qEyV3POaLTwPFzuQnyQCsuurLmXpqbzvqD7LXcHSEoGwXdCoBgTKXqdb
PWEvgXrrzFOLO7d24UYeFeX1biBbV1FWvASZf60P7yLgHsffi19JV32YMU0xNgU6o8oUos7NXB0o
h4rIxfPSZyESd/qpYvND2IYYHVV8IUdyiuY1oSgt/XGJWlnsZmSARLUBEXjfUGJsooVctFEoxtET
mv78fuLZ/AiHnSKLIdm5isziqPCs5ST/Irgpp8Aae5dMxezCwl3DuajO/CtbWRmb//rVTVCIMCtH
CEQyhoUyPrCZlTafiBnWI5Uw+pyeFdk4mz5HSiOypBq0c8YJQxs1hu3IMSHLYOqqrKxaZ/D8Ss25
z4Np5w/Vd6aKprcKNHrisGZJoFHXv0ZS1QBIgRLzN/k9GklZjoSomBmtKa6Ug3F81cwhH4LnKIo+
j31rjhfBlKYK8RxncUgQkiEPTacH7RmW+ayjUZmI3KwTnaMrGEb1hR5xWiyJ4MBOFOZkiOynCiq/
MMFnDrZTvlh0rogHH8vJ6VvWNjxMzya1jCzZfmz9dqHyP/Qpy4VQww+i4Odws8bW8d7yC1cXtgk7
VHcPNbJ8eEOWjhpIAUQq1aV3kIl3aZW7gFvKRHoOxkSuKXcaxSB82m9oDYhlKp6UBwCYuL+qJS5J
yin+WHfNmJEyCQcibPEgxhTbuFnovDAhyD5gKCasHl5GiXOxYWE1byakZLs0IRD+fbcQbircuSTo
JEktslIySy4dKrE7R6VrU+wa/BGfjG2jBQnXiOLKoTEk8W5kHZo0OABYdZnUlTjMckGHl2IFPnh4
bletZdSbZgiBUCZ7/WjHQlsEaDBcE4YwDlHB5Iks3ru+zLZXKhWYoZAo4/9//tILbeXgHcmI6QU3
koG8jKhK82q/7TauJRo5Q0onKRDxNwyoOSnyhyb+fsvMOaSoGiUpvMCPhO65zKIR8jbDn4XU2D1H
G8Ktc/y7TngOJzAYjeNLwXvmbZH7kyA2qPbbH/nKr/yRjEp7AanjQnAs58OLdsWJv9++y2k90n5a
kAYjthPUJj9y6mfDcsnQEUbbHUPDKIXY5PVwchJ0M4ziOL0ZKdz1okdLiaqQYkmV5JCg9baKzt8c
dqhby8ZbFajtjwyfb1A4EpIPjBp0w/EhHwomUZBqZqP+CTrok6zQ+M3ZwuNJonBRTeNLfkU6+ZTB
FtiSl99Rjs0Z2dFJ/NJc0KQQP6KVLf478wm4F0UKGD27n6kBOZM4IvahotaC2ewy98hxuu3MLwed
FILa2dsYG0Rlo0zIFFnZwkvCskWiGDPG2QgpgXA3XoDUxz7fr3aohrOeGa2ENhkkYECSlLhLsDOe
6g3ALEuqY17p3amIC8yf6FYIORPGbhh7IeXsqyo3gw3q7dM2SGC71NWRziT9dXw9W1Hr4ykyDoDO
b1ayoG5uRgkB2RqiyOTEzhBreSWCnwBzHiznfCpu9AFHo5c7bhBi3bEJeU8qnU2tvfTlGr7f0jaC
Da3nV0YeZwj7ga/b0n6rYPlayBtrIiTkS3FRZcnlWnhEIFDKmTqpRUQCakac3s3lCQj7dLCS/GDP
kb5K6i+RdYMTYpPJ9Qj/6klM2J3g9aSbIwymV4ZGeQyjyM8wXoxefuv2yTDqCGLmKqArj1KKvwbR
I4SgJFyTWT569z5n8c22RN71crNSUZKONlVp0lPRxJOLb/JVEKdirc5JVRILFt5RPrU0tO+h5Xio
gu/QH6DMFdoghltR6LDo4gb5WBEcsh+femmFj9/Z81sfAv5xpHBhofCfzChZUZTuM6PX5cOSObas
x3AyWm0J1/af1/cZR+lGNFG27/0QHwotlMiNmtnYtboYSTZHoohrMdFZ9NvCeyjSc9lywmvXwoQ8
O3YpD7LlgsYzMycrcbffzbF39StLKHlAem52s8vF408/+s/LGpKxn+r6W3yjJX1C/mVYC9aCbKvn
+1wXJ3f7IbD3dLc8Ht803DQJaU6VjFS7u8wBO7I/N01lVtQs2ce88YZPhMLYVphYCnWB/4iROTOX
ySuzJna/1J06SYmNRVPeuPlqjvLSwU+Ffp35bNBXGiinWDhU4nKdgTBKAQLs3SLPCDY8N0EkNayV
rd7mdVfBc07vtjtFEZhfPx1gshVAYLvLaGddBArHIIVNY54ptekBWzwuOE3Ni70bgmcZvJ7fNoqA
4xLBZkz4bQBzWlrNQorDvefg7qYj9/B1Pf0kxZjxlPWVD/gqw3K5zfQwcgRKHYjVjF59KuyBajs4
luiOmJpZD40X7ra05K9dYam0Utc0VoY+AZk18ld5/sH9kY5Cove/bp0x0WpBdXmPD8Tl3jGPWy9k
ZCGQt8b7uoK9ti6I4SQ4TxUc+zOgpkDHc6FyO4cxNmGDemRVeDFtPCb568wfAuXDOf14veFsNlS4
E5a7qJ4Kz0KXyQZgR50bXEMUeFovD1RltXI7kBeCcMlgSUAWLldV62hfs+/+SD1q/QtYIAYlhZYN
FtwLu3q/IMNkxoLr5dBLnpSrR65Cxo8x1IIMYZxoMCUVMUn3BfLq2dm4rRPZKQ3qGTuxI0b9NBHG
ehFWRS0cmsychQrZI74yMWhFVPcbhOpDt7GpidKznTSd9iQZjegwbo+DF90SGASbCH7VFqGIl8jk
NyGvrCBXwsl0PBWH5mvvU8YGbvFqHWImVPREKtZdmAC1wcM9T7joQ5nCXbVgsOCe99uM8o5bYXwe
hyoj+oBjIcUYE1RKcXdp4hcb2xfJtg+z7hhs0JiaJizZHXHYsQFxIYTdX68rzfWB79L/xDsqWJF7
u4nR4YioHvSdQyV12SmH0cu20E/hHM9kM6Ro+8xUnPpZaJVks8xYWM1ivQ4D590k5z9tblQz/oen
6pSKpfHz4Dfv/L8KlHVH8RVg2knqNFe1ryz53u2YjlKzFtV6aTVGUPrCcMOksK6A0oYqp+IRNUMk
lYlqmurGmy6FBxEv5rdGeCN3MofiDTTtsaOGYHOyCSTkxL/HCmMe8daQkCQ9yNRKqdRK6oebMpKO
lDgJ0deRRD//5EHIi4ijCKE+5YgWrig8XGz+UmY4eNM/cWb6Y7a8Qzy8PxUuAvTaDY8V9hhwCh53
8Z8gX+3TNuSG/ilNcq4uUnKcFMiNiSUjl96FdZqzwK64IGScMWaZobycZzhx6L88tBUWYhImKXxd
1RLyVHzzwMI6beDs2zz6iK1w1iRNqvhtNXLhxkJ7t4LSL9PvYgDokIdeKXz3Nc5VMG9LnW+HZCts
BaljQKOcv8t9CkUY3PBBKoSpBZLpxv657xenBf1fMWgjdv/f9QwCIaikopk9IElCyjm/8P5FffK2
YUdTH1dLYNUNPgYjo/nPyHXN7AQUVCQRTQ1zb84mXpgy6+NS2BtHsbHqyaZRTu8bq0kGnPToQ48j
ZqJIE3ID4mY7ObGikDZlipTijvHUOoG1Z9HYDbHU9yWG4Sf03ji3nfKyqmdnTuaN4+VMHz4aQZmc
iMY0P+obOkIhTimPR7tdlYEvNUPjnp15FwRmlOTBpUDXjcUOictiMlEwkyiKfdMy+r1WASLgcCi2
Lq4Cc6Uq8pS60OQiUKMSSIn3/kAjGjbSCgEvEiosZ6L6VoG86OIngUJLDxmFaWn6pEAma1gbc/aZ
cB9pROvbp0UyW/Tx41P87vWsevOO6lJ2xImbUA2e86PbTj1g+dtnePCjIlp7tHXJMoHsR1jXjEx+
gO7eKjGEO23N+SdfzLl1B9OJHigMjvuY2z4VJC0nFWIeSepnohHn73NljV5aCPuHh5FZMGL09EWw
YEEDZiQXWeJqJZMS4rqzY1erC40cOnEEyQq9JIj2mQnCu+t5/XicDt7WviTbdjJLgFHz+6FdwBoN
6D1uDi4Y84nr4zqwuwMcrmdwKbHU6gl7+CkQnyoVjMPB/z9TCEm5jRkmbNSLKQdQltI83tWsaTNZ
YwPv+oQR2W5bnjPbnfw+mXNVVFrgqx9UxudbcvID4EmTsrQV0GHNcdjigRJobhO62IxDCJlLfcHJ
FXf1R83LCtSDmv/IN4lIJzJjo9Hgt/KTfq+RT3UZFjOZwEyHnasySr2RHw6oeJqfOsqa2ZxCzmAt
PwMn2/1LzM/dT0H42YQPElXOr5/N5ltZfVz0rUj/6n9lqVCR0uLru1qdApUFRAXvqMJSaZq3i7Bz
V6c+26OuRY/jJZnLsz4TBmKDVr80ZdELffaQhArRy56nEHAS0ljq1PdJqjXK/ufDthhplr62lze2
zS8AgBiiqF70M5723EwXYZ+kMQa80q6/v24ndC8RYn5q4TEK4Kp7zkiewM/yVR0uw8NwDlvcDYIM
dxTh+FzQGiW7NyDQL8iYiCR8G6h8OpT1orL+EhGE6tIMOFbZJj1NXmcZoICa1sFeBSylGMl2sqCZ
O8UfsyK7/jqWXvnEhtoLt3slkbbGEzIv6Ljyv139HbsVlD7UkPTUWGMY8WTPJ6gFirpPOB1yc85a
R9P5XkOCyRn6uQ+YyXqMwVk4QbEuaDytoD60x+xkd7gP8hgknn5AM1+HoZuVRQ8X/6DrD0RG1Knp
Eubngt0xxEUdHdDU1H77C2+zE1PZmi5QZKFRgL4B2x1krrSQ/RayXMvH5sjw/xWiNYU1QatS96aN
7OArS1cckcl7yh3JWUxhiccuDdRvF1Itk8jkYCnA1lKkbcy1yjDthuNpGoWj2dkTLfAD7o1lLwmb
5HpHw/vqt/3L37DKuLJ84R+1qqD8jSGaVo+9dX7yRgO16Gw/wk2KtHl4Sa93aE6J0oA6lVVn+yQ4
68j/f1Eyt+CyIQsdxTHgGu0zdiJYk+qcxWRBwq903CZkhBKREAntE00VvaMoitsC4Gn9QThRXfym
o/S417onZNpDTU60f3TyU3L9Ncw1P6R9kJ4vDkCU0Ny2ReHD37PB7E7tFPa9+bK+LQQhshQiEW1r
xoVdrMXtWEtPfBsY+T+ev0CnHbs2HKBMrlRE5oZY4gQebrtnQQGRnJs2liRxaTYE8FE1tEJVXpqY
U5uFF5MHT0wppUPhATgKa5/8u8WK3CgVnp7m0SPT6TvZK41eU6gISRmAptk4cHhsOF1WdBtfIh8v
w/hAxROpePgXe3acaW6MLg4BRy34YXbBkRpGksu9uCLFm7Bq0s4MdpcYrwyLOUW1Hn8mJ8lj9PB4
4+TPEJBNdu8HB6jLvS5V4BjiicuFCWYip9kdk5nxkajQn6j+j1T3Kh+D0hOqrtdJfYvCUwqWV6iU
PMrU5L1XeUtgri7YQQlZY6sF06o8+XhfMRaDPIrhLsUMRc0wv/USGU1BpRiGUEZSpEPbfC//aUl5
QPP3Q+0G0LS2ntNnVlfgiqWAkJmRG6huqyU6fehcwf3UUoSFxdtS+BflnXAuhumEuPoqGAzAhkWc
1Xd2+IpH4Pdd5Al0W7Tg7i/OgubyQqGPEMhNYnRYqnxW4Qa3txnX+4GxggDCrfI2aDZKuBTJs2Nx
l0L2bT2OIcae7if1YfN5JwL0F0RaY1oO8g+5XC4bMSn1SpLGY9o/sXrfvnbqzce/cyaUrS510nPr
/lLHbm6TuKfdfJzpx84YU6vIE83RKLXnFOx9vON3isUy0IQyHb7Ccyy3CE70TYhKpSF8DOyzqx3P
0lh3B4U+WodBES7l+lVuDRHjmJJ9CGFD8T0qXHw3/aTteZCR1lk36C8CCxwzExinVK5d1iSyq4uz
Tny70ft1fE2rky1bqhPAZwecyEIEFwi8DIcPMNLkzwSV6QcNY5AdaU6dA5uPUQfOfZz3OH60ff7v
6PCyFjAhSRK5hUvfYyvQLITPl5DWA5P2C0lURkFj5Kmmw1LRpU+phE5VNPIe2tQPhhHUfnlqSDKd
0+fClNBW3mj3g6XsQGoL/1Kzxl2f7IXBKSYTCP6R0ZxUn70YPbrcAckmOLzQHtes9PsAxGCkHUax
xf520ttvSwr0qXud0JPsInF8jZ02F5emoO2KkfXUSqa5esZjH0cECL7Iei0unUjNepB+IjoY8E76
O/u8gvJi6K/givtHwFXJSlCmTHa3AXuL+LYKi739rFkMd9JIN/SYPY4ZszrPtkzBVJrrAKLUdQUV
wCQEcE5mhIOe3fAw1hAY1jet8oHJbKgG/VnP5E1RPayGC67htmc1RDW1Cj6LSfBv7MfoKAdE2RkE
YuVtJXNSHsxpDtuKjPpyK01mHfXYzmciPageG9xgUHsZ5tZiddXVe3D4qujim2YqjIt9UgVkRA5m
TGoJAE/XtlW+Ocfx7HLg0NydUX6sW6UPUloYHXpcj8L4fVvrckzMQ76vAbxYM6mprAI82x2RELlv
rNaFFCR8azXxWdXuEB8f/W6+ub1bvOqrRX8MH8vd/N258vrViN/upil57i3W3o7XmmBY8q3T5i5t
HGAfqhrp9qi94wa/IdxHkqvv6Lce6hebRw8uQheaEtZS6uqzhCS5QOD+vcyg/sA/equn6AXd+aEs
1iR2mqFh+/twLmgd1kqVZj6H9+2b5Z00FF2tuassNT7h59hRHBBewkR2mdvjC7njPxjWemL5cBvx
ol0KANwKa/KVgBNaUINqzWLTl2lLaRvZ5+tAINOqNi8rR4u+gIQ/LwT3FhsNgxbF/73sS+M586Pk
t4nBxthPkFeZ/ib7f1KW4AuVDjHeJFmxA3t9rp2efMAdLPyEvgArhh9xSqx8UDC4kJMOeiiPVkyl
awhcsi5J9SiCZ8+pbDLDdCM0AeDTT16vNe4BxX2AC8fRmFV8Rxy96AHu/00n43UstNWqYqrZgsYT
rNrCYkvsCSOl4+vnd+dPGuoOsKC1wqI0EW1IF7u985dWXOaMCG6O5aeAYqkedrYb/Z4Sv2nSXR0n
pLrx2v6geqJItHzvVkapc7Bii8lyxy7UpCkq576Svbl3slj7p09gbJRadTv0tVTbJHci0xYcCDgg
T1eZLJ4PtArF9zWoEBL9V+qfRqpai+JHO5erFWBPKJLQl4vOygW2/KKaqC1COOjCMzMGt9+hETya
XGcMNoBe24C2zBXT6azx5IjE1evjYP/QETcu8qysp7FtsmA5Ru5jYy3BDrqkdXWdSupcjU0i1AG9
BVWJQGYVXG3sPveohzK1cvoifMdRK7Sfdt+h5Bh2oNtgf/7Smc/n1/f6RFf+jSzeP/a7j9Wf9+Cs
DQGFr+CWsGBSbwa1mV65Y6JpfSFxWEwGM55hSYCAUiViR2F7RViJrwY+43ViydIKaVjkdIB1jQh+
LTrmiApRGBJNBv6EEFjxAnpBXYUKrWuOr4jzgbRpiJBOadNSxXsJ3AAOFfVgMa6eyxbMsGCn/rmu
QAu7c+K7a0co3zc95a/HLOh4onqCmlJzL4jd/o73+TNDxSoKkMyfULVo57bqwo6geZyErSE+Mi2a
dz/lXZbfDzwTYCod+YeP3F8inMchpqsLgwpT3eM+KWl43SzFg7t6K7+XLHYgCsuSfD9ZaU+B9mdv
WpcQUZOyKgcZbM+4bCHaSxHVQm3ezkdbsvu4kkqhN4C6AOcgOMO4ueY6Ml0IWjGQUFtJ4uCbQ/zC
SUItDIjHe6wDTRcpq+XvK6z7sSJrqDLmMo5GcAA97/BfbecMtWXRH0lyl1xN+E2nzYrnERF8X94D
RVzraF9nFv4XJaoqGoSrona/nOcKj261i71Eo6XFIsqrr0GLF4xFhZsRXeqC2UoXDKo9BbTjCNF+
hN+pHSt2wR1H+V8qut+W0D+eoGNZbTMnk29BcVuFOXwv0DndwqOJDG4Yo1prCpohTSCqstiUs3DD
sNFAMGjSj8YmXQwqazkcJsj47A9xpwp6BeZkX03nmNeoHcsbeUov753FFNjP070+Cn9ic6zNudze
dHcfxgjxeM0TIFPWdrFUnO3nAzsDOgzN4p2F6Gybn83QQhwh0E75DdjZWg1MzmVroKS3cMpOgx77
FRsfUNYX40EH/HA7gL8a7VLaO6LqWdZr3aBPl7Yr5Fc0qJAFtRi0AzE8uDghHWIwqU3uxcwza1uT
PdtZIutJqKptUY4WeqNXplonrfxwu7SnD2xEo/D6eIo8e75U0DFXh1o6fmm0n8XhaL4SMlz+kljh
7jhO5vMVCeic52KvLPbtL+MMKJ6Rxp9xuBQ/1s/jGZ3EjqlzewqTC8oSVCB2qrz+ZSTENI+NA14O
0oTAqzWx8asqsKcxoZ3o856MTTWrFYoLw4wW88czf5+qvmL7Cmx5TQSelblqg1fip98Eyu+W4Yq8
Tp+djtledpoPMKZQi7jASxt7EeUVRS5E8G3E1fs8E9w/Vhl1w5L/Sx8f3KtshO83MQnp+d8WygIo
E5sBo+mKWvl2RvPLKqVyR2UJiam05RBCVUsq5HWzMdqFitCmx70BnvB6knqiMgLJsjXU1qWBQxCY
NAGSa0UWd9pZhElbB9Afquq6zJkkiSk+rkdiIamBXgTnvcy42siEIyBosFCRvP3hIne4YOt4L4HW
0SmuaKx6jWBe9CbwtxHjuVybkGva1uTK1lnRs63dUrpai4Uanbm95tVbKmaMmcCAtXaplFeP+LgK
dGjzspsr0tUOlYmASXeKHDMg+DPqzcQ1phwAOVywUhdS5epWgaCxrWepdvC4DaKfsyGdGtBGDOYa
uyRsIsyL9vEcTl5AsCYj2W/JJTOKela0d8xP5t40jzQOe3XWodCAoXiYvlZxRVUQnLwvREq6gGZo
gKLcpIh4hfXrbZkH/h48/ovjdjr84sLpZY1oFbeJOv+Bo1LtW+j7ZVvFiiCkoKZCaMT8f6RYbBWV
d5ehcDrgQDEASozUABSo9VKut14CnCH+Ac1t3qwo9tTMtZE5jp2opAJLND0V/ah7VdrZlHeERWLM
pzD2Y2pGsWP8F76I7AGyJh0rkyXVZbDdd4yP7sKOAW7vWkng/TY29Ni1VIaVGFe56Y2dwnL0ha9P
9KoEHOAMcfcnvBYPHQvpICNhsD3t0jfoOve7Co/4+kUJcvHP1pnMAZ1wgGz15Utu8TsR3mGI6beJ
E+Ji5E0vd7qbOW1JHG9ZCjl+RSb+ibQZ5VjlY6jaSedkb/I5Xkd/uTtdYMIvBxWypp0lpfV0fxHW
wkXAomeTeoTLUbCADER0dz4Se3SCUIHqfvd1APGq/Qqtg+SsQEwwBnQIImECppWgWxQLwteWz+kk
0stR0HBW2qgMtmCNUG8QT+lbhCiEHPEJanH3QZ0u4ntS4g6oFfcDl4z+zpMOCC+udM80cwfzadtT
YN3UttT7shIVnip1UOIR7aFgJBZrhH4aUZJ98Xk1s/ZLyT/pp8+S+AiRe8R2v9jFSVGpBA92x+tb
Qbj3UWFu4DvqXfuEzrZwrX5wy0ghilCAdpSRvYIWFFiMHbcNoY9lEACVTGsKFxBMkZgMWbRGU7gl
Y3l7x74yUUlh3s5OypvOtmK7jrcRYE71Sk8kK5WjplHlvUdfDoTP0STwTVs7djkUqagrUTOZucLU
0nVQF8UaDcN715/Z1r5F2wyh9R56XGNu6aR8IslgofJHrmjaGwoUkHtiPOuu7XpkrhOBQm/c0Q76
cInXf7dPuY+oKdzcff9bW2DLDBpP5rllrCWeaI7iyOMi9/+Q9vPz9GLsXCOHnYktAfZSpSQP6fbO
91Ns+ITgDcBFwV0dyqfxTuPCr3VBaDAqZq0MCFYynCfwUmLM8uWAgkHBF6d37DiTKlKdr/l29UMl
9gUEFOY0h56Tjc+Ij4tVDWAkhg/T5QQ2HzCGkvjH83iutF61E5ICPVvh1Tp1mRkivPak8QJWINU5
3zcfvI0+rLo8R0zC+v05aFcoqH52lMqWLLrWUefUQUgeLAmkllWTFAMo+OAcEHZN1jmWg1CjvyfW
vS55GehvkqPii+9/I5Zb0ZsNg+ZbxWrHUv9gwXt3RZNvuWGd+xwiEgFQBiPBMEwiyYv55qXrvpMu
Gh7MYdPWbK5mzc+ISJTZeCWDHIBv5QvBCJOYmPJ/V7m69UV1EHlIBBMODHVdyNMD8gQDEE8KheaK
eOYTwvKX0vNXxcu+AskoddKSTOEOL7HMFpGIXY6ekcPazSwk7/ogawzmHUSR5YlDkAoVxho52Qqe
kGF/WFRiVb1vIT14W6PvZDShbxIqMN/sTNAHirQw1PFyp0lMF1glSfB5qGoTFHwi1B82PEHtDWgF
1NvLmd88EQKOXzf9K158VwlCay3NousyiXDOkh+R2hgaNySbflEVsWPSVBmgWo+Et5GMl+LUAmwo
Q+CHoo3H1FtsIeGrpoA6EH9J+4hhc87XR3E/0JCT7u49ugTe1uUKI5ZZEY9YKtdCu4yd4ZOtl6JL
r08Ya9iVuDMJiltaGhyDBbDpveH5JueVNQ1r+jjW1lxy15VF5g+vHEoSI4YWxexHil1WtfpxKAq3
FYz7TuwOWhjh1WBAG37FVeS5EPXpq2aR7zWnj0oIsRIyj2mF3Z2FzdoBeZZZwtS3zgb2V6+6jnv3
dH00jtQQhpEpeRPeudujf/t4xmD+4FNFuxrQd+xwZ+YNqm2bEQRqYRxjwvSSR6Mq0GMZt68+JHhP
s5erGWXWHF+Bwv88kS8kHEhHlVXlpN8sXm9KTkE2AUFDl+uTWjKlTaiX1OiFCep3H6WEDJgxsHSO
jXCWXbllOCMa6VE3poMWvCtfxShihZcRg5C7p08DCVyI+thIi10jUuGzMGq3+9xj0Qy2apX53zfP
VV+IEfQWCPwx3e3OJBV8rr4jVNs+nPg6/2K5MvUtJmxrX9/dEhZIwerijw2pE6uZu/khQM2D3ESd
+74sbJiTJkv0RpFkaISmbnodYhIBlGHr33ldvMYdJQUFI/9ohLqCY49+0dCltsYrdVKYMTaaT/1m
fwwmqlkEugBpLWHH70dmI2h0OHbi/HWKjjK9DX+bqe7sUlRvt6UHR5kmOgbTra8zSbc12ragn5aI
JLFDSr5qyBwR3YLzfnpZQdwbAm6PRBs4wn/LZtGHgDsezaBujttkRhjhan3piEu7L1s/DXfwkXef
1XtqTuBE2Lwu2bXBnURbYr+390fu2jtG3XyumLvCQF4kBa8C7tdd7hkdFi7QbGTMJL9eAB2yOwsP
FDys66dc7AyaaexHLVmHxyALGXBkWNE9xLyxJflT7KemAENKDasuw5hkOcXlBzgpTmh7KVsiJmAq
K4yR6FFfEJ6HenjcV6AjKlru0R6x0029vA/rEos2ZrkIrdfanHZ6UKBkvOphUEHS2i1jqdIu2php
fcLgfuzibC29vUDARQNOYDT4MoqIOL+dUPlygyfVLy3/j7ZoREjKfmpU1NOd6eE+2/dU2HxiJDOa
eueJ5+w56eghNxxPysFlvyo9J1gECYhIfNDDtaCuP5peLYdQJtJmB7/RI1SLE9ki4xS6G5YlKHqo
fj4pLhiYzbjaU8pYfmPX/JZyiPTGgp8LpwSzX6sQn7Tyo7CvQB56XeY462NKXlFO/bYrQzZk6pU4
Ejb1SZphpKB41OF4ojy4/qTwNLut9VgBdhCvX3ERGJFogUXEmFH+eqlGsPquYUCKWp/rCMZIPWze
tFgV3ddQ4dY0mPp2mMYG4Ayl3e2qW8QeyZ+65x6rk+t/7NXzBFOhD1jvBZk8FergreIReGA4hPx2
ocKRylETTiHg6nGmBBACjDzzh6TwKCBHheJJG+jvI9aeFeK49ARcnodwkg/7nCNeWwlYiey0KPQ+
BdeCztWymbBaQs9YQlWuFFAWjXpduWskCCIgE5VR6pdelWp9I+lLRTNhG8OQA6pHkDNEl2Puts7z
3JjOOqFkzf1WU9kuIMPmTz+JktsJXXV2ynmarbKe3NrCKBgw55RGKJf6cxH251PRXltCzS5+CBAn
q+82a9BBbBIsvOvyoTGDBu4dmYaKNO13YYRP66zpvld/I0CE+ly7C1j8kDloMofqmibo1kr15s8Y
j6ys5SHSFk0UMK23GKY/tk8F8V2C8PcE64ZF0FdrNcMM1sevK3tDr3vEw1XxBUSZyuwDeyKaauk4
buqHWibtHR/U4PuQrnHBF7tdADT6wyCjIaPkpqmQCOekYsD8Z5/pSpg4uHMVIoEq93I2ljPvB7xn
LmYkik41SixA+oYGejxKK5QCZzIrHq0v/8WcORhiSmI8RuLDQF54KtilzN6wVxRBf/za+RjxtYnd
SjaWycAj588p1ZskD+YnIEDRSXuI8rrRKjXgwusvz320pLwnfF2xYvAmeBInUE/hylgLbl9dnuTH
9FT2sS+9WRnul4ONPWSjQuIL2bF5FeOV6dmELmYx7tdE41ac4TbSGeFdkbbGKDnfmHlNkRE4uN6S
Oydy5x9WnRXaSSorK2c9VnPjIzLKdfoKjq7MuHt1sEsX+BaNEQ3RcPi8PmCUaO1lcKQN+MOqMx0j
BiSxMLJYVXvueZ0GqYz8DdRPHuzb268HaMkItTCkcJfEo/GRO7Zdkah611EmyDOo5lP63GfnLwTu
tVVDrBkWlCFmmTt7yKvMoe/lIuPg7iygCLQXOI/b5OURTQ4fkD8HCNjnWvCigJd0GtAot84wTGKl
xwZPR8vJ5kd4Fy3SUh8MTr80u5PaMBJPrb6uHEWh5osauVp3jf6pCnsWZszQF/SPHqfacElsgxPn
gE7lKJ4TnZTSgXveCab7cM3H6t+JYoMfKvOKdmXYxQLn4axXweRrjoz2F32LmzhEk1uBzmDbiVYx
nomUsuF4r34YlVA7yB8FfcvyVhLmo/KEMQfB/kHhMTqjb7fTw2qZUkNv6saeBOWR4ByMDH0QSyp7
VWuOk39y+XXdv7kXFxQlvjMXbBVacTNCrfuc1/tRZ29l7PVwGHC8nKJLxv8/XIiJqVkL3s2ZwCx4
T6v5+vZa8BCSZ1Zy3SxIAzGq5AAmDyE7Q87ZE0WJzxfWJCz0imhoAg/BNTfYDffdrdtf7L2LBIoA
3P278y7WzNDz/CfcYO4VdLXp75X49vLC8fDiT6No8HLiCViCwgmGYXD7U0sG/BeaVhAA+BHHTm9h
0q8YLupEsp0XmvkFOVNID35M7n9ZMcRcvadX3ShDNYCvocZVejuakNPbN68mvAZOSWf+kB099O/R
SsYBWzSOuOcE+7qasp2jF5xw6IC6mynmxzlzkeXep5WmKu39/T7x60LW7snTVDt+7/Ncv3Fw5ENq
204x7BKQPOaMPwXMQX+JlsMNH5OiJpGBzaBDc748M0YFpA5LZUNhurFTeVZ9CDX2+UXRIuFTnNqk
IUVA23ci7UOIZJyII6b/nQbK6qSIIHV3yenUSnMt8urltmXZJul2EgwcXZ5K1kKauene6xMNejDE
Md2j2p6XiVBJKYU6vwLYxh6MfHVu7+bsY/ZPaUCs+bbPSiSruxy3p7sBD0eqz4Am1tbHauijkkSB
zTmVVOo7zMvedV5+ALXBdMCYJjSgaOKGo0HyxbHfpAU32GRTPiqo+BcS4daAfwtnYUz3zmoNrXmO
gUxjnHBpUrVWbVzpL09/b3CAbDPQ1uPyuateVRa8vbrBFxfATf28q5GvjqvlSrrqeF/egIR435ZG
R/r9RwxdTUeVqBwRwcFvtzpTwQSpPdHU5ih2y79mUF/M42t4Qw1rFik8e93gE007pD8qqUbmiMpe
ozhd6vRd/U8CWrJoplM3KARPEJBCA0D+o6hqpaQZEQ08x5J2NVeUG1PtGU3YKUu8hqYr8FwHMlu8
PSUCbuP/bafJIoP6fUuxMorn1ji8OQpgRdD7VqX0aRhVzVwALs8d5BKtsQlMos6oFPlve2nEHOqN
82uARqJHvD4atBOlU63VuFqZUxUox2KCBA+EMlGSWtKDRLNZ4jOFvEZzaPFTyMS6dhiBAZAmfGs0
FukQTBdtd8Lg2T02CZpUub74ny+Am/Iejy7l8xaxVpt+z12Va/lvGMKKXTs7BiR+CtZEGbg40RhT
pk1/6DYRMebKYPc/v7uFLIagpnA5SwPCnHRfaymVHZBPsMsLB+ebact/+lrkZFGDQKNCz3SQewVu
KjF9HJDaYEcfPL9V3I2APHqqEyuwFzshrKOptH/23cSdzvYlC9tgvA8s6ecgSLqWmH9waq5RUA+C
8NYp41GpIrBaRIm9lAX92DeBKqy5KZpLk8IP77XvpU2fBMb1CjkvmhF8Fs5YQdY2usK8Wu+WDVE+
aOuDBe8W57kewFV1SCJJiJxCanOaXWysywPzN/ZgH7xV2h9U8zFfSznoBe00g4fuMucGCphXCqWe
mjK5aM+czMjVR+hzJIBXb5uLwNs5zGdAaNHYvjtpVqJnqfpsygr0Qm/wUnmMTn4Ov/hxotjXKFU7
4t0KghRB6kn0twbi1w8QLGshofwV++dhAFJ3haqHVY8/tQejho9GWxAJJETeMFJPODs4/X3DCZCW
lQydC1c2qNoXNkPy8zAPchEPXIZ1wMJEC0eKTtMteNeBty169Jzxsat5MMmV2NSaXvu0qLMxs3it
l6P5GrOIRQTbmFfYXW3ApMPNh+yUrYFpP+rDoW9HI9zdyAygU3Bb5pR2pNtTkaPxM73hUJTt51es
u+fGm8tGUhEclpMus128eFiQP8ilStAmLcbF/Z8SYTXvw/y7bjux+WKUPAdFZRWmyTNzUmf2UJmY
QlF4vXxp3FSR6zKmhv2YWmzBBhOH7Iuxzx+QKdkaxiOUhOhp3kQK0myHJDb5UOJbNOQC9TXcuR0e
XPwV8p7aVN2ayagcKeLXqXclSkVEfC5u5jHVvhgC3yC4H26bAxVGG1MR7pKmcbsvoP2hoXC9opXc
q8/9JJ95Ntidz7xnI8gIZ52RXSZWonH/8YEbhE8wlNM+DP6daqGyPFrn8uEH4W9SnW0YmnXx0D6U
aV7QD6JeGvdJFyBqgkanczrtZZKAhpZF6MDNDSVCGI+ZxhgzwsSGK+QK6r9EyenMZHyIV5SqIheU
q+LbXkt5zqcYa3RwenDc3kznDVI+ucGC1v1XPiaS5JP1U6MHG5RUvDrd57Sn52R86RASTsFWuK0q
cWsB2kYOm+t91ae2HofY+jWbKxiBJ1jyMovkUt56cx5FLstbOPcL93ryknkKX7d9HnxGYsymUwVk
/ScWQdeUax+hAXuYohpga6iHiy9W6UWnJpzGbrgxMa+83JvrxK+o75gj9dmMk8kPA5o8M9kE+pQ8
24++2Lgx59coprqLWT70L7MZIrLppKmkK5IAXqt/jJQjyePNxEyHEXcclHF3ww8dfOzvBtsKv/XP
OVmr/7au15+crghUXHsiQLlAAmAxc+AhxI98daNv11EXoVVyL4y2a3yZOUkyAN6XdY2ShFY1qVVQ
v/Dmc5ZnACkO2OAlsJqVNQFXJyOQrMnMeJzyFhH8ky4czpWTNIscjV3zNI2LhIY7VR30HHX3wQH6
/QP2IL3XY5lcbzhyth2MKGk9kJmUYQWjMmgJu9cKsnH3/ibT8tSKKhvKLk3wCeVNMRUgcsZMoppD
TSBR6TPFK/RVLovkcCoIGNQMv9War6VYfx9MflDnvkTW3AM6ECBTnt5g8mVdYdmy/ErE28BsIuCZ
ps8u8s1hxXsL37ptkyo7KtmirLVvBUTpVcVr/t/8UBFQ0txL0sj/NXHXGZtY6b6aA9eC/HmvExnE
2QSioOqFMvMphiNQYJnD446lqWpP3CpK2d97TZpewT2IEYktB8kdjBvrN/KJ3di87ZqKc515caTT
32CXhJgr/dwAtEDd6Z4cf3/EEyLiWBRMkoX38MxBmrXxJgjVlSNQ2bErGbqdUdVzmJA/+P5ZS9Dt
9AvGZurC2Y1Wt+7maRLWhyzRcdQOiNuHXHJq9TYOIwoPjtNfW0wlKGpCRE5QJ7Psd3S+2x8DBlWb
tF5/uj2GybNY5kRv764jkkX+G1jcCdAjD9lQJMn2tw3XfNl1i6xfG7ezB2mWHF0lHmXqDU9Yg9NZ
C8WfKU71ptpb5ewpZVmGpunNZn4HUEtM375aWsp6Id1Cs79Dn/xuGSZWiylJSlPD5GcRHuoxS6X+
kLCfEY+c/eI2S4UNh5Lc4dh+hgOAvcp23PENSLE0VXAAOOHlmA9dT0W1Fjy++D3jMe8L1qcXmEQk
mXjERNVtwQFnQtexauTnskxV2GGTjTwlP4cPxLJLcjT9LNTvVHOBtlGhGw5vDZzOQTnSlQ7ck+DN
tw8IEmVFQj+YCJEtP4lYuL0fG+sTIJk5m0IZyM/kLI5ib7fbutosKe5Aw45OIF6TXbO+1hrIQl/3
hhE2o06BmDgLLE4W4efoJcHRU7Nv1aWK+LiKj/IjUcD+vAN5bvmOJvsUn3234QFFmXKOMJEi/H5A
dNh2qsTFbKb4PdOPM1qHCrmSyPOmey5pYbtHkcVEtvL5w6oTgu1SC5SbX6ys9tyiVEroj6SaAmaw
b/e7ELQB7ZHu7yRR/8fbZRzZSnzDwelH0QSkCRFMLOcv0HksYRai0v5Evi8QDPDaY/ZZo2wa6aIg
sw9bSqZAyaJshu1hJKn9iSNKUVTJ9DZBp/O/wB6XfKxvX9qW784uWl/GN0fP++8BDLvDFjb/o2Uk
YY3ifWGc3ICq6dUuCbajGDmPBkXYzU/VdtkgSFXTjMKbTDrlDqrPyMgzvPMrRZ36RzgaPaBD6NDt
ZvcxmIRAB2NulEdB+WtgVnVd2WLFNbe0ccWkDPPBlA+24W9E/zeK97EZrfBMnGT6GvwEvXzeDcGH
/aRwx9fHsLqrIXP4byj7G/8qAQeWyulhbJh/7SFNqZnbRSii/CvvSfSX69sivvN+eAfjSCU82NGg
ZF41VmVuWmeVd4QtXLbCn80nrTw7N2Lt0Gnu/nRkoGOGZhH1jSewn58UOheYSB2Seu9oXf4gR5XQ
Xw0RQuEhvrNGpE0hp3SVIFbkhlQIGyOSvu2zO3gDzFsbJKFnSXoZvUd5O3X+gQJ9QnVkYXTJbf9/
hZtuHX7aIb3prbN9PrRfpitf1a5/6FfDqPaFj8VsnaRD6ifn/KkiUP8Mvxv543Uac3nLHFizQGlK
Za9sSm6colxfxbLV6fvV9pQGil9keH/aFAcYWiTBA66Pc0pjU0qyJO8IfzAEe8w2HlwWctTcJRbt
wfv/eKEBnz4PV7kfy0Jg8Z33hM6mRTfcozwiXtN7m0xnYeKfLdFVL17A6UwJ/4zc2PPfUEgHJR/l
3SYpnQzccOjDqgaQ7zCqc3ircz7Y+GzFkkcexLZA9BzEVJYKJyiTBCK8bNoz2D/IH0ZWfXQdaCJ0
HXjVV7vk7FUrdJjs0J1KcFcnKXJL467ktNOaOsMB2qWmQFjgB9XrzTab1t69O+63axX6dLdBKtXr
wZfRpU3C4EA5zvrtsS6RlqGfSG/4nz5OHSZ0L/l2G13V2wPGPTcZLDj7nYXD/t9xVcrg27ZRRssq
8bJGuMwjlxP0O+RBUlZjrF2PsNYv1HHyX23l1GcbPsWVhyGx1tEm1E4grRAqFzebe/EFSM9PKqIH
WOIZFNnDpdqU9KEf46VVM41vrM6bD1OPiNkSPEddCFMz+l0taUp6giqy5fieFE84KsCmM3HLi4lx
XUeWztlok7/P0yzWvgGLu/fEbMUDFDJ5qsLrHdwi53STlWMn8OSy7yT0TGcr3JP6gUNYva0AWAPH
qRuPQaR60r4fXu7xOP/gUj66XZ8QBc4bRhFggYOLxGVWHLVq8YhZgIOFf+Jz88UhlpKC3hV1T1cL
98wx8DL4AtzVACXsgd+VZ9rs7aAHDHFhqVIIpUR+AMy80qxRJGtMd7nKoctNaWp2chIvBmU25mOk
d2DIaUSVwe5SYy6n0f3s6cGJmMj3y4KchA6Z/BTo3TlVPMEuzhlxPJwvdnTj4RG5+RnjiDyyNjdx
IfhKnGgUK8RCRNDK/T3m2AHR6YtT7p6c/XAcadzxI3LjuDDNOyFbHX0s/iJAkacXFWdfdfaVWNEV
weWePtY9Zh6DC//s/8O2UlsH8APMmjW6u1DlvalC6DAcLEIWy541bADyGKmVSvMIzgAn1cq2D8ds
AeGkg7GABRd1POzWVM92JuznzSNOyW2qiGvur9Ds6N4+MJUAOcrl3fReOed1L6m5kQVZSVn5H/yA
KR/F7ZuuzAO3rEkAGRPmhhzWvPVzywHaKAYTxdUkU3nVMg5gPSVfhyQKy1o6gj5QXw6x9R3kPvZ8
fPye4CcM7YQHdK66ZYsAnrizV52Lfjyq0oRgumo/61oPYo4AlBvQmR4hMFu5Tzlb9peTaENMpUvB
Hlec3fwV0Of2OTiGbaQM6mdOy2K7GpmCsUpkHgWqPLtIvMGgXdCVfCJwIyNpijx5s/ZYUcABhEaU
mBHgctXKz8t1ZPdwpAG5AscSLptyhGzA8nC0mOuqHBe+hx0jA6ArRRHBthKS31CESsc4J9EgmsfC
MB8x7Q5qdFoyHfEfy9DDbffCtPbfIXTYl6rdC4MsaKrh4JpBoEXiPNRyDnkB9W12h0JjhKv409m2
lCZFJlNhZoEFljD/EDeECjx1wSYFx8vDTstfvL/vMtVzaNlE4+lIzKW1RFjgfn3AfAj0eNumpV2P
I4aLPCsOy10lnBX92A+cRU/W1l7MzoQnvVpru4IedETzle8i6fArOrO9oAvqf16En4FXg/RlL44d
zR9FmuEBmx+DN/1ttVxtNTc3Ptz/kU+X8ofRrCH/DrcQqv9UIkh0wFSgpM3GOxBzpeGAg4+gEEjb
fAQNaZOZc6ibQa10NiNB3s5zE935NsXLzGVNRlAuHUMILMjZ2M7L04Rc6z8GW9tDw/YoNfCLZw+Q
xbeljAEfNeAGLyk9rxHal1rYUM/xSm/Ws5fKIWJVbDMtxzXeJiCd4izRqBevuTdNVY4j5kSedA8O
Mi+ZPhP427wHWtte4MvvKF/eekTpyVX+MfLMW/MvcP56IqrIgBpM1YcfSSyHUHCUsKy+VoNXmK3Z
ioHB3otwm5OiA7Q3GiciH/qZLmk1rTYkz1Q3wtqjCB/PyAQg95FD0AowjVZ/rwh5CWTpAGdDblF3
A/wc/SbRBbC741z0G0XVpl2gzAP2BK2MnGd3844ws40TTUx1Gh9SMrvBlTZ0T+cNaL4yjURgOmtJ
jTt9P35bfEID7NAZtHG/n+XQaweZHYP9DY/AIirxhrtMv+Tu5SCXKvo95DqZt/shY0phhwtyLqni
jrbK0AJmzXQQbGTIWS5cXAZRrI/go4cK5rYGWKWIJhw1iVlYFb743q8OJ5uDuNHRKHnUS9Iix9Qb
f/5qkz0z9ofaEp+7Q31DCwZdxSAVkF7icZU3ceR54Z+8AOF0Q6zRyEaMb2YCK47Dbuw+DiXNZe75
LAwAh3C4KK5dD9kYAF8PETehyka3czInZ5mCy0C+NDTF28AhpaU3usX7G/GQ0+XFqFBzngGXVuv/
xpVdyAdF4Up6dRnSRrBIC/rGQnN+zkNAABtsf19M6SosQjJWiDwLBBFf/kLa+VQO48pictRzukD1
NbViDQ8qKmL6M/ri/D9/QAO0UZ82CTZsslBY2gggbt/PRzkG0X5tvhb7tPLZmYI07FFWIaIVb6yx
djBACZbQ3NXc8aaDpfELJSlLMQKUhYP2LAobWwP4XhHQoZTY68Qu8AdznalXnrMfU5cSjgjkYB2r
y5WNUlMePIySjIGJl+EqHErOkD2YLrHU+sl7okBeILmXCZn3Liuc/6fTYsGsx9e8RCOOxJ0cvCet
8gWVXwOT6mEEwenCD5QcdxPQzjbRJBiEk5L36uGv2rwJtFexbxDx+w8j0OQwZV177yvU8c7PtMig
hgP9c67OKCIqC87AsH9Jll96qeNgPe0EJVfWlqXtXbw2kV/KwnvW3NB1fzzmuLjfBFR0FG5xx4Ec
MbOOscDrvNEXxPVbpf4UOoVetTtSG4eCr1YqY+kInaoyhdJBVZXsbOxKill2vHbWfqfPaeyjei9V
RhlQlONc+c6lZwog0HiWweWgQTKkdAcuzHQk5SuL/k74eE+Lyw72Q2ahAigv2AF2eXyh6E5Bt++Q
01XAHbULvsnhyyKC/R6D8B9QwFPGMd3oZTEKhl3t2LiL7lJwN8uXMBZIZC3pfBIW9atHxPyS1y9h
qKWUv+wpmZ+7OWKwNEbWDgit73h2mKIhaUVQFTCjlhy1ESH3PJse8VMOusvVV5JsOIrwDSnQS1AH
BTR3KRXvOpVHmD4ygOEV4q/kxD18vA3MrH3OnQDQbXUU64ixr95CMIRotwnYi7Er91qVX4RNiUzs
6ltT0jp6mpNZ+XT00tGsGO/FENclR/CcFkD026NcERoHwhreQtHvwrvRdgYc+vNlRt5Xv19oTTfL
IEGtrc9HaCtzTbeJMQEtrThrUqwnmX4crEQ9KUJsR0flftzXA8TfC4RwbMDM0KjFBRZdOPhKPzx3
9WFNWQ9BlDJBtkG1lp0CDshPZ1lYsnT1uiP/pHf+VsaiI1hIluqChJo7IupUgcsVOsM1U5clvE8s
pLshA4KZj1WW+nvk5geDgjYyx7s2YYR+bWvGYhu1Pmihw5/LiiLih1Xm9dSjR3hW04VIpN6sYy32
a8XXDnIhC5PDks5bSCTm0jolrkiOIjTTHNyuqgD9hLQmq5QzvaJig0K2dC7HJ7qpmPq8MCkrgs8q
1jKVWaHmSvHJ//8s/eABCcsgcXmLOHFzfl8993jhB77IlMgeuQwJerSMQJlKVKalpVnE4TSz+/1D
54ZPg+E5NGxET5kHoRNvM9aMB127CGD00M3Dm5JFkXCC0MXDuBtgFGPsQi7FMMqDWy+7cvTnN9yB
HHWLuJWm/eHfBt/Yk+st59CV1ce87pMPk1kLM9vErXFZLaYUBSEQVPROq8Fp3SGB5M3oHcJruEkF
7vNWBdEop3ZneFx4SUzysoVoTq+iJ+VVKBDzwpQGp/NQRDamXPwh+yypAgEGJOkdhsjd/5SFOV3t
CipJuDR+jkd98ggIr8fFXDrWD1KgQdB9cG2Idd8DYii3yHPQGBSVSeQdr392D8Q9llkOEVtJ3ZfG
50ixz18D51x3iWiSW0UfqH0RUEsw7bwvf/gDNmHopCMrvjL2hAaL3HkTmC9PALE/3jZUgz13vz5z
YmfutgimVZnfrOiu7UP2OdBKle2iE2yYdXW54+7cLdnXbLw2qUjXntiQHlk7/WjD+3Hs7/y33GYx
cZPhchylWvVnTFVsbXWV9401E0LIhzzwi20Ohe9+Q6iKqLrcX2F9X1u+Y/4LiKzhmaes/Qf4ccLb
QTwsoj3RI9wyA9anquKUZsWr4UPp1Z7v8Gd7TrnFpt1JtCmHgfRMINyyHejQZtZFcdzNDht8mQfz
3q6qkalYxsfmH7+qP6rVtE87f81xb1ri4je3yQGcLJOdvJm5b9KGetsRpmotRCJWZYF7uLGHcxA5
lKONMLoqWgcBPQpOURU+RT5wakeDZthF6i+3EMcItrpDPLMDQyfc208QrPPAQ4NlfaHjWP+9jK/4
q1fbpCSPuhgm+YrXv/fWNZrN+P1YGf4UIppTtt94YaEPW3bkTCOpxxekfUyoWmFnR4Gzlusr6T93
BwYHcmjPiYLtbZFZflyn4OmffLWNfTJhighqPTtk/lYyYPgZxkRzYKmK2HdJ2x4wmMk++KsaSQo3
fVhQU6HQyIMTLUjQpjco9bXRbQCgcAnXtf52n1hRCpAIaEFa5h26nEXqCqe8TfCuskZmkJIF6C16
AvX12NkTJ0Irwcz0yEap6t1VCLYBPVOIfgb5mBfkAyW7j7uaq2Nz7ssWeP2lpBcDWCQfHftt6kwT
L2dy4VBuogmh3rjxp7z9AbbiDZ+Yfro36Kxsr7dlzVLywtS2bsJqMinGUr4O4iComrBp9HDoLEzY
lI8gBuFHb335hJI/QOEOvaHF+9slK58lliD/ha93sTSa9ix/pSMytNaGfgypak4DfAA4395WPVjn
5tuhOWafhj2G55+ZfgbTeoxEh1L2Hz0nKnJaHEAKIodzH2tueSc4kgUFy6HVYaXzK9bw5HsbVMiB
RsF1e4nQpHBOXR1QJvha9MMoANUwvyRoHHrof+nuRke5uGMcImjldpHPMV3iQxbdxletiF/VOrjf
QgocxTkQ9opxoPCVL3JDLyLyouOdVfwIlrHLCLWcLq1BqmkA/biv/FgflKliUKCTdV/WXNpTv3GW
2J0m9FDPkgBOlJuZqQoS04AK0otHLO+vJCQBVSMm76SbDlkvFbvju+/X0eD5bS8X389jktebk7fO
CRZTvZKqDaFZVAa1JFwU0UTn2UPwDiTc1nn/c0MxXYAtvi0Riql/B+JI9djrmdFsUwZWOp2RQxD/
zw+JOkA/rqLt2dcdY1tblYuMI9t80s9grtYrMuSKXVUidQS72Z3+cfiZxTWNE2biBtKkZgQLOwBw
phkOFX9g0s2m3t/RHw+KGeRhYC8O7bfOUnvqOQdbwW0VP9nMDY6XPmB4tOVxe5frZnr7y4cVdweX
b0yQ1UcBp6zvgN7Yu8Hi6PnTTR2uBty0rZCe9VbRrBOv5skcCuoSg7TdeDv4u9tx2fmCti9jr2Fj
BUIZelB6bd/XMVqoiuH5wOxUH6E0JLW/XShelG/TpXkZ0lYgAcYNM5z17XPx8PGii5ZV2EGzZtY7
9gyl3h0laet99sGjvSq5NnUIIWs3pMK9iXPz6IgDFEo2P6iujHsu+39esQODpOIAqMwM6FsfS8A0
uHXK4o6HVuMeV9qBNZWocm9s2frNnsAiVh/YqzEWIn2ShszAwuzyrdzjratXuOkivS+nWvKXhD0P
/P19+UpdPWtqOfYrvmOGwCwPAtII1L0I9fSEEsm0xkdJ1hpPFc4tjMgUVxxKqpdWf+RPkMyBkyzt
htOC5mOyFYT6CbEtfX2LRsNN2LHAYtlHUGyc7SsJ1i12mWdzbI/vZJZCnXBK8pIE0h9ECfTKrr+P
nh4C+RGui53nnj+mVqH3JnoMW0RzvnaGIcgvFRoKCMt10f3pPDFtkRn2/ndYU1NPG3wg/i3AzZxx
uGbxHmPbt4yhSc/Ubh+pPWU2RKF/lQ7S8QPZ/y6IQpiWYfaU2t5iR0DHuqv7+S76zG0u3+QGP1hD
0UvVpb7JC/fZZmGBr3ypENAdO3GpQUVxbw8WD6YCQnJtKWGICszIkI9BwV9gdWEPHCqeTpI+Tpol
ifOxEd9f/OvBcNK42Oay2E2dsIbQpXLjKaxlffGI8zothsplirEMl3EZ1sd8FdpybYet57pGbyna
UTt1KpZsMM7T+dOlLzyHT+hvkdFG2Ht4eTUA4pXEZDZ+Cx5jBurdmPssxNm9dYTcJ/86SdixFzCg
vWMufP4bL6NrVCZ+JkKQpD1d+NGQXHPI4pCO3n1Tuk/lCLIrjjg4Zki/tSu2Kg+esZRiDg4lh/Z/
6DO4zK1fxcmNxrIh83GMs7rE5a5tiiH54ILCyJjFaWWsTy7uSiWE/1bCEIMZ1Ve+nyAqUCkRzqZ/
jIwxGiIeTjUJctbG4+77RhyWjuqe4v8HQoBsShcbd42M6efauAMr5f0ZdlgPs/t2OhxlyazYvqo5
vVjl2qQcJjKgOWnZqLrcj7MAnQwo3vvyJhl1s++cKAdutwhzhkai/TuviRvuxyWGwj/5lCkrLs15
yblMV3N7uRsumQAOqb/lHYmYkV26NTpnGNwD5uJs9tzSQWBkhZx5nqmrkSW7WprQDqpPGmJvs1ZR
bo06j1OUJJms5MM/V6p8+XzApYCIFFTI3Y4Dl2DjoLUhPPFeGBOcEHNyKPVyU64VUfVQJsdTTGei
CH4r9rbq1vuPHXkDnfXkaFPrJzI/x1eEfn3f5Y7NpsNTxpMFLoyb61SC+JCcnvSnmuzw90aF+5N+
R1MqMphN+8oHNrsP768jySZqMHrcs8erkoVsnGhdx0fvljw/XOHGXBztxMV4utntcig2FXzjKAq+
jABAGgAWRwaQwtR5BFKy9QyCs3tN/7t8C9HmOG3nySVA8nXG7/uj8Tbnpc1T5+jnMgNSwddMHDmA
Bm95+ZnDbwuwCWqhvXtr48o7dIzTuLalgFTg4kzUm2QK5EcR+VuSC16fAeeQzMjqXzjAgH7ZoOwt
JUNCoODUUx3Qvh7Sd5ENouxkdfeZctm8G4DcSaB6Z3m4JmogwelRL7/wIduLFflI1sF3P3x1SU6t
JVaqvBDsCWtfPdnUE394nTMyPCAMXh+VbH/RttZne8YM+69QlqiWWnkPxZRDjxq0MWTgR8lF2dQ0
9gurY2b5gkBljTLeDOeQfXoyERobLpT4Ae3wCgNgHjnugKZgGnvMX4pvy62Sc1wTyea35m5wYadw
JjRvtNzQxnK1tiMvOvoUeawiMnlVjg7WSGfeZWpzEPUFGGmsDCNQJUXzlOKYXwd8EzdzrvlHfbBJ
bbu43tG9xcpf2mvZwXXL4+vEhvfXjNqgyEjyj9xeCNXPac7fOwemDV6gQofRGa/4dkqqQBmBekds
KL/HdH4fudRfsaV6w9SoW9BxpoUwGsXjsnt4z75AaICmdPIxJGb9yzC7PhJJNmVh/7uzewkQ6a26
hMPq6NVzb9IBfHYZlKy5p2g7Rfp2uezOGyvQ8rRTgVQReXtGJQKU5n6xAuQa7sbIewQlCL+Nljxn
jmmqcdgssYa4vGJv/OXc+F1GNIEqReNjiNFHLXQVt2oZ0Gw4rDdGMy0T4Ve0NEqvw6rDcW3lmpsT
T3ekNHCSQcc34F9OEkZks/wUM0nx0plx4RLBX367y9yTJPeMI+bHtOUys2uEsBUCOLT5v4OfQNVi
ccFZDZIPXVFnf/jXSdNd2ypRHiN1J6HBgUmbg/JybCAz578/Zut4FCPPY/QUWST/cBo72WJeGQ0Y
S3RuO2xsUT47O2PTSHYZrNZWH+g3hBnE9mp0mujoRumBgIGPQY0yIg+AM9U10QNUo+DzfwdTNHO1
UhMGunG252fSDtifOT0xtQ+Ig1HecxzGjeyAE6pisrVk0tB/w7pND9LuR/NWe9HJLtBpM/p0jVAY
23IIWAmSuOBmGj/ySusl7fekWpjXFq6AT+WilVtIKGRLPSwkJnga5AHaEn0kx6aJP7+rYAuMw/03
XJWYQ9UwZSEzthhBUaVNJpCwFg/iKfNNQsDStPFPcp2kSVBD1/cush5ykc6BzmqH+N8PV+8qdZ6U
U+m+sKP/SSXifhNfnQlr/wM0rV0/98CDvbGvvXhy2xGqNmGsveiH+Oc0wGipTZPmY8rQmv3XsLzw
TXZSzeaC5whLa2A9asEClu3ItxZS+W9bPwd3QAvu+d4KvFTpTByhZVNCE0x191MpavLTLKl/aHY5
GgWD3TZsibZ++wqhOgVMh4M6sIL+1k9ROSrLGgozCK4CDbkWNrrF28Sycg7RtS9u1Ljv2iNXra6m
Fvr/VjVl/SoGUsjsVj1ZWy+6hdantSxoLuvQtvfJJsEEfGv1Hl0r4zGkeIYCMCnKhhPVXyb+OWC6
QtEtHt9QYrLv3iyt2YVHEyQzzvM8duPy4vLg1zf0RO6CrnEYPJAVtkj7GKKbYASU6Z6raquHvPYi
QY8aQVOf60qURgH33Fr9aGD1nCI8kp90n6yudStZVYLLdzTnIP/1PetDBIPlSDyGh/GvOg96yjAQ
yjJ+KsmU/MjmKtXLIfx75hOT2laq0x2q6tpgH0shtU5g74wlOU416bG9d65NqEBVPLQW9Fsh36Ig
rmfWUO1I0uPwMwjt2987ZAAWeUh8sNQfqWtUWc67f5v4qoaPUf0/3Dl43Y6KAl1Cl5t2WlWQfxxN
I6NXADsETSI97oNKMcpErJojFqVMP4unTGj3Zedrh3hIuej1atrF/W7e4z7DiiD+fEyJpTVnLpST
MW5Nh1oAo/rIN7+GmCvEGTTw/LG5Z3IjDutGeaB+2belEwGuwesxY/W1yzogJPLJVcLppB4PSGTH
qiNtskm0NI1PmmKozqqhQhZevMuUCwztfmqoX4xXauvx0i8QLGxWEHUqTp/e4Uc5PFMsUtoYxroC
tnZVf5M53DlEb3CmF9uVYDKIDnosH3UmPfi++25ek1bTatg5Nrd6VLu/HrY1BjQfUbIjjY/wKU90
68G8OWfdl7ZPrbIsLc/hkeEs2kMl5j2nRyitm99ckQoRpjf2z21YqIl76FuR9vGfaO9xWaAVcHDb
WQIDRMVyPK3zxWc38MGzhLPjkRWP3DnTG4ryBbpOGCSWHkfXf9Str2E/epk95wuuFfHqWkZneKhS
7t5dDMIFNwGlqdoPN0g4RRz6q5TpnM13Vkd7RzBr9X1GigKelztnqEQf0vxEGkYa56DqKV6d1+o6
Qz80GVMfKOo8/0ehJ+unMMsDKd5V6uLBD9J7T6v5ej5+JTItv9SzacPrg5lql33lWQh0Ezf3+ifj
a9ug7aORaVZJlTakoWtsN5xvns+FwZuGDzlWgZefQUUBICs5KxsxrVFfdKyt8ZrrvnvGUGxY4+W9
BTEhZepkDaxn8/g9uLb/ewwOPnIH9KKWWdfi1tryrcT+qwNDTMKTzzoqp6u5ttKaKNTw7nSA64pL
11wMnMfkseWY6QuDCU/gxpp9LWya5KmnWqjXS6u3kzm2BO6HWk2xNHaD/PnJAZqWyB3mW4IEDfd8
XgEGMBbZ13EmufN1AMzFDaHz8Z6J+aWvWeVD2tcURV9KxtHALPOVReHG927w6Cd0hKvny84U31Ws
F2TtBjDv5RnRQ/aTwosjGMFcwnuKZCTHruXFFLRC4yIE85qgA6CvfJWCIa7MUcd/Kna13Z3IaFTo
z2rJCkft5zCzrYXcKHzsXbBvsNTnnMNdNtsakMnycBIW/hriU2/ezeoBs50k7W33gfaEXiv3t+EV
wCyARhynYyutLu2uQMkPqkmcBkQD2M5S6ZKa3EIj4uYbmmH6Ltjqvrv1bThmPS7dY1qZw2vGBrCS
61B35yaHDQ2k/5XIoGlahr462Gbtao17mbz3n9dtoc3O1f5a09VZYoOA9110WCXJUSd6N5WYuLiv
uQg2s2k1VGhY5P1ix9CYLeAGWN1285+rfQX94MTLXfXEFmqBam7Abl3sTz1wcHn/QdXAsda9g6fI
yLqXXFu38PLrDPLLnYeuSfbbMF3MMGaBFSvLCkDmVgfSnWidgR0bcgpZeJvR/8RdV1XYPAWFTik1
dJRgMlc+v+zQBVV7d56/Vtg7gyJuXGOrgWhnk2YpvaS2l0MzW6s1R+dpwDKMe6NE1H8U+m2FpN/n
0CbhmW/ysclSrsBQ7hbyTtr/2elAQxo/yT4eWeFRaBL/vVzYLXJEDewTsPORVQQNzub7EF9HGNcb
gR+pTHFHrWCTNH5ggdTup62gL+Q5QVXn83XyWEnLh0fw6Vaeh5ANYenpU7SQDOR80OIzzemJHfOz
2qYnuzGtFzFJZ6LyATpDbbeqa8Ai0r85O2P0vnYP6ic/TAwLX25Ainy3CVuyK/w5uoRz1XgIpsic
dsbOW6D5qZem4a5df+9aTmREYIv3ynXRrLglsvL29UtJAyEzFHisvg7DEaqRS1nbRlncet6XdCre
aC9Jb5u/nFZsJXq2zwnOh3ts0ds2nYWTFwcYb9pK5lFhEwkgy95CKABCZn7qy163jn/TBZ1o/bEE
GoG06LnkEhRSeJk4/UOdq7fjStf+9/GVm4Ugq2OR+veE7Ut3gcaY3LpaYmJ+epl9g3cw8tPfqOI0
Qah3VGtV8EXqcbiI1f0H7gRDPcDt2tLcLIJo/GhBWiDk/bXbQ148ZM4jbthCj5pFr/h0iMDrdybh
FQhdyqiHUx91a5QXmk2tcBNZ9N49R2NoVLx6vSBNsmnQNquVL5fmSanfz3e/e6VvP87kIdIbprJh
4kwZ1l9eSmDT9YFA0x9gmINT+XhEuWBdOJX1C0olllEhrHip0qNlB4aWNt0krOUpfgNVP2OZaQ5t
SpDzDwArJyEQNrtNGyJmlZmXVESSf5W+mkF2McJlcjpQz5M3xjEOZVlv4JYhlX0VWmgKTKj5CotZ
AMLTWmrbcbkpmeLVB34NWNEeShlQqrFrVrD4yxSe5esmk5MbKAegHE2hIIb4uom9y7B5ncBdkxXr
+WF/1u6T38eLmpbhSaoIUr1CNUZyEE9kPG6GnVMRwg66+65myf/237t0dGmznNBfkjR5GlH31PwV
DAmYDVODb/oL1jwy+nmZOsJzSp0WVmo8sjrE2PZ6r/MFpnByR7Hi0xhC0a8pfbcR3eKwt3YXkxrC
992u8/KYR7+/ct925pWUSiPvcyl4mPUgyjss2FwPZ2e8l3C7H8p/i0HCKIUq5kEA9gV7i8zvvQsS
vYXp6vhT77f3OalnDWJPOoXc2UyD59Tk91lvKaL9l55OCm+DsqJ0OzWEjUKKlqhG3hMcL0LOIsNk
kqHDUrE89u8j7EL3mI10l3V8HVwnYIy/F3Oh5/t5GjJBIoJ77hjoT60enyjWSZrt1jARMQ0EgFLX
6ojLGFoVPRyBQrZbxkHQO5FMkegfcL3cC6BEkYsw9xN/sBtBSeX76G2HItWrMxe3LoOOcaBfLvR4
KWcJFGs4Si/0Qk3JUTTXQ+18TKSmhcm7+CaWU6dtoC29aS4TBZZZcgipmajZF1ViNk66drs8ejsF
SkQiScB1X+L8AYtOpZtcygyqT5biDgb+7QUEKjdRKRBZ+BatiOgW/iTmPuRET7oTE1gNrelZZx5b
EZR26vyUXTeJvcEiCLy+vhcm8+t5D+7XqcCJyLDAsgGmPHv5PPIiD18R0uxhDMb+WyMoidIvLb6L
N36mgmG4sII3G3PC6AKp03xBlqZfh3k7RFHzBJaAFNwmZK6mzM4FGVLzYY2hBbvILNPGsSbgRnlK
vEG2cQXLkkibrRCdWswsUevBVryGs0jEUyTxRWhgUi3X3OQ/njnWsVSRodqkceq/eXanUAsFGD9s
GPBCaUOVQPB5d+EIwQwTApxGPoE2sM2dpKXwAW8DE+fDnzzM5gneq9PyZ7T11Zhdzea2V4un98lS
yw0NvZAznVhDiZFVFlSYAiS4AN1HGYd/6Kxhk9YWTndYkhsNFln1+AmCqUdJb72dOSeXoH8pxaO+
RYtmiWb73GWzWbgAnzpHo+HoXxvW1d6+haW4nUJ/sntGoW1PyalG7lP1HDJY4L1W4gwi40Z0duOJ
IKMyy8UEe/hOg1LTQpak9UTwHtVl+tdtNhEOeTeuq6R23mtC8JvHIWG9nvZ9xYvEprXztyGJU8tc
30GtIN2bkr+3x9COcpw1h8TZvwSqMpZq+gu4PyT65Gqzc1aEmZzGRfGFCMk0VazPkPGoVqDzdBC5
nTfEIZ57+K4encpO7qx3HYnUTTXL4q5k7fCj39D1jsYgN6To+DfMTBTtRcHpMz9xX/WfDiDTkkFX
g5fkGF9pc2WAvK7Rjx0HNt9Qwl3c2v9+b/Cor9Qleqe9kKXPEA2HwWPVkhVMiVfY0I3YYYmYdt3G
GZJSrkhB6ZIgnKKS9ZDXeFU4x4y3x1rWgFnmV7r6UcH9QsyKTGXt84dR0W2lW08U7FZWa5Xhoaex
0q7xVUW28fkO40OPwMA5pmKBYKBH1BAMBT/k1g3UvOvGCmnlSqotLeBdFk9hPeYWOzjoSWb4WthH
p9p6CaEZ5hbxLDe0Q8Lbbz/HDgmrf54eodjEIbx21gudJEHsjt83xcCbQslmZe86lRT+8fZMO5Ru
mn2xE1Rxy7gSABT62uOZrkWCnqSZHONaCiWcPukoBeMYr/W9wXIY26UF94t5TiQ8huGggPMdzd6h
teXrcVH5Fuk/iN8M6/oqHBYZbMztn0qlEHyQblHAHrI/WfV8YoUaNL8USs2EhFJrEFS6QpDY9q8L
f2I7qBylnyhlqyDB/O6pXkLOo1t8sF0MFFH4x4uJ95GsGzSYbRZ9+u859+aE/wAJXQpdggkqg8ih
s56Uyen11oaqipbr4iUMO+Rk6+IjpwMho0tQDyxCWQFZIu85LbNgwYdAEBMfpWgSWrQEH9/p9W0P
IiyXW9Rl9mwWd8nYV5lkKzptCoMEkjEavvUP2kJQY7WLYAsmqi1ZV4wHvaxzRqMvVv/8UFbhVesB
BlSHQfBLEqEAjt4buz7T4NPcds7rKpJbCcR8neHvSVXVT/uPLoT+Ogk7wHGJWJ+dGrHwUjxIDJxK
LWz4Pi/LfjyRiikb7W9JL818MbnX5FzsnJs/q1YkH6v+xyCAf7FqXxTe6R1xLzp3qRk/ruS0vGCA
vTSvL7e7V6Jqx1QbFwytdl1wXfZBb2NkjWphrmbJTmGEY9U2mh3HGwtCv0pH0ZMPTtHkiqg4BX+8
T+XrqOe1HcX+YUVPDhUXI22LQ7qPlDHliZqCYxFT8NcZGoOPTbdCe6pU/WDyXuqYW9Nl3fMWkX/Q
ViwpwyrlGxHstYyhDcgE6oNrlErlYfmwZzzH7bjLRKDJM16oRSyjMSYel6m18DKxRp6MWIkGvnan
1qBx/+6CKdl575ubZxGAYKEc+29qjbKjGcjnLovpjrVjgIBfsTM56AiqSgN+xxCH4HOnCKLx/yHo
oVwAu0nXOYjG5aiR2joHM2svu5UApWnUm/C6JaG9HLPt3wzYnr5+qYbd7CwKNIKhXwBRL80l6I9g
BS9ZzpxaKtGl7Fygq43SLY+7OUkr7XpOI4IMDHuT7Oq9g/XEO2iVpZIrFKodlb2F3WzrUoBflLYM
b747FXjr92wlV4HG0KTA00kVRvazliYz2+yhSamtD+igi66OiWu0Wkt4tlja3E3cBKnmsqnMxtlj
QiU5cqGnioD7g7FQ4nyYxiJPnFqvoMoQ1d83//4Tt8P9bFRG3lrHcrND9wVKhbtpuW9GTxrT6YKb
CTtuhyRUgLhMswVnSihXUvzpm3tOx00eJ05pUdGOBDWhmTMatLO5YlH4z770jZn70kZ+Hs+G0ujK
8GU4wunLGgED1iiA/2uyDrbQTqBeJ25KSFIGuC29Mem6DjAhHZoA+mtA5OsHxQQzcUECidMUYNaP
A81bP0EnndW8fSBR1RXsgWbqkllL4sLKKB88PKr7VqxDTUtgyE7DVpQM5BMvI12jRVMzDChijBiz
X9pDI0ntjkkIeOhC+vW8E60VLn0pvgOZ0TpO37lP2/lfY4QZyHeRs+1wLUojIBIyWvJHHbiqaw+1
t34bNRa1PbmG4kLluHmJgEcG03pNSN46QKaguYINpSxc5MMH4mjKUlbyoOl4Qlqo1vkWHIFVgU0U
I8AC4+iwKCS9Z0f4SuTa79anYJq8BbyHTPlJ63N6VCMRKkBIN8osC8htOicNwFTXMVnCwnrZSo/A
5SHrzGszavhS+6eJHl7YHUVNBPLRRrn7hHUc8iV+QZjGrDvH51VJdUKgVqG3XsFxI0imNwj/Iamc
cOTlYmiJ4Jy5vTZXRgt3N3xTfUpnBpjw8VemljGJro6BMrLoxoIpb7qkApmy3lXfgzyldpiTjmWy
5W9E8e5i//AbWspB8guOTS4KPkLBqOIisQOL0kpra8AaY0i9CdZV+C0QdJnwgZI4wHUXzHiGkpb/
JEQQU6DCcCfoTWXBHiesOXeNSl7VkeVylNhb7PHLwdbcoma8lllLME/ALJjv5fnO3P77egEus7P2
z1O/D1XBwrEk+ZnjsaC9qGQE4GZwoxvztgWEdVhmuW9Xnjb4feyXcVTf032lec2qljvBKjyjLWWp
BKj/zMFP9brLWigUuRV8DmFfzBq1tj79znTYOMjqohUznUCyT8YqTIyBGyDY/jPWmUVNpDBVQNi0
E1/ReWaJMS2N0S76N5NK/5PxNQLX30IeZZKoR0cFqNsaEItCdEaZYVcqF8WojLY/ILxaa5Mtx2c3
jFwagahA/Mq8X6aYELVgJE/8KZaPTwGL4pfYGRgMhyhYNdi9r3JitmBiAV1YzBjVghoxX5VSlklN
Pj6HKaTyfMp7SCWbhscbRBA9cMd1GJpr2hKn2hZy7hhAkOQzvX4rjNEew5o0tEXMxjO3vrolHuKk
8NpwZUW3IzzxhO2MZLj1si6h068v29EvCZUQ4esmY9JsKbtkdH1Hg432JisDbphor/Xq+e+yQ62f
Ud7PYh7H9GOf6AXxeSYu9xfpItbJ6VxqBcCkoBjgZnPv+dU9Qjr0ZQXdJvr5QsWo6uAiWs41I+9+
3TW4FKMvJYEiPEN7LwmZh05x5uFxsSWfGMCCL0jyA/o9o3zokkoy051VcykoXwdLnFc5L4jpc/l7
3g2t3UVGL0WfoiniROV3shOwlaC0QilFFFfcrg+bLLCzyWVMBkV3cGkab9ufQzI2aI8l1EXetzAj
48gr7eRqQt2dlCMG2BfgMoO8ku+bEaw79wVPUVJTjB4ApZA1P/khmMOB1CzzFEPtoPXH/lSO+So9
W1QDow22LMmCBf3XNb/jxN80qeaBR4BI7p3vc1biRO7xmCVy1R/5qnXX5vamvMrGtW1CkMa22zx/
40OraA7Ovof/mFq8+lKw7aQ6ez8FzUp0CystUbD/XSpA5B4ZWbJnfwj9FuoXYPZs5K+mjpS0yXv3
vGNP9/EzuoptZNIPtecWhNIo96mXq+ZaUS+mTO7QbfFfk8Bv+WWbHXllOKg1Knc40w2uok7ENgnd
sNsp60zeeFrzXA9SHVqxQJRGUSqwQGksWXT63bGCrerajuBKvx4dYoZENP0JdA4fQsUOZvzmsJ9A
NG1fo/4hYpew355f7r5stKHgDePx7CnXfrvg1RDBq6BZi3nfWCGi732MoPFHr1qIf6eFz8xLe0h4
kAMdzV/0RE/r2G5lEePJJ1UdqPN0azSDQ6ro9SRf9EahAJmwS0sAk35YOmpVTy7np1xDQHcvIJN9
fX9TJUkJat56G1NmrPbvYicfnCvviiKi8jc9f2ELMbbhKyL4R+DWYe1yBY37vcrx1QT+ui60lEqY
pW74fbbxY8od5GGpeVM2TVnQs5I33lbO53VS0rwcq/HFjYKY/X9y3ID7R2BZt/xJzQllg4H6hboW
/z6B4C1qyWQEWrNtjIaSJyDIiInq4Icz6sTgfFhvVCI4yzSQKvZd1JCZHdXlJI8/aeCZTC8CAYHl
u82pQyoMHDf7YPRZ0xgL9fPmDgBOgnx/ATNoiOPx2TtRNwpoBSa8M5dO97BolGSbx/HoeTQydgSE
8WpnVVHrAy0hmCCF6f+fx94xlh9ToosenU0BocZSKLemae2S+M53woxItHOrkGbt3bxGdIbFe2PB
63pK+fuB59slXsRJMhvcZ6CgAJXqaSUIhtHdO2iUWPOzO0jDKEyNyGyBjEPjmOH9iOwKHjZp0b37
cpwYcKLcpMiP44ibdi/MqhakMts/Ch3Y4ipSfhgwoa6bBI9R/FvktRNwFvVOQZN56UFr7rdo+T8K
imuGE1EmmodDt0RNiinD1Zxpt1xVfvFpBD4SZoK/zF7NW0yl8Nl+ha3DV4DxMdhysHGZYAFhwxl0
UwcpHtcLsB0VmZKQTpj1lFO1NnY6zzfi30TP2dloUVtdXQXQQXxxy1nf6gkruemjVTOJQ4LqsnIW
qOIMJpob1sWAIIhB0s5qShKtR2lvWfUgfvSK/q0dZBZ7Zt2IRn5yT/dAGxxt/QFq7haEKm3grF2i
TiirfxRjipfP4hpc9ErbM0qJ8Gbxg44tOkJ44YzDMtPEnlgU8YfSVac8nYv0rrEJM9nLLy00qTg6
grvtsSVsuUAWFK++u1Blmt/E5Owb+JGGvL+C6/aMfBerkUFSNvGny0s6y/f9BtQVg3sEXC4eRFhJ
HBmCBGgTnubmWxi0osuQYO97t2KcpnisUoQI3GKFF8DDrF6ERFDkOOkODxqwLaGiuvNiom4XoMhe
rE75VjScef103+hB8ftvy7nSjh7kawCfGdPP7HCCPGBICoycxcuxSBTbZFbe6HJyyiXSm5bl4BFs
czXTmvdhIRMGHYFDe5e9cMLCkp9HOvh3KixIJp556BJ3wDtoRBb1MWaNLZnh6+a93sB7elbQD4ge
uVVOxpxrN4yNz4wyzFQqIXa2g+zUgLQKxPy9plSxLvZqMT5yV2AKJCbzQAf2gJDTg4AIXR65qlZs
WYux+LEm48K0GheBnfhdG+tOM9tGrPcKm5d9fLoF1BY+3jgrOgjmU3AJh54Q/NBnjeaPhGIBVKya
kjebusfIopRe8gkXbwoUHQX8yGiMTFgElkakONPJnUoW/p10CqBuGhOE+BoYuKsHANDwbqLnGU3N
/M8h4/8uFcJVObIOQ4nE/iBOfzDQaUAxRwVYvTwrOXJj2XhXVYRiE9Ev5LMi/aa0+Ny16dO/ieeE
whR2UQ8jhDh1t2POIN0+pAEbeS84Pwwslv6yD6Mf3lgso/Pb4OicFV0lLXOg/80Vp8fFT/HgjGb4
XklywAo2bqxJ8PcaQ0PZBX7Bjw5uvWi5gv5KyftszEUgk/vBKRZucYJqdR382bcZLNpAwkYXafqr
50gglX49lpRCBnnkUP7a5PByT7nVolCBEn9Pmip88VstpozmUwRYIg18/Y0qDw+GGUZSHwk7fIMj
truEF9BexFV+wtUP7HHweNi3OXKYcP86CsDmov50JM/ehQ6l7iR0kWhnaXbCOw9OKclWG0FGgoJi
wZW1zSTp/CiA1IEVAvsNHxjSF93RKY9OJkPIVY8v90T31lfa5R4BhnNBvsCL9X6fImn70yXBJugc
lJRxf5dbajDbIEb8mR9RSXZoABFycf5zKYZ/gkgr/GJbqFf/+tbCSCUBsEETHxEUoisGrdg9SuNA
IBo2rHz7ipQPkiLvImxwWBopsfaH49HQ5KvTLwua/2zCn003BK7PIkB+p09qQ3FPPhP/HhGjxMuj
ji9LTbtQI/IMxINjx3sEVyd+k65UKsBKJaAX82cR4MgMgav4rE+ATlf9olwRLnpyj8jZaJyidaW/
TSdyuOMR/WvlSG+tH89+r9Ta0XSH1XyhPg08U4N1K24r0+Y3dzf55qfrKlo6a55AxD+L1hPm8fA5
LwO8OMNPF+N/Lfab1J5SB4yBRBaqTfxWqwNlOxGgdxqNGGm8fJBT+GihM5i1QYz4HSQMRputZmn+
cwmxPqTfa8/8wPJnqdaqRrgbFkP3vWDFhj4rJTHdehG6zYL1P2W03u95wyY/pKBVoiQO8MKHDGC2
VjR3kFM5H5SqP/dTvVFvhNQZ31xHQ20t4967wef3rl6QY661+M9JXZvwtTo84cafwY712P36dQPf
0UZh7VNs8yAuIBjx+j+6MNynBmJBbhxCJ2IejbLy5JmDtP61VBfMnITmQmAwOtWyt62LjF4XmlRs
2uWj5/eM19Zy7WxFQMU99p+UWpCD2u1miiEJuMO8bableQM4RYmQ8qc8YQKbbesExol4adk6HB+o
f9IhST0Ef0Pr5LOxd+p9h88PUQ9mdBEhX0PQ28W29eGZ+GZjvuKdcGMjfJocCVQNJ4vKfDugxXR5
40IKr5EYf0Fpc8WKbK7Pwtm2XjKGGd4RAk5Yqdj30aS16AoKPHOG4OVs26R8ZsnMBNPD7gr94LEG
1GNxu+1NeuW67fPljloyuKYDFIN5Kc/ieaE9kLFao5sWCzke9L8+qZknIqwHE/7p6VCkUHISMUPz
PRpO48cCqNbSzTX1l+0uNK1oVjlehESGQbp1kyOwp56P8RbIuZEvTtEf+ELQStMOgE9Wk/CWRbc6
EiR5DbSl/M4SgUpfECkwfvDs5rDqaf70hc4FqBbI9mCB230Q2yb3plQTWEDuABH/uhzUQjNzaGf4
EfRjAIRbCVnl2ExolpW4251SMauFElyhUYPg6eAymJ+UewQtTcWFFhdcC/1Oydm79lHnWE5ju95/
A6oEU0LKif/zikx9x9c1U+pfaQzdXzTZyplQE5dYQHhAe79sQ5zP0u1ZLO2I80gFlTPubvTCpTBM
C9CAO85hEfG8NSFId3ljqs+DZfkeThxv8My3EQ4z7yzN6DI+V2tnMpJfyLkWcDAZcDuD01WCsg8V
/Tjzr5TW6iihyGmsXa5Mf/WrLD6dn/pJZF/tFiS9SgtxO2uiuNSyGu5FnYXyTL+0648t23I4q80c
GUjNbNZU6NKaWzN4kQMLSfjENYrHZovd1kyc/KMcSWobK1z2bwXtA6pYx4HGsIwFZCd27wAak7Dg
Z/ap/l2RDV9jIHbxXHuMDl0CEEE5dITJ7CASXICyP018ri8+1p/D2ivO4DEGrNiuF7Eq+Ym6xSql
a5nywZcin682hCqFRlqyYFNa1uAn/84exIs+rx12tqK3rC4jNueGuie/ayJde1peO+pkSvXyt9Ks
m4IhVnqDyg+T7vGQ9IF0TQnfNERsD7qxQ+cVUhMfGFv9XTAopX5hywQrWEy5vt+cpug9BMUr4CGr
tyxLwnM/JuHnVPb94r3deM0yQi0dkP546nuX7HNYEVlD2jMknuyYPQ872SS6MQJC7wRM1skmgZ9L
6KL0DQO//BtKiwuo0O7kzVoqDwP5f5mZpzztM5Id06t11k5yUCtxWUIUpbJEOWXoS6k7I7obq5jP
ZDnnzaR+ZlJkU/4Glx2sDPwAnZKkVZE5f2Dj0sH3E9DJIp6M8/SEPmIG96dQQVxfmRcMkEW4ykq2
hzurp1RUEusL0dp9y6o6VzgNIb8GtIshWb34Nj/ryd7zF4eBORIF3DHMuAzRb/FuO9Df2idINdx9
J/pN0dW/v5az6JTfVijpqaG1UuKsiEYOytt8x+GRksCv8RQBmphcGx7DiFdrfHkOptIcD3Qgn0Hg
dTT26OAg2cNe8WMyWCq3pFDRTZ5f9T07ziZiZF+1n07lLiNO/0Jj93GgBN2D8l3bnul6VuAPpxzC
yGTGvue6VvrEXmS3KVaaO0LbESkVtmaCIUjz77ffsSrQTQLSOUgefWgQWvyXJWS6l77yvwqq42DK
Tvc9G13g6DVFB9MAkgzkEI2FcG5FajRvrNwQbdOh6HbjFFROg96avOkz6HLVYDlbMttaz6d0lqIU
o3VzCrS0yABNsB4YQWPG4w9B650qvD2yD9nFER7lD4aGAhmHEyblundPoHlvQ7nlJTidfFLRRbDz
LZxcYLKKV/v7S+ztwXp5xmTFU1JUgDXfOwyZUhhH55XRTqXlvmErjCx/gbikP/iA1MNoqnuDbkv9
GheeKqd/kLcmbbX1NxZvW2C2VaQsjVhl0Pk+7v1lMTyW8F8DlyR3AuUqcBURmZZmD1ITl14ZUBm+
99y7Ix94JGzNNWYO0vmffUA53naNn/bcUPtJ6WnINcoj36mpVTTTvt81t97q+5088ikdxtJiAjMZ
hL5Dy1cyXzV3MnBFbZ/WK+rC2+8MeKTSxShwNBbO6BqQC6CzwkC/C/iHQ9kR36+O2nxAmDsriK5c
F9Yf72qMEDHVwBL1l09hpUYOENo9/IFEtCYzAeUY4K7sx0sT10N7ASXe5OaxpUDBMaeR93z+hLBL
oVAxWPLrnsU1L2NQXTs22QFaFyB5903dD9W7bVaVDxEvS79BzXCdIzwipA2y+LI/jvzEAlOMW2I+
pshhfkuZj6sfZaIrRyEA6RjmOKL+h+4m4EWRklAQTTlsW6reJtUbPIrCp5bVsTa7Gk+GhQ5NnOTE
SFe5EqTXtnYU3yt8IOVId1irDL/ukVolNAzCcOlvbloFWgt1KDlBU26ofsyspKNh81wr40OoRzHa
14wls6lOSInLPX3FWE2q4HExcpfeg18GCtquMjJ77806w2k0O8Daf1qG5FVpb3itakDLj67mTLwd
ofEkoSLEoTwdLVzHhu/6rpu8Cg4L1csJOvGqajmplb0ENBHrrZlQfyR1A6CulPS2svPZzsQVd8mu
b8KwOe1mix+/Yircctaqs6o8A0JrjIluxz4ROjM15M6oeLmLa+oF/vy1StL9xH3cMPVYz7WmDJJY
TdXdPTMK6dzOw3jlL2QcHdEdSG+icJ8TCgnyLRjfeBU1VjpPMyppVVQ1d8nIUEiaqEVcp80OyrkE
5lyRNk8UaL2IguvLCTL7AMw1dKbafziK8ImL2fD6TzEezmYs+b+EGHhQggyGiKZwhlJ6RDNRdE0r
MOGIUWCGwY13RoI/LCMmV7Qz5SVLVx0Pzit/rEm7OE7WEgNgxs3qNE66mTku7yRDcchAha0YDrk6
p8jqXr0ZicWXQvW6iGMCVZ+Cy9AENmwPSPI+7MiEfJi5ID0dpZI++SxGggIjo6HxhGPEzVjH8RMd
I2A38hFNL+d3GHAhw1i4t7VqWgYHj4NwoTaPbh4DWBoI1ZCpF2e71/LhE44S9tSyTOyD9QFn4uAj
PjhF+6WFEnwDmAw6I/uXbsBxuDhgOa1kCzzrcCxUyk7t300vUsxSbZd1CiECdIqN2z5FKU1VWIA+
VZr5jqF5ABj0CniZoMmKFEW8901K07NwFEXAUp9YbD61On8jMyIvheTbgRZo0WmI2wTF3eoEKspW
oAGQ8vKDvJt/oH076CdVIW98hsQvdc5u8UPrShD5aXRFq+rvs7YgWo0kQvXP4Ezebk/HVyiVj2UC
YYrKUvdgdyflaRN6wJgTPromQosFtOzNgm0fIIlp53tRVjmA+mEDhDGFofGo//3xBGe1Y4WUJXCS
OwDDK89ty+CL4oiEiIqjITvFoDjnf4ksxReH5x6uuJPbBiuap5yzgsNv4nxajL+nHHzDrZi2OaDC
Kz/7j1P1sTwfdHjvyoXL4P0amEZEwyFVO3SZosDeQz3pJRnsLZ5c3Ra1ePfcH2lvUK1qkQMovmO2
cuMpq42DjKjTOpr6ze7oZnvhvAJJcTmCoBsJQYKn4W9jIVyt7e/koxcUCqVXDK27mpoS7c2itEtk
1/TECy2+bjjI+YdOQQR+lkHoY8YTAR5y0eCeOLXaKkrIsf4UhivKjBb0GwkKqfLkOFF6LGmK2iBJ
njhfE38aIKhGVkuUe5mrIxqyzhE7+KE5xIIbWBTIvoYBJf79WbG3kJQlT/KJ+fcLCnPd7UEND3bI
/pLy6lNhH/P/ulVtJHsoSr14DkrdPHPx0bQ4R6+BGMdWbA92IzXqxoglurwAiAyoZ4ZR1xWIeeuF
6RIKLLQK6HonF1qeN6yykJug9fbMttW+WfWOxXg2Ea9g69a4HUrlGZS4KXZx9M/0IxL73YSANpN+
M8Sztb9FhUCBxX+WJhqEBINmN8poFBsbxUWb5F4Q13q8DaraRfJPIv9zTmYn009G72wy85HlLsbF
jM1Uvca9ryqiRBnmom4lT4MT+daPwlN0E8hRSrIl/D3UjPwuCsmwoAc56URmK308CHfAevodDB9/
TciEL49EVbkDDHEkm8t1Mx9GyelQY0svRtop4DIwmVV/D3pRbZA3SFLZFAvZDbcalrr2VgnXFKxG
zsFavn3rSjpUs4RJi/X0v0nu3dM2KOORl+5qnl7DSZtALtccolsXGKQawFwLNdKSBPYw/+Y0iYg9
Eblc2jlNb97S3V6Qn09qmncG6EKBECBYzVfoTwH4LtB3rRUhrqj82wbBX6UqO4Lei7EPDyx28zIB
4Vljjp+aC/On5jPbH4mFstBcO9rPMuZxzON+VBppS3p4esYOCXcWPGixJtvibRlSxlAZjZ+72MNc
hSmAxOrwHpM49wcd+3zaqFmWRaRpImyiZY/7lNhZZORsfMNGA1nqOEPUx3ZOcCdBmNEmU78zTLBx
dotsLpeIjmOWM2gah4q8a/orSPw90yull4/jOTM16qOrEIcS1hl+Btp+rbNfZNJQPQutwfrhskzl
UNCdMO9gvxaYDqTRWvm5KpeKMSFKyyZtXv5L/HPGbVIZevVybZ2pZyZ+qXdkJVwUdA+iHZkg3C32
cyMeC/D0LUUZuUrv9k83+WW6VhR1ZdWPV8ezyXbvyZExsn1gq9CoHOHoaUn0AVnsBQq6SiK1kmN2
Idkr5DyjR8strQdlsod+7CDFlpptowQQTniIZO73ARg4VJ4nT3GdAeNroahmxxs0S1PEet7K+q+E
oDzP29bw4Lerld4Ww3Flkust6f8+DBFyyABfN379mmscIXk6BqYX0pz5AOUbPfQ9IFqc+9tUWKjL
Ri6Og1+GYyHhhPzeRWKI3DyPtA7DrnYPi0LC15ps+6CLjCnL4zVrsj/e7HCA+E2QOGBmKCtjqPCe
8SOvP10/J5KPL9yEYgdWVjZfPdU7aleNbpc+WW/2UpxCZBb3vCbK5RwzhpVekf0dLbbKhNiDYsNY
gEbe+Pb4qIcO0vVXz3JKF5MtWM0QaTWAIFUWDjwguekV3iDKUHygQ6L2s3d8+f0Rm3dUuyNF63eS
MsHX3dCoVe73Na4jxewqaTMGqRWiRHH8LN9tqPhcRVoPydi/PimgogqtVpwwP6/avexPOo936xXR
U7SdmJa1gzz2DHCzdSB2iaXsV4siibsMx3luZViDMf8n8mI/O62tmu0Xmm3pETeLnW1kh44w+Y+0
LVcVe7i5ptl67RAYpTdZsO+XAmkPQplNW3oYBiC5Z8i9awfhzbbOOUGTjSkVP8h/K0wHXADYP1ua
HKYXZDUxEckT/wNtZXUC/g4jSOPlSGA+hRhUL+DCfKndvbqdY81g8nusle9ez6sSm1joQXiVbqvN
pRSosyz79cN2Pj3WTAXzxxT89JTEZV4CqEOXxpE5EoyhhJwOnvHpJvQkrCr03sXo/ozrGh/N4H2o
/SYcTVfGlg88VkF6j0cU+Bqj6OdVmvlTCmKXJCBsk5gg5SpYF0mJ2IQ5rTB3p9gp9Az7vf82IsEI
8yD25Tas7pvLdMU2e2VvNs8NPe4bx3IVib01p9saKBjYLpXan2ixdGsr2Hj0hx3D6UAZ7ErFWLHP
h5YkWDjpPhe801/Q5W3FWm3TynU6DzLg5efohtwUL7psrY7HwPKT6iOxu7WSHjS1wTTWlasrOlCO
gQpafsJcwzDaV94MUBOgJhHOD+VCe1miXZSu3q1S9YHmUkChz+HNZykp7hoQKo9MnDm342m2Vce2
UkpcUxdXXPGvfppIQzU6DPG1YAR9ZV+ob7G/ofCeEobbHL6b4W/Uq5uWFA3mUaAR/Fdkfr1J/vb2
KVFj2G4c+heK32jITqNmHQCEitx9deB6vcwvs+a6hfebwzD0+SQLKBWMl4HAyLC63RKQYkhxZy90
t7KBPE+sF2GUXfsw5WUOlwzksiL5MuNJhvx0Cy+WYSqqrBw+/b8pywc2gya3816sKYqnwU8VReco
1JItX9mqZ6fgdr7wpfbSKZsnPdHx/K4iwB4jyVe6qMHx3OK5TNI8CR7Bj0b2FXad/C4jjZ9XDZNu
00T3Qyu1M5JpR/Qqbgqh+9ejkAFdw/NVOxSZHyYJFUbzbOaupdp4mWg652kegNTYw5zYqUIiA3Nc
wys+clrfi+OsH6uauCYWP99cDKv2HT5DPEh0sGLkKN2fbPrHRqle8K/oe1puPmKv4axTc8IXudcQ
wFFwrNoii9rhdB+egUTfIrtfbYNYbVbUhPzpJ/HDg3g6uRe/p/8YeQYNMRk7W2PkRl5ZL9F53rDW
r3mV3EyA4y6lVd0urYzPaQbn/fZYapDO1T+oLXN4dYS644GcVD7EPdDMfgCyt6Et9/Vf8v0SdS7l
xpiXM8AyGiAF7C2kgWZftwBJ3DrkzUSAb01sMvhiZlz/l9dxFambEt3t4E1L3TcjaXY64imkKs4r
konamq7/Bc9u4MaT/zR+XUiDTmd/5qFrIIBVAez5riXH7k55OAfdYYhoNvyJZ2HmtTPK6VtXrhRR
eTQN3iP39oWAI4UjUmjq59DzCbLuBCkSxki6yg3saW1n4M0AKvxyzpp+IHdPWn6IFamWaf0aIczX
2Xz+dsv1jY78w1oEIYxP9yM3wkfYZV5fXpq5VLMkEoO4lF3HD8utdC9ENA+eA6MGzVk4/YS2F03V
DyKr6FJfxZaW9vxydjgaKnV1Yrx0YcoUFMDS9gUtg2Pkg30trS4faeHV50clM2vUaO6FOIaSyG8c
mx2oooWuxT6IvmhG0GoMgCm17X9Lkn3hKnBZDwWFI3tgVGL9cNSY60gfU6UGhaqAjYDjC12E3GgS
ltiKBuHbYV+Cnb2FTkJwJr5eI6iC7UGEYolR6XGj08J7lq3YLeE/jXnNMvLWAJ4AD8km8Ib7awmf
lgVUov9QCl4LcWt35WWAcJqM5C1yLUmOO1E92k6r6aeHmjTPUR9oGDHSGM7AxwRcv5sGKDLyCoBG
ivjVj/mBqFexvt1DIahVBCti1pvmWj8Lxwn1IYtQxZhu2SZuyFZUOI8loVc90+USxprQhrtX1P20
pGt04tYCMVNvxPtNtc6kCTxFZGhJAIoyf+EVM7qguxBpWuHOZiLpNuxnDzXSZ5Wscc4/nUNwE3P6
f0zszfNF2E7/JVLUwy2nOKu4uBMkV79xgR8MzN0PvNARPz1UexE1Md9SSZQ67y+E88szz0CnRjET
g8O+tH4I4XjoLSRwh2FvYvSo+QzfYUUtKLfIUgrqQBC09k+4XeT7UZOg/5V9xTi6s+h8mCEKV0gj
m5juHEGnhAflY2IrE2/xYb0fkHvo+jKofUGBHa5dRGbdH/zKmGkDaum3Ngl/oP/giMHLdG1BLlJ0
f4L7rt1DEVlwSnsUL0tHLRs5v2vfAYU6j/FDY6VmAfhuDKMperHH2k+8QYGEYuZE33CMSpqiawbh
1TPrMoCsr/8hFhPbszpFTOVT+5XF+5/jbERhnlPeAfQQzo9bKb6+ErElzznRZVwvwjF2NRZ96ql7
jiB8xTI62kMrpj2sIxvzYtaWo02QfuENAnozOp870NkGde3OUC7ZApUMJ2dJ7Zreor/cI8RlQTl1
19slpgcVvS7mjp6HWVRAvbD9qqvjzk55qwDbECorzEY3a+YLTm+LazE6XtV+av57pfTaCCh+OWvf
NIIs9qAYRGIpU9N/FPbRI2YBwPfgacTUU66dBBY0YKjddD0bb1phnlW5OuzJE5s1LNh+OMSHBzDX
SkdxvUxctrE1TPKItb5F+uX9KtztXoWHgypsVi0623cgckuDaWLdr/pbuQzth67KcPEU81uG5o4q
rC+2NNBDkoXhOG2kbOsCta0fAnQRYA9MtBZEDdj+RUb2YjtyJh5wvlxFTAsleQ2574pmHMCYFcco
a82p9tKUlMS9Ywu+WaP7DorjIgERCVzqv/XkMs81qQsNrdVmgDKJlFEkd9XXo9ciZsfHM2XMKy0u
R9F6+JpgJ4Y48oCGS2wSCTTBlw3JCHy9Re4HEhadWdb5O8SQ5mc1hTRJJhEO9DqB8YQyYePujmOw
yXkMs8kb8Fss9xiG/vHhC5ivdlaNgXmo1XJzwnGikg9HmHXL76I6v+7dGCKInd9HhAvZEw/0qdJz
KphI0/DD+3RjwrksjE+iRgc8+MREJo+TGrK/2zMMeNtsWWv1Vy8HVVPDnIO9+aJ730D1/41VAJQk
pkFe13j4BICkl+FP5OXsQHejCafw+vObPFhqWPvrAgWGC6PZP/BMrSW7mjQ/OG9XvBdyyIa5Oipe
mob5zTZlmp01AHO69SDOL6uyzzynJqFtKv1zsSs3G0Z/RRHSSdp5hWB8G+gd6hJNSztChD5LNDs/
hAjPsLc1Opjf202tUBVsO1USAcnNhLZ7v6XGiKm1BKGxWorkJYNsKJ6uA3n6NNVaKNprKtZSY6rT
/kFOGha9m667oYJfR1OCzkF7i4Orz7daQeYz7mCsbw+z4bqCWN6gk9e+Ib+xDOIP94v6QJ/bIaVr
R9kfnZ4c1tQKBFhB7D23tl7dZhA1g36EI4VZI56+UEQDVo0dLPN0eIvQQWgw4ACVSOZ1U2vx6ZqX
wjtaWNIko8wYFdSvrNaxTlspsNqyjA+mz8a5D0QRF1oezwaq9G2g8NVpVEUXJe/+gR99pUkAlvcZ
bOJVqUEJcA6agh9bIADD26MWLzuApWfmrDxX4HcoMlY+pqhli+CGKhBPDjEtvG2pL10XS3qG8m26
ISVsJwJM2pI0dUWF10mK8OEGCq2GOGzm14F3KxVZ1KdVyV8pBiz6anEeADryalW1NgjDXzzEQdoy
YNNmVVu5ZghTf+Fs7QUtOlyj9NeYPwAmH1kbk3EA1tn/wkQajeyYYpCJRT5KwkowiywivCckdgZo
h/id2TKj30dJ6afHZua2mapDjKqSa2TjDP9wDnPPTwPtcfRmtl9JR1b5znwx5/nXQ2aKBOmKUt9U
4frWe92D8Jo+94mJ+Ba3BdTkgSS1NIH0PGINfNgSC0p6QBiijYwHVHKJXCe7i6Z+Yg9/DfmAALN7
jRp/ESZA7zdkXSY1VMskq20uamo9aOU68FoKZGGIq9r3NNudFERKMhiaI9twfVntIxO27/4NbepC
C3QlQGO8/Nuqp9aMgluH2OjZdMP4TCXyWTNWC4SnLXmGsr7EBhnw629s0t0T6JTF4RRGJBnm4VSZ
nN9Se9FICoj6wpqvfz7wYEJ2EcgaqnR7q/GFz9p7Xso+NSJYtFRkCv0pB9mg2KwHjCNCThdtaiRf
lwBY8Bkw1DFGrNaQrkFmkL6Tm6J5ULtMmpIdJ0drXjSysgqR/qq1Z9jzk9HyjNjJiu9EBXaoj3R0
jno+jxI5Fi+7wTahUh90yBDGU5Bm+9JrT1QKwbdSpCxU/DyjdjOrlEF8s6WvhyxtwWq9FX0rygPN
O3fAgWJGl5ZhDcBi36UFDUWrPG/7GJwxgRo4FfPTicU8vDawSg5dg1ZyEJYGrTlk6cWptbpAsq/1
H29vRuV958kzqGU/IUttKf9UYXS2fmXjyvFZxPV8ed7tF5AU/m44RippKdlVSwU2QJEzDwPq3k8D
/Ww9JFNIv2BmmFRsXzZnzIhb/2t6hPaqysGyDe2NbZgUegRDTnDbxQoP3/J1Qp3WwMSz3EWWEU7P
48gnyr5fIK7Nap+XQEz0QkobWQG9mByhmnxhr+Nb7rtvLtOr2ct4RC/6NUftP2Ulznia0TELU0ZK
SYyb/5yyPL89DOP9pcJQBKs33dSZ6tApu01VWbwss9IvYAphFF1bUw+N+4cYZvQre80iAycS3FPL
OJ1Fq85ti9TiI2N6REdKxHuQhSG3qhXjUiozZr6Gnw6JqncXcrpCd/gOd/rqrH1uN/8mKu38UkZM
Yudp7UJkDVet/EqqpxjFvLdVUV/RvBG9+4Mu9LoA79yiKiU0vI5ZH8BhuWQEJ06599ZvofwwpAro
S2ik9dApz5zvlMk20x8QM23U0vIG5IBu7S8OlBqgHaC9W4Xzmg3w56WsZLdfAIyuEH8QLI5ybe5a
38ia1zBidEQHcmOUSNgSU/jRKOohPg6x3irMhRXWQ6sfnv0EAxghmNYarjNkrIm8CX4Kc3AMIp0u
PkLqNzaoWDcwVHLiBGjR5qxknmW5mTLN8fbcrmLus663A96KuL2825yKdLrOb+/iQQFcoptjyHJR
PSq0WIiNitWlxaotcBCOuJe3pcxLi1jbFAGSg3J5ZST/f/LfB2lgkdRb4M+YaNzYI5XhlarGBLJk
15j9X3kEK61TltlV4sqNCg8TUtuqHaECKSde+F0z98rIZkGhRXD7HFkjv7HXCBBnBWvkM1IdPvmQ
ZvAjLYha2H5xNrj6X3Gmyrhf+33CbEZ9UkGqatzHm6pZ0VLoL2DYIkEaIWdW8jxQ0ZU0SulhL1Pr
U5d3xf7HnGOPb6mmFj5GUR5abeg2MSfye1wvHLwuCk10+AA/pLE77eoSxNBzoVRie4lk7Aq/T72V
QheDVEZkpOfptD7XiB+BpCGpl37H6geRlCow/SxlwuLQj+H2og06ntz0Bgz//7kLt9ZMkyiOj1uD
A9rn3TcdGHNhYil+hBGr02y28BnFv/qXmRdOx6zP1vy/cvymX3TJykNrfWht8AuF5sIi+RIWokIq
Ud1Zi2gXaHsZaYYPVCMXCk8+t5kt9kWeD5UqmqUd2vrq4PiV8ko+F5OlOMnPX0eeNsHrz8uopQhQ
RzdOpEScbvy1vxK14Mq0cRsdwByE4P2vKtPLjFWO8rg+0FYRN4zHvhgY4DaA5cje3ggFJtNp8DKy
tDE78LZN17DRB/VVtaZaLBnA8EerxQX5P+r+2n/SU3xC+SmkAw8ssDOiTppggvfRki9wLIeWhIym
h4PvxOo3OXK4c6FZ+vVTRcx+v2EiIO0/F6bf5uynAbvV08ogE98hCXT6L5HybixwZCiFekxty0+O
Wpg+/bVU6WpvKhRpCt7YN9HqY5buuc41SuwQAQSnpEK4s9cRyPrRVOqVIp2LBzc2yWCComxWfOAZ
aeslPSrLDwYnU3h9mqyeNbRxbvaWRvXkOd/oFxN/JqePw9L/gXhGxJS3rmUGSDDBY6KSElRMI3eq
EjvviKqbVefe9VDMzatzzNPmtWKiXiX48lEIOTNc3tBgIFbo8GupCDlCPXTvdpcrlxtOBlRLuUde
UPrXmfuzowHpDzyY98XyReNzkbkncw4fEP2Jp6JMGASPadnMA0GIj58AhVBPl4/8PNZGRKXsLrm1
r7MOKaoS5PfceOeyZMUSJm/Dw5Zve9I0T2E1Y+83OoLM9bqw4zDcugznJ5PmbniwHWG01ceePEri
nT12tgCkX6bc6WAAtRueUIVskZpsGVnMCC9WTe/XGLilWrKO9fHliJrHtPqYoo2fARKEQMI/IvYO
htvMOJZyWlel6kjPh3xSQzgXzNVRss8N6jF/rFsz+r+fSQpMw4XhmHLdIBVghGGBNhVVdGjJYStM
GlWbTJZFg62vIZlIsZSYJWHgw1hHdLDWCbeYNV9tIcQSnPLJHqzwGH0TpFpQ5F04wc/1clX3xcbT
/nJY9RvMBNSrrPiAhP34Do/nJ4nbCSfVu/l6I7bTYpg6TBB+VXDf/OaZxtq/hGYDaA2y69vkW0g2
C9Fj4QA3oBnpUR+oT4tTrw+7bHL3Fz+LnjIBPWtHJ0ojeXmoyfk7pZoUzULeoGIGvOwev5sHZVFR
mYyqMFgtYQUi2yJAEkVec9pYyHomRBdYx+lKcOoTM55E3TZCTQwN/5BNYdnbMov+ew71payo9X3i
ZVe84qCsdGjVcK3ShwquGAYSQNn2GGfN77/eA1ivm0CMXcHgFeEkZ8l6lbZU1QUwQjJf1A1Hpe+t
sm8FDedId+hU8+qdaDwhkFjTfGHdAh32aIYKnYB2iU5NFEqDGhszwBwOY4KHi6Wda1H/FR2UWPeC
beraVLY52370m05zGy1K614A6Q7bcfCJxE4rMJVCntiMGNto9s+XfVvl0l06iRuMuHwc6L9ShbOx
d7myAdtpTzSYude6HjWv1jtqeD8VssG31z30gOFZtllerBBRm5MDAC5Z4QZIdVxqoARL7LiPMkrv
TtLg9SjNoVJNwYD5FbbmjSaU2EY+gJsOi0odphXd3NsBXL8WLKans6Dim2xF8bP35lCMmDQ3HvLT
eTTjpEs8SnU93loLR/LoJf0HtnriLzI4HKepliAhOTnSHjXS1xc5o7qm5ifV55AlJSiyVWRsQUaj
V7LJjuBBoweGyAEBM7i0J7ivUt/eEinPNFg9vtTo5t1GB/C3DNN9xCcGZ/NvllIrj/QqW0Xr2mNK
AGK0Ik936eJm4WsWTsDfQkCZv1fJKt78WhYGJp2z2WqFAJ+Pc2MmgAfWgjzvArJwcDWhE1HWj+Qi
slM9NWjyDJ3Ee2r+CQeWYnoZYXSYKSF7LluIDhA/yXJMrZQ0JrAG6xRfiDzjZnrfjFlY0vnpdP/E
NQoUL/CfdLDQS2MRhPmNnXMFdgCPRz3zVolaXfEtJcEWZdTY5q33l00DmQICh0VL17mMCxoj1KxS
KnM0jiitPEskDpIPPV/8RT3dUe12yV3yABLtIUaIR0xYuxixeEEjJENP743DaDV0kTZbPsenps3G
xeiYEtEJLqRwxJlNSnfooT9KWb7PJrVQQ+8SmyyUcWf5Dao3tssKyqwujLcLiiD23fT7UvQsW8lV
aeupnG5tuF1h5kdogliAwqjUQIWGb0opPoz8DkZZZn8W/LogaFD4x2JmvcEjBMTBKH/hc19OPs2d
CjkGFcxPKD0jZk5Dh0plV5zZxr3LkI0eDoOW13gg/rvbVrJUPGR15L/C9tZ9dL7tEgEEUkjMwdCE
ZchuPbcBJCDoUcOZfnUrpuTwokIbKdmKavt0A/BKGpwDsppzMvHdzoGjq41cmEBTwfmXfKXOVJ/I
WLTX/NIX77TqyDLwU/0NIKg8HtaH89Pwn/AQOSos4bc26fxywPb/t0hp0ZTLtK15Dq1YzmwZAL5g
Lr/5UxHUs0ilymSUl04PrNQgrr09lPgipoPNFJRmaZFLFAAi6dUVV3LzwUTmyPLNB230dykx7juV
Dxf9kWWZ8mVDKpw1AtXKurcY48Lu4UoIOzpuQcyHbqKMlpnYWC0JmA3QxNkIvp+/iFFWYgv1s8jd
SPtch+XqmP1hbXdxYK1PJ+PzEsBxcP4LKm0/cL7CFXL8VhF09oueeSDcxzsN2a31iuEX6oL6OPDG
nWuwX8wNOWByUMb/PAJ+2sasrGHKZsgbvpOtCONo52r4h8XdgRja0lRwiI6sz/qesUYWPVugZi8Q
w3zVruX4NVwkV+qLgFg0vf9uzlE9kp2f4uiS1p/qVStwF3XtTmb+2XMqu2wlbgvHpjOaC/oXSCpt
iPI1rx0kEd/5LbOXncDEkfdNPbuiHoEM2uwQn6dbTtTS7A/sQ/t81a+fEQ6f5HSCR46OXDmh/GsG
helWbkwLao9bYH2eEgxr3HKSha0ssSak86QE+qvQv7loxiA15ejbIO/5ZtbBRZe+Kkqchcxbgr05
CXym/ab7H/h2bGk2aohjzVvf1DNyOxIPPXzvmU0yULNe0lCWyfhfjhxkIGle08qk8gvl/tH9BaYQ
63JKh8nqQNIa9ev8JMMpNuqdfNaxLDX2WvvgESETWvmtuEDhJMFhLBiq3INQeeQn7dXllhqgZWj/
o480d3RRg+0Me0s98tGzhbXL0zjRVNcdkrfR9VrN8eQRE40yzjpJ9YDvEiN4ETkZAeWAcUmME43G
qpxiRbmRE6pI/pHbbf79fw2n31gbaGaylk8cheu/lyUxsvICCd4xFQQ0nYmYK8+f8BthnVg4AZJK
2rO4hADlskPgV1gPSQGuCFFrY8HP2d5Pc42XSEPTOXSBazMjMfZGwBlKny7ChD7uFopUW13MaW2V
PhjcjmsWwj5nGcdHvKjmR8AIyfNuNXFou0j9QDjanLQnyS3CVO4n125xsKX7QBTE39L7G4r6VwzS
nY8uanKMKlmxq66Ty1SrCEu9qYPlzC9rjk1fhusN25GKZnrL9nM735hNhEkv5FTdIsuwjOoBdyGG
93C/7VW92MnMRe/SV0tErtLwafW1kDg3TddaMw3CvjMHOAxo7J9IubPovMgCIycYMLLmti2eT1nl
ZwZUZE5I0/+sHMFGb1auC+BSsmRFsCZQQJKIhuUvWCpmEgmXOAPeWutYsxEm4S7jDpPdKCNa5pMf
DWdud6dBAcVrGy2UcNPuEYWrr5n40vCHFe/aKoNr6SxLYLBRMa+cZPYdhd1436+CzpKZKDpj8/U/
7DRWv3RO2ZIESoUn5kHnxxfqpEi9ds3EgrmKmQFFRHFtsHh44cQjo9XbAlL4T7p/+M5dJmkk5YNq
bG5oHS9xKoJJRDeF5gy/XbHZTo3WGFnzVbcKx6ilT2XjlEFNCDk1j2ga1DWV07vSANmqo6EFhvVI
71IAV4sHQVmDhsJnZevCuPiDzSin+XjldOKauuozeUSgfkz8y4/L4yfxeaOo2qWco2xY7nHwe4V6
yfJIcEF3/1RRDAkZPit0PbYejKJWEWIVxZWMJ8cFCjlKT4y/+rS8JmT4y9zzAxyumUG7x5O2xEJ8
4k+n70i+062UOkIyYustTfbvw1NLPaoBR61HqZnNpbpl5vcTzp6q/JgVZygWIwD9MrN+Xo/zdT4V
iNeI6fuxztaCx8UbhRbvMllW7iWWR+26rsYM5sM2Dg9wFynlEc5v3qO4uy63u+44zzk/CfFp4+CS
Ibnva9pFiEu/BtYT6bDi0YeZzBEyRmr/MlPRQEtG3ikx2CU+Qh+HiRo6EmoxAY/7FcK4K5nkkNvj
K+IXRN3kAHJChYXgqq6JsRzqBeg0/4tD8FlppRnug1NsjxvkSwvik8tYukP4sCHjL2+l5qbJMVEG
WlGujLMmO9F+KYY3PZulv3AijPbPhJzYdqNAO9dW5WCqboJD+/HpF7EsnGO18JFSvLxco+3yOD95
AJ2vquuzUSTwWMC3TekmbH0AtoroWpk3yCwwncXwAxH9HcLEO25Y5sHkY0Gfsbqy1Rjvj2uvMm9f
F3pxzLGpMwLzeUUnSrs/+qXKDAGNBV3izKNww1D0VtrKPsQo2txiwKFBARMNyYOWsCrfljsBggYS
HhPeB31ceQoHTkp/C1FVPO91Yf4gk1s4f1dgZKNJ9a6AJYSFVLeTg/cZZriZ4STB6BIZxMJmQNhH
L8pgwnCNTcGj2QMaeitCBt+A7/IQFhNLO06pbfo1iWdCZHtAJseP2yE8+SASis4LdCHaXy3pNTZZ
yZcAroS9gP7SsZziFN8Krj17l24y23hrRxiQpR0O8bK2T7+UakUmaphzbK7uNacOqjx4Vr2kGwTp
YuabOY/l+0hqKKscuRvppLdm3V9zLebURs+olX2YtItroO7GuvTV3l2xjbgEJUC2cFNsK1DcgZyN
lLOzLRoRGpCtWIuX4Z4Op9407fh4+adPz3akV6uU9NbLct2VYm/ndA7GQ34surmHFe9W5jVnNTfy
cImNtPH7pHufdhhdQh+H/KdP+kNm54byLNYVwAoNvzD5ypkS0tJJ5iwWb/c15NQ25smrqSGC72f6
Pvf0jpIG16DTnm7J0efvlwGh2nMFEpPeAZ3WDRECTSlytR2I820gTSazqirf0j17k5YG+3YRwZ0H
5hhim7Mue0Gjck+49Kd2ouMyNbvNt0jPBNAx6f12Jn1Ml1HM70Az63M7EEyoLChzQviDFt6RX5Bi
zXe8lV51a9wukxConKFL4FsLcxSqXVEenBd7Et8WEh8qWdRI3ZBDZSR9BCLnD47ZbAoN5MqEpBXx
SprpkTyPJqljy7shfLhVlMm5kvGQXXATrNmx6Jn//SuJ7/Zzw1o0YauGa4nYSjs5v2jsLS+FaS1q
vIQ+sLnL4bTGoFGCLrI/MujW5KCO8ZxJSaENE6WhmFnSf+ZVn1A6A9TwZv8lY7DZrs7921+eVJ9e
RDqO1n51SlBmUbZagjU0w53NQGKivkqsbvpe6LnJq6vCMIV+ski3y5NkZdgkJDJzipQ/T3lha+wt
GkC1Y26pQD2OZ0zGQYTK3qbQX8vBGBn5kS0K7WbSgPWcCh0EFELwIVrZ5rT9OOgey6YoSiD3rbMD
tuWeBmrAluxN2wlPh6Cy873eFKaio2yeO6Rf9umFZFWVxxfmCCak/Wcwx8pGd9yeuBXC7rEe85Uu
qxj6Qpq6EVEXjgr+RO1SCHnMqNPX39bUXoDzy5UrVoIyxe81GLnZrQp3xhIGnsteyOb6gEwLqKxP
PORTYEyOEbyUnNx79sesZpOLuI8JAUGVKBwSDzONldHnxDTM7IjAlYd5iVVihHWEQZ7Nv1qG3ry9
r6xuq62cb133ezDnHf4kDD+5soWfEFSI5VdOm2ydaPig6ccwVo2N4JB0jezRqxmJnhVG7KDzqr20
uW+fY+XesIhjOqRVUsUiixu0/gwKIMHJCJzb1hz0vCYXpzWnhc5JFdjUSwvypj8kkn4FMsw2UeNM
G1ClLUeaaFmIH5ZTApzWOHZ36tOF+fBNz2RFzjsHucqXnDLf2WLmgxGFcfjesFu8ml7ccWVmdtio
8vpsoeEORSQv7rsRfIOCbsKQRqxT4nouLtDHlKLc1DQea3YE4GWCFZgMNISdtTbG3JAfummVaw0m
FxjHBzgGrxqdQB6e17Qq/inBB22B9A0UYiCQXgkaQpucOiwKgigIApXMSIT+n8iGS9brHJFMmaSW
xqLa1fMrQlCwg4Sk/HxYVN5MJc+F4YRrDkS2FOlIRSZ29oEnjPTDvkKnqq4PWkxt6uENjt4sDJHn
ddAomtWqY0L7r1MQNXSPW85G5uYyHACdxtwYQyzHEuy8UYYW7Kn8nDEalzhvn5ZIv1DBX0J9vbZ4
Tppz1CHaGqDAv4k0wuI0qyBA0PPC6mDTuQqXT7fHAczSdv/XDB7zuKpUNHMZLVuFWIFFkETvpfBC
1alQBKitlFiRvqtUV0Lj6wEk30tIVF5LUIEXGX83OSluDd5lGN0kM9W5O/zSlxgm1YPvRPOFqD7a
79SrYyp1X5tsJjHKof21SgDsGZraOxDpfeqqCG49jfrqYhytlK+BImTFWbc1Kkis7FNu4rzo0FZF
iIiZw72JTT9HVXARiZbPzLvDp8MBPdaMNvSjWkMZTzS+qMRf4+N1snJFQHjs/QLniLwJMpTGiOUI
rEkrBH+NOA4AphvuBev+NLwrUnB/FXL+D67d/3X1ia6pkkahzn0xcrvuDNqZ3pJDbb5rwO9TWgNM
g5al/yXPZksonuxu2MZEuX1xvWv0GbGE0OlN5fIOnpSfA6v97+WxoUjGni8HgpN7wpev1jhmTYPB
2RMfZp+8kG6jZg7rzAy0PP8VlCx6j9FZTTROJJHkKxxoq0LqF5hdW1W/Jkf6JFzl21EgJLLaMhr1
LJn86MFZhmMdkfoLufk5OlQZGyWPhk5bDyY9ZlymjFsU9co2cNb9M0v6JIOi8NIKcWVDoAzsUdzp
UcJIzRNjhOySSv0l9VrXTnoH6PV7map/bLxBfba8C3gxaQ67Nbg8PyXlDw+9GEeAXBOg/MlaYayA
QiPFvw7BaZ6Nm26pcYKdQ82jtWCFvQregg7Qpo7Ax1/ViOuLq1uv7wGRV0ks/JJWn8Wfpn9pp4bJ
c5HUbGrIfwjQ5O/GtlgNKKpWRqmEA5q8QwMJebEMRD4scQ29QGhAt0TESq5RoqJIYRkxAw4iFnuJ
LoSFDFSyaoEXB+6c94NL72foXedX5WJUJAEV+/l1vMqQz6x9RLz9dbQfmZp8ye7Xsa8yhfZxSAsB
cBz1YEbWFHP6aT3uWnH4muRbVE+1WQfMtXX7AH4Qr3pAd8ePNIuZsuyghqoWFqM1dBGVgEwYqJbx
Pj9Qm0s4GZb9R1YsZbPR1C1SbaJdwvvjdiZaMqWaKPNLRF+r6kTGeBIr1TYMe6lJi6mF041HABTl
ZRkXRjgOENnslnn1PHLjI9GnokMoaDlUx4wFL2+p3nJ2vzwTc/xTXyRis+7Ep8mil2vzXhHf6F5r
YlZUbWdEcPWC+sM0zvMADozTEgNWI/0HjSC4/cY9jMLwXVItJNG8Nztnqn+DAPaR2yjsnk+HziNE
nbLssG1JE/PJaTO0I4wK3D4p4bisCXBTTrUqJK8houfrsgnGQgj7+pQyuy3ChihSvE70STuD8jq8
zxQd4dLA4GGPbnTTgcBrT64ebCuNxYmP6nsTfz5CfWS9K5t+z0r5REXO/NhzQgd1AVrrro3CYej2
OmZYtVSrxNQaKgPdEyefoaywppZovTN50Ktq4N1T5DdT9hZmV+5yQv4rG9LtT7DRDjqhkPp/u78f
evxBKpqE9NgOCElXADf/2YrdIdUEcnh2burNi5Rhc0SpUI0exzFJ0cuunD6O0hzj/P37UE6pj0ke
QaL4EUGirW+X6UKAgwxwBEwEdgx+GYzmNXcJymxuLC5Z4VYc6iHacezPFxsOf7Hzaao3kDlPcaLq
A7OSPSIkaqVL9fIK/VwM2bWcCGlcreYCSOF3hVPV5dlrpbF1DgU3e6CsPUmduPs1iuGLJo7rl8k9
FMc4PlrGEGH+dVuHpqobsr4GFe3lbXwPJRxJ3LXvmzOhWHwA4cdSIqzT33Md4YatFF7i20gYezeN
B77keKECNe9M02GxiGwxtKPb4ryoAiLbaA1yw0BZvhwNQ/4J1DB8ZQnw0nxhyeIXGxpT089lVxxb
SObE15TfFn3hOsIc47BySAI1MXv/uFR6W1NQKbI9icNhRXkVe0qhlIg3urid3u78Hra9NlXN8Xav
0+4QOlEhgiBzp6+b7zpcbL4wJKcinsuW75vW2A9NRHzGQjhuGszUwzE7vgmcME2itcWPVxOnyJt3
PLUnXSSIHUXzJC4WL60Lbk6J+iNmfbO+T6UvYcNMN1uxqu5854atJImgwaA0Fta6uHn6pYlD0CUk
e4yRS6ZH6Sd6Yz7Ub8C5zCsCg088t/AI3xP8QthWH/oZo8T4RnlPPUYo8GUiGsiXza6w8OZF8RwC
jEzd9NqaIEU17Sql0n6QsbAE4itAjFfGW1Po+HQ4U9yDmym2fqbvQAN3rx9d8kFvg9/Jf/C/jXqe
y87kmGvIEeDELfy5DkfCP+WaOrDZBGlvryt1P8WHcqKVpuMNZmW47doI8wM6t47rnxftO6IPuI0U
JzVPyApLQTLmAwIkoy2k0OhUh0Sbo6Cq7Rnf/JkstzScyY6EJFRWNg/pksNjfVwL7X+8OsSQBHSM
L8tIXC3a7gjPQXimszlIRXXm3QrNgsP6iEGNYfIKmZe1n3rfpVKv1IYZYo9r8Ha64Jk1fpy5jx8W
INpuYB4wMheKSATFtSwERfhhmpKA54OSTx1J3E10jC9J9uLiyvFxBj5wu7PRlmablLokCQ2nMabe
QWp7zrK8IhhnmborzntbW/aa5w+l12nQrwmYTKNqDs4RM3Nf+ZBkkW6qXWgrJail6IVFcV5Pv3d6
dShExW5cYxVBlRN/ADA9tlhmxGJwoE+PBAIlj7/uOuCAUHUJuomggG83fVp1bXG/Nmi4ts914VsW
Qe7CnKwMrat9dRlpsv1Rf3Fj7++PwN3r7doGBFUbNATNrLap5i5lOnaFRfG5u/WgSdiC2zIlswJW
qfEIglyzQqJYoC3bvLcEZvL41QOF01Eje0XuhiCmPmvBCA8cpGBGScGlHRrJwhNwtdgSWp7Y5cH6
ocURBgk5Ik+fZtk7kKwluAtJj9ADhuL727En2IkonNDnHyNn+5TCLWBBEYt5sJV5XfS0gkr+RYiF
qd11MHD6btxzCmYsH7D0eia72HC5JL79XN3QTeJqc6935h77DIcmZf0jWnonejueGpNpBlbuERpC
VsLrpVdgtJBuJ2Ly3NT2Kh+5jbCqzWoQRkFKVh7VtgKi5MZbtfhwpRLDaYRFLhwb5u+8ZM/FcfYT
CDXiP21dIZNluoC4zFiNLsugoPRXHI/MyuGPuRhJOsC1ZPrs7MCQx4WbBoQCtoWlAYqid9RJOqwT
6ZriNIuHPMKd6yT+BA6mI2LEIv9BNhwAHQyhKStKtBs+lwY8C3Zw8jYpkk+qSZmjdLVux1+fa889
PdCV0W1WLUvsjZncUfzzKEtpinCehOFJVsK6NYITPEwCzBG6SjyDrD+sHIR7hbv7g0iwxaSPow7t
2sKcLSLJcr6rWcPH7EcRmHicccPHK/GNu8jgnYKxgQgkz56Rr0WWNzULXKYiKMnhFt45vgBoUgjE
ZuuGKD3R0YECjTXaa3+yqIkzzmMA+sYssBhzNyrpXFO3jXQbamqY/UhW0eG8OVDg7LKU/CzR4vGP
51OZy2owDP03VmHZ6DHytnYfs4VOIXvDIiUAZpbi981Mymy8c1MfqTXF5qy47AELWOdSILsfdBCl
2Oln/nzvbr78Bo4FfygzqLdUnYesG/jCCvCfm2MQ/GxvPx6MmpubPVVG04jlu2tOpVtSjF1CBIiQ
c4L47neeL81YxzddnZtXOQbLakvGRJNFFgi8hVi2rMoMB/gBdlAvuvK8HlzANS7JqFrpFjqCnGyt
qplC2hzXPY1VJxYPa7AnwmCkj+PWQhTBRqhUCvJyr5gmYnzJEG2FwfwZ+VzDqvivr7Q+woqN2Awj
uvDATRWCnsIfv3kO7sZbJdv/+V0cwfFJQ9knePgxY4+ZWUzVtQE6h9az3KwZ2M0Gk8yFvJCHK01h
3k8Zem9rTWFa6AzijamDVZUaDY5O6MKRlC5mREVxXoS5N32cx5c2nXnA9QgfBafgG/zDR6YElUBR
la8rnn9l8W1RNB9q7/L/c/qY13RhAVC2a6yQ6xrPOwyyin2d2fTgPYbFfeqtzMXI+oC60DWNM+Lm
/MIdWBuOfW3ol4m5cNdQUuURrFFeScgs0vhSSqcoAi8skOx5yuZXZSylbpB8uLWk/seNUL9gqVzV
cXeCqoRH5PwIsqtnCECZaQHA+8JrYOF84O2/Hu/Q/PAsZgPDVz1zbHyCyJ63VGnQWSFXg8LxlIcB
wOfoX9oB1Gi9ghPjnbBJiEjYVCye0gNN+VU0CYiuhN2iXja67VZkjAcsNeFEDfKcr3H8rvTD7cNh
c03WtaIREuSUE/ARNSACHiaej1XNzJQegfmohEqUqzYUZWyBlAwYmCdRYWhdiAAceCTpDiv0g/zy
yjDkVwWif5AkndTY2P6oZpo/IZ1/wFIpFWm6Am4gaAw/585wIez5rY0+xlawCV4M43eawG3yzIXZ
QdFoL+zSnPNS6VBI68tT3LUfFrKIoPKyUCtkF2xdI963xLCRi2GNcDKSjR+KE/0OaNFQzxyAPGpG
hgtY8oCk5CV5ySSGKuL6G5JK8UTylNhY/OzulQisd3qLvriNXKnZPFXqgR5xJ4PJamVOCnZ2LvZB
5VYkLJdzLG79h+K3Gjj1Lr4LfU79W0NjBV8+HcMBqoc9jkFsCyuzTygdnr4HVYrZXHVyIPZm6shN
wN4cdl8Iosh4ikuBrIxRDvyXsIxQ9tmpiYEpDVE0zOJVvRZv0PXeRxda2DxH/+isg4gy/oKlj6uI
7PzoWqauOWkBlXzSSush/yhaJud7RHerhaR4Ke3f9TB95B+L5cHL30yeSyGdC4W55Xsql2DGmBC1
wuGsLBr8+jx+TgFTLGEtdJn8zWGVoS4cZEqCzEGbAWqt9StgjwzRyzipSab/gEHmaUuywnI+KgqX
YkgIEE1TG9tevpbYBua/FN1Ui6zS3T4uqJ1QNHcvbS5G886U7kkcO72pjp0fPS7oM8t6KjMQda9r
kP9yTMq7v9MrTtP/DsFhMy9ZNxsP6zWt1INeiyYCTcBMQV6bUJWz77Q7tiANFZQuU/YO0N45QKUc
i49gQmN4c31XII2wSa+R1NDb9Sj8uFp8XvWYVvLPJKTYTPepTB6WKKu19mFHVCdDT8kPjBRSM9Lj
PumzjuFBv2nJGMEGMp0NeZdYcSv43XfR7RazEmdS4ygm2mu+UVnFFbPfgUXJZaot21ASCSNqi8zH
jf8WTTLm8y7P7joPsCkiuGJEOUOZVF/GeclS3c8A50YOGIXf9bp9zkFvEzzH70E7cCITuS1pmysB
QPZ4u8SK77ZpTlDiEz2KY4x0+fjzq/VM3bV3TYnZyydo+ZuxuSckNIXKL0uMyCI6TulMUoYlswma
H4QSHmTQG9gqDgE21NG4QlebCANgl/IR+9nu8ymvvbJqQyy/dbYYpWjQ2NBV8PRHCIUeyKkJPyWF
27dMcu6SvvBHQWAofgFbr3JtKYj3uquB3un42fCHyVCcAcxzTXI595oyWCpxkrGUOMvC6mVggW/w
nM/0bqgRqMzDZPvcQWzaJEl9WhAz+rm+C4Ql0JKH5V+EP9dIqu6krIX9cdkX6NVAko0yFvul2XkU
5AN7fh7SrMsQTZyzoCRVWyFBTVhBayfJ5ArEkd6RPz/Oug/oxK3akV+eyfemuCJ00C/zFdfH0mzi
oOMicWbvpUYEHJc/i3LdsFSYW5E6wjAxvb+YhyrUdPgZggxtqPQJohBhiLWs/xQeWaPp6FeMjdjh
HJGsPgEl2/CzaS9VvU7rgDTfavurIWaCJcqX83PTskU10AYzmfDimVTV64yeezZEe2bEjGTMgg+K
kDrN6W6LPWycrYL434WVQRd4wUOWsOUWMWjlHRj/KGNnMGcS7M7K/xxelEoeaH9dvbQ/yUokUdY2
SzjqKY1vTBESXrk+YDnNTju9wdALYWHEX55j9+VYbdoRHBCvf+1zsWpjCZWwy0wN4gjCgMg8AlD0
UqS9s88K13z7dM6TkmATbCuzNdgN0AvSHZBd/8D0ZZsNjdh0M2Y+0AqQf1sxQJX2uvdl2JyKQx0N
pCqGHW2RfGVJ86NIwShLV1g3LdtK+WF+A6V5yygb88Mt2PBcbseHJSVlh3nnGCVPg/oiwc4t/goW
9jwcgxXf11UfYeKS7EPv/aQUMHPwz5FhlFjLLiYAxHsfELLxZR/a36QkDtRE/rD5MGPyqnjZ5eMu
PHHSH2MfK8QLa7GRBjDDzz2aHDFcLUVUnAXGulT/IuWfqIcoi76EjngBtNGSnD82SHTz+EMfq6oj
hK79c9fouR9mBUAaHTrISpJy4azcgG4cutE/OrwSfkH9mCqbC5aaD3Uz6sfHw/fcxcaKhd4i/0Qp
81XoZkft0hGQk8Ney8tlo1R0BWM8jOy2ZgGftvwpi3Klhiqw43KkfnN+/R7gnpmSmANce1hKMnEc
9O6VzrLtK+FUhcfUvZ0t61CvGT2uRPppSTIlRaj10oUg6UiT9//ekBULS7AVPobNY9dHF8eh6f+q
PPI4AxjYwPWZSyXGSmxyeZ+yoDEJlNj2ZilglwRU9xWLwP8VaplN5b0ImEy1MZYiiMantjFecZUC
MdA/kpu4vv+MnxDggsh2Om/GXxq9PKiMggr4SyUyiB+I1kbZQxlmjEtst8EFDEJLAr4mgl6k0f5p
Bwtv/KTWINj2TNcmNQZYywFT2kiZX7ba5wt1ZYfBDKwvc5EsPRMv4TXl5CXD6NU95owiQjkPT109
GtTejAJKu6yvsEBfxXosgYfEoZVIsbKI6Rz/Z7eU5+hNcoentJw+wdBctdTyXfyBtZZ4eGdWhYuh
3hGbZYdi+YI1dxfdTQPueQRG0z8b/ANsj8yYtyVQpUVtsdHzMX3cUvAQzF6NavwlAcm/x9TKu+pj
NI2ihx1BuMKKnd6rCBK6EPnoidVZfeS+/LOWjlk30jPHDsr35Qdjzk9xCXCfOitH3YpV+hKIXRqf
yG6AjII8C7pPHh7ZDZjMkVsxBDEUstXPuuYrkLEa7RFZvDndAXL/utQ6o/FIbpwSHaK1VJwtEF10
52+s0B3aqC3lch1xXvW3MEW92K0Ju7W6vgQ3+PmctHQCwXp9JQiZAuuh79OMM8VqMLZS9LIzkRio
daviOH5PTOVbKtiaLb6x2EZvWj6+nc55Q4id6LW6DhVgEiMYiWhi2XEDrbQV16+uNkvv74Ctm85P
6nj4uhlXHcrxXOx0P3FZYwO8W6ytqM7UPWBWXhPmKDOal/N0Lye4TpHwXD4XWIK/PNyQcVqBPwH1
WDFzssuSeKO9MjvZN28N+O/NTbY9B3+gYPHMHGASarcxgF9VzVnng4ardiNGSrKg044Xi4nFumZs
vc41l/oL2tv2KPkeLfeee30bo/MXyNqMtX8fliCN+oUM3Dp2ZsXay+HSJFrcJLQIKKDk/Ua9PB6m
p7VKC+Op7EGBz+jAifouxSh7W+a0mo+9vWUhbQYpMGyLS4XSjeju0pVYQwknbqa4okYc3+ZENq3g
u98Ft/lyu0ExgK4PQdVzHtassz/2FWK6RmqR8ETS74ZzYHFA+n4mt2quGLpXvVd90vveqO6FxZQL
u7kdiP1mVcrxS32VWZsX+cUrcTvJ35hv0/tFklRHzmci6aSeXmnEqgiUIH8E5yZOq3NNkR2KE9t4
++gdSYExzX7hQD2UpdHhAKB1TeEMzPYUFabosHAZcP5WqPkqCqmyw7/E2579bMQDH/nasZPNWljR
58xA/sXYAeXUfGm0ynl7pbh632/KVBH5tdxJdibEfeBw6R2s+TW3xEcQUOAZZftmgSov8gyMWq+Y
/lXCLABrxNCa4fCR5lLOn1SV+CcV7kklhbVOlwvloLA9ULHSXfq/yoH9vBFLIqNi2MDuMcRWsAUD
1qrsc8owuDjI9C86e06xuTocG8et9qrPVKyC5AAl7S4auf4CV1/DpGhE9Tzp4d+xk9klMhY0fYbf
vBon7Suo3H0hGITkm9q7i5qBFbquJHJiSDlWV0cxSUnM6wKb5HbM8fdbEzhFXpTdwoMjbE7PFNcy
D/yBJP1KwbWmJ/+p+s+X/ka3ndPX38i0NUqpIrwMyRM3ks+FaknJpCZ5vXcF26NALIT2hHQ+q1nN
aztZS7ZpQsNUN1gurpx3xM2bd6v5ULvgBdzTr8KsP+a+Y0CIc2YbQJJlQnEfM5ZjfZcSpL5h9VOT
82/j+zUMGlzOWQuAYxqjfOBCAW2lCZq3lvXNwrebnih1bdVdrjSuwz/X88lsrPa+2ZVKaWLdp2cD
oFgvdFTCpEsSe0VdJ8nKVf1GsNdfLzl6nyooIgU2bIA+fixiuvVTa3oHLIYDrUshRr2dZolxm5t9
gUHbdv3ZPjDZMJbTIsfGq5AiSQLcEBcB2Ep8Wv5Hf8T7rYCw4EiFA4dHfTBOjfkL7cE5+HKf3hAI
FJHFQyu/eSox2nYfzdQUEvXJb0BCqg32mozl8jSyrCzhZcGsUnCr6WcTzLeFqcHKQfnlwczt7F/v
OuZtmnSZrQB4pqDhIQ+FpOpbrgrvzhOgcz+8uWzkHPwMSV0AgRhbznf8QST0ICo2GVBEQAdmB/oB
NJbWeWerObVIK4LJ2Qj/Rq4Hur9gu/0uUsHZuW8l2Ht35bUnIicBf5Mc43m12eD3re6H1Oflq+y2
IFWuYXXI5dslGF9l0v9qxNeEeAJ6ukBdjW9go/TtHW3m4zEHuWcoUGyuZGkSBEdiDRPSfEPV71v/
riq70gyerxpuNXr9gMDgrWzOLcezx+ctCXRw9kDwjeo7YbY9wdIn9UYmQkNy9CJPBiZi22YbAUZ/
8sIJ98HP5W91q+zW7weZDug6nAcYZVS+zCYEqAYwTnZrsO4gjzs9h17uh+U2m6WyDAPIXAVpQXh2
iCcfUxSddtMIRUO25Vw/gwRFZrV0cfY5fCh7uj55VnLxRTtNfNFOrZ7GlHhebwS9CPmsUnVFtaGH
ppGi2Vb3ObPgqcp7uxXCcoHQoaW4rYrCKDZUfuljfxSJdWGizY/E/Qb6bbyKK1M/ouwIq7iDW5h8
jEwBXVQnuI9aDAj1QX7rcUVxlhlo+Nirh2ZTMSLT8p/vF7eNwRAM1uT823ZTWudmKUkanJaE/FiY
CXH+OpBMmXiEWHR5FkYdJy3HPkWR+GDpVU1ASQqDEMAfjO9MFLxksyXTk+crcVNXG0N7VTHN7vbq
ZSjyKldgHUfuiklgkd7NElpLIevNwxBgOKa9sADQfaKylBZ1TYeq8mQvVgQbnbl/dYtB0iOcG/2N
ewI7Gg1FcMryScfsxXBAaT9Gd1hEYu99oOuRXuQ0UfDzVAHnI4NQUg81Wyk31iBE4FmB4h10xZ1W
gTOsfG/BNtANcFxVWpGEt/OVZmR7R0iGSskWVQ3bjgrYIgVXQhCjGY9eZX89nGbILgZctpNadZRZ
Bly/GXbRJ1u5NMnjIiyQflpaO/Ihi5+cZRJOqJ25WFPXJMuoYEiQUUlzVspb6yaRvuTfYlW05a/P
SSBGjWGwVd6uzHCqVCjaRy/INASNLFfwxK1gO7tpCVwKOBHR4S3AIPOBg3Bll0ovjB07f0oWsjYt
P6KYYUpzXAhFlTdZcIM4DesP5BGoMF1pQYvdz+5SYXvZ/DFBsiDHdJ0PzqjYO5rgEJcfLU2WB6/i
IZeKq6TSbiRZWlgCWD5ZWxuH/Z72Ez2MwjqMkEf7zffsz3Mbj5s7GXn9nvlOFs+v7H6xOTLpHPSg
kc+x7NsC1YkcVz9QA0OHpqkv7kMqA7k1JZjTsTtmFdq4gbswSl20p6xno2oga39FaYG/BfNtASOg
FbEfScuaLmEIEFv1ZaiAGmEsR/qRwzGzhJKCxfgt+CkX/uOFdkGlj1mjioDUV7smjj/WTfs0XOcw
IiSApsVtqjdeBfzj3EZw3Srt49f3aYEnBxB+sYeUAGT+C9nUFKxqiOxdoGCBZXUQ0ZacTqEJ1l+4
UBg634uJ+9qqBzOFZQ1W1ouNwEPtVFK/h9YQctZRpUIXuKgMVcVw1U3zJ6p1Zp5BhNVayjMDk9Ux
tEyaHu4zwrMystkDyHcv4wihYoJjH71MpdFsIGxG3Nvi2pqZqm3l02TDv9iu/XKbwZ7m6c4P8H78
870IWO4Rj+R5AZqvrisBEcTphO71ubudVi2g11NOSDtcUu0vaTf7B4xjs61pBy3h8LIYZtyHTv23
obATvbd/mY+j/B66KDADVn/fUwEtlrbsjeaMwkNNUWGBPmgdSiOymMsbmmzs8nQ3awrZwVBUxtte
MKwpvz78/028MDThiLt+Q3Kv0mTPDQHu6G3uOJ+KRevyemBOeKV/W0vPuEbHyMaA43M73stfi7Ni
9NA82XHQaw5cbqL1PvaYgd/+xrMg59CEqeXA1FAWevEJZkKgzPgR+DdJLoC6ucHnmsLewrX1tmou
oAVyDCvgmh1rFku2XRlGZc9pHN3wImtD6nYhtGBoTTnYuUmtXv4wE+iyf7g/WWyJ0TgxKToQo7j0
B9pbuvc/bsS0ccWEAk2m+yMZkOsnvXYvZNRnTf9LACpFCQ0ctfDMlM51Zg13HbrUmjZIu2GmALgE
VAbrgzKjPVMcrL9N0N7RPYuKWQ2E01BWe8/J5/E/eDEjIS/FYdCcbRIxu3jAYH30HRfts9cPN4Pd
YnVf4LAQUmrIYM9NQMSJU4IygbcMvw4j51jgALWmBQA3zQqfgybSlpeNOj423U5x+UuMPrgxhVMW
h7b8Gk88LBs16EYkxQyVUMEad0RXreuBy8AjIlAb+giTt3Sal50FM09oo+WmpuyzZG1J7w1NIKMQ
MGRqyseQhvaB4kuqVcno26Jhrgc0cmkE6cwzFNN+elHRZRYznMnm8LeEcvYllTLeKS/WE+YOifPh
844fqCJicd1coSAZROQlu7DKMg3tTnwbQVEk18QB+2aeRA08/g91e1Je2DR8bSoBT1YnZxswrVaJ
VW7vjd5HFqXR8y5WrKhfubgN/K0cf3reJ9Zzg7f1hbZgH3rp4NhMxmSfndOtrqLusXHq/nKFJnzY
p4BGUtL1jflNUay9iMrJiPbS52OdNNdzsQxDKxRJPAkoRQNB4VL2UoyHQLUjvQ4dfvM04NC0Xngo
aYQaJrpBywR3QUCcsjAlsOBxPw46GQVndItH3rKEupA8yx6/XSVu1515rU5DwmEBUaUuDJCV7xn4
5O1geM3uB7U+jK+EQbueZ4wMauMPcepL+tjzXOw4I/+1TiJzRlrpfNleztYxFmjuVbPDKI9dkW61
ggfzGw4fApaFq6EuDdNGxTVaxgQnqEBNQw7QI5lcBrA6MajkpoojGSK+nGw8B/wuNJ+9OA23LHzq
9TSxwkRm0AkRfEbF0Z4nUxMXpeZhOwFWPOeNKv/trRMKg23Nrk2k2T0dvIqLXjAD+fAtbFkvBX9c
WSkMr25lG9XI5nV7wsRhAqP3L33GtwXuxnk+hLDrknU8yo9pTgUVuES47GL9GRzYwHIwuqTJJnPl
CAAl+4xPOJzSpCjqO3fI8t17pr0g0v5h6GQr8Qc4da8+d8wd86NQeakTWxdfAjaJoFKPQ3au2YcJ
czQ1qUwuKUh2ZptWRWuu0aWHvmovCkoE+8wDfCtw93Dl7Rv5MyimNbtiqkJ+UN0DS4MRwRBlmjHC
w8q73U734Icj2tZXKRA++Q6vslj6yICIWZvE9UIgbzIpIN7IV6EFDE/3KIDchtuT031sr+OvgIF9
fm3BLNec94FErB9Iu+g8ewxWzttRapb0/2Ht9hLNVT/PTjaUelxcvtt0LIHR7a6oVwAyLO4PfksA
AD5M+IcUUjeQlxhZBf1pXYiAbESb0DtgbPOqDk4KW1OUfUitDIvFMFzs+CGUCKPRi0C6UI8LhL95
cAy5pXkvIQJHsUnEHPoK4Of9hGFKDrNtszTH5S6YGQcJ3yl2i9+q/UnsvBUxKYvX5pabrFv0ctv/
pwNMPgZh99Lw2VRqaFI1SP+gODsgMA6TmolPALYe+fqfRls69u0nnx1MFSFTtJkUYOr+KRjusP8h
CPyQ6aRG8avG7Pw+vrZCjzEA6AYJ+KWq2rq2Xg1O7x7ziPemz5jTr69v3qLTtgyaqUgzM8o9qstx
5T+aTN0KGfKZd8s5z5LdHC2nmijDeriaRgqjk+M/NdncD1SPbSkEmr1QLtW0+a2VgRT/aDir1+9j
flFAqyyXnYACn4b8kpI2WxlS0uPZsT8objYA9lfFSDCyhpRA0bfbhRmtcaYuaLEv7XV7zkwy/NWx
eVneiAp56xlXCwVhYSDGhxOQNDcoiTKGMS1QI+kgpYCWoz4ABIGoxYhRnhVOGOBDOFXhbOQSRDBp
pf08Eiwuwwatg4QJoR3AwsFYrqR5f9yxGEasHwNZ6X7hPf4UhBU48ylGNPFu+6JdgjxK8ruJZ2bR
49fqgN4BcM2Dwu3D15qZhBOROH/HoVgyHLjsNmhwNBzmKaLEqb7di+rFSMd/66ZHxjPRd7ofNlly
4FsfQZmlsIGEdZc4VptGxNZYIff4jnPHdfKnwvZt64ZwdUVzrQxD/KaWMdHIzdMml83wN3S1URIN
3zTEeoxLfrWj7Ra4lXDjnsY2X+JjgnEGbB92x9RaysJ6PE+IdDDh8IgEEm8ebONds1BN3Ap8uu5W
d2Q3HxDToGqZkm/bN0ClxDlzy6PBMnFMc/QOx3p7HZgMmuIPpOpsxejU/NUV1LeCO63dNetfKzel
RroyfnadEla/drtTKG5H/ukBmcg6m/Tc1JsbSKS/U9kt4tpnONQU0d5OQAaVT6X8PjzuZj3Z2naD
z+r0NGF6SiQ+afPWXwXOXvTYOxqJJ+sgXU7NLdYRs1ionkmJwSxlzEJ1EnDTq6UWN5lPTjAG4hzB
MnFkR73bTs/jf7Xq1Ymj8WlAuzXansX8nsZ0P4oBLM2SA33iQQFG+nlQm6rKFyMMMhW9qiCMDwz/
ctot7SpQvJuBMLApy8OS9AqGZoGqWYuffdqsCl70ot4AjlO1INaGcxIXKyAFt7G5eo2XLnJAZvcf
YnR4i9rwU6Bhh/nUwE0rn8y+FvzF9h0eBAP/enPwVDq0RoI4WCnXclhtyNf0zlH5DK4GmHwtgfQ5
jE/6q+Rsi/SDhgOPMhh2NhO/qju8h8Ht7/1aIK6E1FGQpsT4/DCQF5E7mpvRQ6tICsmaz2bBgeMu
3n3suzIpsZ/To45gfdCxyhv2C5mrEIfQwvZjGr4Z03t3uCwudosHoI4I6Jm+kVmTcO3hdMRFeAuA
W+qiyGOQhTgOMdFs0BH/HS1YbG1sHvDVeVYO6fOmVk35RFGPOIrV/+c6N0tdVkWlq2OiKIV2k1Wl
KR78U82AOLSafOVfa6IfYsEpdrM9MfVrQ+JAZ5cJgPDdaeN/b1tcpNbHjUJ+mcfcJ/C9hDK24JB+
ZWtcdsN2c4j4GL1jCP4UOiYt/GLAYfJONBSVN5oMUzhRM/gwCSHOAv1pRdgWhLLaOOztIcScCIlY
bjcQP5bDgl5LlSRMdVhsPdx96OR4dv478Hq+8/T/GUCx89GAUKnvnl5uQlpw3Ec0XTczRg7Z+O+j
VIxwovJmVmkMgz+7bQ4VwHTm2Swnu412SWkUhAE73pppBfjqm4JhLW6j0EnXa6lUpYMN6/kKGpV8
Q7JSRa3UtbT1nVpjdoH0+RX1d+SOr5Bn+nuyvhqI0O/lKoGVFX+xA+7oDahTYb1Y7413kuh4qdsT
2wRHLmKe/0FE4lyHbR1BjkS6uYS3obN0o4ZiLhMbQvL4mY+Ue0iw5mBrTM5kjdNCaOVwcn5SD0eo
183mBQPxQn7zK1RZ01tKmqpX2wpu+u1YtzUVx9s+Cf/g/WbOdP1sHmP0ixLchWIXWk54ynfWyEwj
AYoHzwqNMEjBBIkrNZtpH/xqsdSVgH+CE8GjLbRGsp4meulntiF5mqX5Tvc2gaZfOvbyXhZ26NhR
HeOogb8669AtuiziwDHjMTizdI3Zm7+oQOACjQ/UUmQNgTB4M0zoQHfE6ZcBPVBHcuQahIwYx8gF
/8fXH6H48QVGgWZZAfOlviZ7GYk0oClfp5YNlj8h3akQQgfHbcG5YnYrg0uDR94Hd6iWG8XTwLT+
s59KOeSiCei8CZJa7LWY+s/YUNq/lhNohVo/HOFGpj7LsWkdP9EAVkfYwvgTiAH8j6gIo6nEXd7q
lMTR9ivBkGRtml5HM2pRMYVyr+QOsx7IqbNZjU+cYZmi/FXcSiP6uDMy0LaRAZwTpLqsoiqZlBSe
G4pORRelqaBCV8yZlOIzaE3gdkWbrSQOlEYCetszCUbDadiWl6bhm9slS0g7T8wJjp4dVZkbA1na
QzZEdFH8f6TbAOb2DRO1L/pL1zQBu6tMPIJWlfnzvfnOozGFTmP59GmvZ1KcuIIkcJtWKYtwtaDS
b78Ysd7BFtebwys0hPhbW/YL8q4VWdKMbvgCra02roJwH8lRveEyu1Fl62OhHAqJKY5zK3ngxYeZ
o1xTkMRG3Ti9vNXhIcReeMJnJ8AXLDeNbkORPKXVUwUiJIMo72vLmjRZXB+cpojB2oockUUPfVXM
xnGFw2HM74GgpAlf0bqZiuUYeKVzIisNKc0QGWNvvF2zb3c44yHWqKfhBFF4Ul2n3VVFLgMd4U1S
ny0ldSDLTFN0EjCvNizyiKJ/uGvIxn2cecqoHkxWMXQwlX4NGvkimde0d4eaubobZIxL8VJYknPu
kkNENaJl/GaEcpIHnsPy2WscW9MrgULgxhW2Bv9F/mYHQw4hnu9zjfGuhCMGZ5VOghZ8bSRq7944
1oUoCkivdRnpFfp2SSpelMs1EHy0ZTPFJL0xSQmkXq5YVVZDzqh/jMqYIffGM2GGdSIyvgVgw4WB
+EeEClwUF4ysAPvUt6bFyIWbF0rmF7gB1dAow6jTWeR7MzF0Ib7KmvDWz3KpRleD0tcahQsiwIdV
WFQlJsEdykv98xTKRZs2otj2hFIkyJCnFQoKi33irwNPeXUzCyVcHQQ4VrgSJpeKjPy63Z/03YWb
p6YsSvjNNfINd+d+k36PuEHhuKRJrKQ4jEv67v2CPxr+rjQtUInHHHtdqSmeeWoyhTspRqv2vAPG
b5SQQ33RapELI6U20yZOLOLLsbEufDb+WDkyNwBetPcPnRTiSymz7NlqNQkd3tauptR4yUkm1bUm
ieV7NT7lizT/cAuh2Z1A8rm2JwNvrm2RpXn9A0O2udKxrlVaGVUSDI36oKAQZy85o0mHSnTrg8/C
PCZ/VQyAGqIi2YaH8WQ06myA/Wpjn7ZFafjfzb0PUh2wTZoUX1cYBirqA0cPxEXUm/GYa3TCw6Ev
OdiAfMDFUlelfrj3tscUieAC28b/LjsrWUFhYXokI8yVvYiAbMcqm2IGHF00V7cKRGQwy2h5uPvt
BDVvwAi0ioYd5UL1hZ4f8FcbNrtnhpiq3RG17qWsIkPS+tgbiYOzwwjjL28+EWtAtPOE+7Q9Z5na
5lr2tf+9wedZ0FIfUiSN+ReIJ9cKaGSlj9y8J2kCnW+qXFfKSekMs+y9/KdKkWttVbt9gh1poEZL
hnvgBX1/qSmkdS3Lfexj1Qhgfwrtjw39I5GO91reR7YgVRC8guLKFdq0no413kgomHNLuDmfNgrb
Sv08dpUFaAjp9b0Tk3svyHKsKRGu6Cpg/jpgQoP0lBDSaoEAuywByVsiVh8sQlxP/wEK9hg7UDhh
BPCKHPjmhVeEFSo9lbgQx6TpCLUrZjTBAJE7j1bU1zHzw9UqupJ5dDSq9YbQdfkWbpEN/bYRI1QA
cTB1xzbDT5XbH9lg34YH/INJMERxW8Yd9j5PV3Ut5Y0bwyAvWPhPRp5cytMb+99127Dj74P8NmIU
cLKA+f5jveh1iuhw1WAdpCLbLSEjKOZM0cIBzirmzSQmnehaurVPcMoDgf0ZMZOC8UxmS4aE7FVp
ACtEJ8SM7ExDulYuDbhRBrqT9NpCM6kZljtXlsL4upnqWN4CJg20wS7XBWnH8U4hy5MIGA4ijU0I
M2y5jDVhLDdVZTQDuGFYNeSqVxr/TQVNPxOkEz1H64nYLIjoI6PRMbjUMmFTBESSOGZODxeRG9WM
a3BMinBI5y2zXX//6bg5l1ESwFTM2QldrbA8Dn1AYtl1YbhVdai2Fxve6KCa9vkO3MpRGfHl1oan
pLt0fX5IYB/fob7+zRFSL9l5VlySOQtqiO1TcqQVhQ9cIGEahFk263Su8dDIS+lqiIcgyKGNCWrk
puM/489HRbWS8C994upKzGLwCpKcJ4MXAsIABRXRt73HOjHcSGkPjiAU78Wd6m0yQEftWszgU8hv
2wMwg5ZlhlgI9YhpWlBw6uGbo34ftTFDr11dCTSxVzX1H2K+yVOu7euZUqTBCHH0HxKu9n3RfHp5
gYX7VJa7A4H7uHELa8etv+lOCuWTDkBe/7PFbmcZgr5i8xQlux4NUk77YndiRhOnMtOf3h01DwPk
zDGRHXuWVN1WWJDf/q8piYvV3MJWztyJ/dmmcos+uDmNYbndMbXSKO0Yr7a9IdmXJD+R24YI1Q3t
KNozvlZeiBOCrv06dwMNtl5WbKU9QxLh4h0O2k1nnvPqc3/AMFDXnRvOHAUwJEiuqi2CEMgrJQFm
jyK326MrpEbnnGAGr4NMATgP+19dJI/ShqKnIPHAbrocyXEv1CPMyOlVfqxNFvaBpCWZo5RZT6FA
lpkdM8qXUj33ykoWOyb7vOWH2aiHK9pWep7ZTje8eVni88J08Bua0NPy10rChYkbyIeLE3Gs0EUu
cJONiLhAJyy88HvjTmZzwDG0keRQeNOjvJsjM3ZC/a35+iDg4H8CXDgkh//gV8xEUXkXrtcHIxsp
9g200lhopJPohBKV6viKQNF54b7Kai2bOulhRSKeZJZwxkT6Tu+1zra/9VVLftHbuz3iPxa5Wnu6
2rnKnfLSndwpFT1hnst8f//eDm4N+4tnFnDXCH9Y8uv/UaLRluu4nteSi3yD+8QJzPUl87IcaEDl
P8pTz3DEtWRQxYJBvyub+EFqrH/X8maVEstEsN8xQ+Zk8fnxE5w0udOhZ/OYkT3jDPoeYzGelTKD
exrmm5OIVUTDaMCZJ9UBG4HxNcYm5zkKhnZx9JV47EpOPRsNeYKzvne65wvmsfdgLUb1ZUdv+XqC
IbH3Dg6S0hpejUotD9jp+iiCnLifbzQHiBr8dcOdkbuhqSlUxe9d5KyYVB88dClDbFuZj9UvVd0O
qBqFdC2BZFu82Y3J6OcapjgW5xcdbDiwl+9bZljrA/eebjz8DnLc/i+HQUiloixzRfDRozSIk/YP
kurwKP5Sxcpg2ziAt03j6+Ry+HJueDA56/i03TtsaY24mSDtzmBPgB0vTpODwCVytQXwL+sGMZYb
ci1ct5erQLnnHLHQdvQclcaBa5wZXEIPRP9rYbOo6Y8pCnV6Ldlol0QyxWvzpMDfzyV0SM6oxArd
w1MznHuR9YxjRkl6NrvT88o/GL9AwfGgNymN/ahye8eUeZWpkMfKcODwrRwb+r9GpaoSvt+EejlX
NJQXjzSotBgh/KcjwNZz/AZWVaqOQkEy1jXKoh6r1/PPrSxpYQpAi+haivYF0m0RkxBXriPgMrVB
yUKnP0vWfOrhn431V3o0rVvDW+mT+uuRMwzX2f5fnZRsoRzJC+FJJ7mzqQ40aQx6QxdNueJ/oFP3
OxvR//3v7CHnda79wYK1AKPpkwT0VlXojGKO3IoRcIC8ZjlDexfP2U8NUAxDXhAtZFVAExCvCCU/
NDu1A2vL5oMDLf+EsHfGJWeUfDbJG1wzQaJxvq3f7IXszqACovmZeHlIC2pPNUQCa3YMGTPg9F8H
SriuYxi0W8afh7NCXQsrVFa+drDCP1Nzq+4imstwm+HhKqN0gKs+GsXgpIfXMUVatTJo/sqGhPmw
NekHuFVh/KWj8QgKjdaJTpD15onjqgYpl7ysoV74pDBXLLVhdlK9UJz4gUx6peBbGfrxXoSfLNzB
M6vLkyIl6B7ENEtfR3G1QwSwJBazsH6rdVuoZMzLHQekWV1UCDy14gNFnUVpdp61V7ND81ayQGFB
zn+5a43iCa7oKf0G1B96SMxVBm8tX0aidsTDgPgXC87DWRwwzVqsumQpq+Le5mZD2CXF5co2Au7l
rspQnyXCuGq65OM49HyoUGRUMVlWdoL6bssqdkRgKa3VHWiR4oBjoKMR6FPcRiHgwlaByP3kBpyX
m9+lpa6EpLIWMqhdXUJBkSsGbNZSKKOE1vxyiinOiuDAdjhJs9JR4qU97BQksGwtRnbGjRMV2oJE
H/BBZqkM8kV0hUziCI1noR/bArD19M2rAUWeCrgOk8/GDlFKi2VPdlszRFw/xWaEseMjvN67d2sW
YoNb9/u/ZKDqdzc3oyJjFtzccfslW10Q6IUYYJdnBbfuaENDdRBKBBQHhe/uLrZCkgaN8fUFCX2G
B81YDEylR7Z7jBARCU9KQWYrdXUit7sP5P/uFjoOpF3B/CtjAieObX1+0xA2d8IcZR/QM6S7Peux
RsAva+GVc7r+KDXMxP+hzewksdr86ZnmwTjy9wTW8dl5a/Vhkw6xcZekuky3zhj3KTgmttE7YXFL
f8Oa2MjO8vgr1tVIE5kM7mfDYwGwgADuyuuOEHNY6Njnbk7kL0IqCGrKqZnn7RzjwsKhPCGt8gnX
jjtp0uxYgAxAI8FRh1VrkCbyfw5jFvh5G5sdwKV0abuH4oDtdT9HkE4TTmLeXZ2K8mGFSxvBTWGf
FRZQC8aya8YolHEnl6pjthVzXGf2bgB4gkajPQvC6nRBLXHHcoFCwTfMGRKNpjxGuSg8L3JkVqw7
wN8e0GtwIlsv9yNXMTs6aCWeVJ2Q33Wx+ma1Zfg4MWq7qAZ8w22LEDYMnjrmSl+6xNKiLWolxeEv
cblqpTwiH5Ai8ARa3+vSt80YQ22iyzJN2gfsEyREjT11q6Owj5Ly7ySUySxioazo/kvCm5A9Gbtn
Xuso2RngfeAhTvg9X8UMq1AGQtGo7KQrIG7IapQJqq7e0qCFCWAqMGxtJOZtBKKzcMHfZouI7b+B
0umGQpzrdOWLTnjpe/8wR7nrqTDDdni5Fav2G/yX5jEfZnKhOGgPJUq/36LYloIFqXajQRv+So7o
7R75pA+S/6IVlOs4V0d2Mp34Vt4gvGkqN6IF1aslmLt20aWAuytbnh9KNs4z4eOW4edBLexXOJHL
7i9a35b3zk/j9sFW/9egB5A2bouFk10TTcZk1H9RTnkgbEd2ISjGY56F4oxBZ+zxtSfPU9BiVZmw
ETiCW1zu6K4SGEI36E/wRdIQnSCo6/GOc+XJRlxHUrrdRdjrWe6tTiVKIzpUUFw7ycg0ulKLkkxc
v9hYxSvwNyucs1H/vuu1piGLtctl5VYPEYqimCsDKp5qtVa+pXgHUJF0/xK+hGOfMq7LMEkOwqQj
+x0u1w3Dk32J+6CCUfwZ/j64J6cPxGDv0wohrHieDZf4IWlNs3wIgGu836D6fpiS5nbwyW4WJWTZ
/OIki2blAj0ML+y08T4KerIzKgF1WjYzJUjJK7ZDKGLYhwXPnh5uZDewI5Y3WfIkmqRPw5CcxHO/
TpXsqyEsZ0IMg3Pws9z0f2f4XuZvlt8UA39J/puUn/ov3nVdHiC9MKhZm7/wXVNm0R41ZJ9UMRhv
0r9z0sqI/tF0bqFO2H9s/dUo5oek1GOxcoCmoiiVssQU2MQFN9yfNCljEfFOaI7gbbdvzMQSBciU
MM8OYcc++xKnfYNhnXzLF8jN+VOBLKUllPofbuF18NR0QUSTKUY8iopQGAJlPlnTjvz3lUB/kPAY
K9PrnIMhEVKQfwEqqLuawOxKqFkkmp/fhodoTHr8C/d1jLIRKB9r/9+Tq+l8ganMz4FPqBPD9bOC
e3GbsyYCGgYzlD+3Nmt6WnkkiXK/lC0QNtVEvfVZNR0xUEsYrdiUzkZEU29jMjS0VYinkQVvywQd
GrBF1pm+2ru25Zm1OUKUV8q1FtamImYCORVzavRJQvVP9jEK/d1EDzkcgubb9hPqyX4gAN53KY5w
e7SFEyEQ2d7lsAf1/bwyxeaTFmp/ijeMgdr/xaX3Rz15h7e4BJ2IuNC0bP0yjzIAvy+2HkZNlggB
np4yhSLofecosELKC2tVB8B29nnaya5SWIqGtJTCVBNYgzcg195yv8WMGUw1uGig+ZQZjGPoqH74
cOKxo1P1jeqSEtTPDWd3wXUYWr+FYHyImdzb7bLTBuNcOko5+4P6wPWn7Q2GpveRxzk5AHdivxjh
JCDJ/o4PlcHSkKyxaABG1EnUrhR9Q9CDgrSl0h653OX9IK8zHIvEpoh3Q4wR1+P4q8NQCiZrBCcg
n5bL0PbRHuGqnDH0RFhNKSblbEORrodTnv2Iomw6gukZoMTjwGnun3XGQG8drh8uKNAwaMZLlQzP
LiP0vrKVgcpKH0HBrHOTo7Rydzu0tmaaw6z8wD5odez4mj8VuRFra5bCR84AlF/HPmv5HCI0YyAi
TMCL/IBJOUv9xKfnIGLKuHGcENUBK/+V6gjW9QLCcKrQfaHcFMoSUbHnEoRU10mentS6cWPcu90f
NVaaFNPoigccz+SX85g5lKaljHcTsuRL5/KiwPEwXnf6Xasml9kG7mMJ1pX3aBnzXX2bYSZQd43I
yaLEDU/TlzpkSZTTVpthtPHYwW7U5kUsst8E6X7a9KTgjGTdYlfmHaq+5w9U0KEPlnUh75NhiKJ+
FiiFICgzFD1CZglSh0BbCR87/jgq7EPBYFZWCk6TN1mLiVbx4eL2U5QDSgKwIo7hLOQD3UQW/VLy
J9+joCxr2QA7kK1uuTQ9OXGgrhzGMle7UtF5gG3TdeU/VaZiQnrnO1U5ygkm2yHYCf6ACVlbNWPB
h959+ItOZXYAn8MtkDmvMvzYi4RRaB/3SDSlN7smD/pIEBa3sSl8L/qw45Pdm7UB0i4hQb7quPV/
l1k0DUF3Z2Tuv81JzzsWExVHvZkz0qDz4hLdm8hBtXiy9G7caYHG5Y3/Mic8q6NNvLj2AIkkrSJ2
S70/IPSsaCx/TpNmxpW+NHQoPtAmep9vjQ8UTATcD3WI3xjBq2+E+TPXxj90xKIo7Mv7iO4ynm+N
4le/ZlIFKVsl6rgbCMeXEAIQQW1onzwzACbBXpYQ4fzLKx6tUxN/L0BFFn4tNdddQJlGL7q3LnGR
kLjUEvL4UaqmshgTajlY91e/P8uQjnA+0sy1+MxMeKCKXP8FaBouNtBl2nJ1peANecp8SXjSOGMj
W4hSCkLi6YndJTKPihKNRyfSxh+lWfyvNPiEGzaGdFxPyp8S41TLGWdHdlXZRpx512fIrqb3p8Sf
HYgo2bItiFNPdr0H/nui9QYGliFduwy6mHXUNd1fPMVDKkzf8oCcefj39Ivyu+qZJcGF1nG4m/U+
2TP7M4sLmZ4o/2nRqEthbA/5dOVyv4cgMkIuKhLpKsgJP5bXqjeg/WX85ZiWWvRM2KwJsdWy4vv/
f9lo4UHsPELHj/ab/Pth81eyVSfD2P1qqJOu0pGYJJmuTAupU+cQH4TxXKoQ6+hlkaNHlL9okCn3
v82/BEozocOYEOXFiQzGQLQY7sxJhGV1QrrRPXtHC5FquxTTruAn4xlzEAhaa1dcpMv7blRqxRTp
6Ya25lR+mHUQk2KP5tl8NtocDihtjC5uCXupYP9Rf6vSZF7DqSnF2ODPMC1IY5Zd6RYK0m5PxmGQ
v08Z09HbsLP4wBA+F2MnQ5HWlMMo+2rh2ybt7qDcGeDj5Y2oNdMYjjvuY+4oy8l7/l+OR37Qvf3f
9TpdAHv9Tq5/fuh1PN7JePHuHMkxQdjf1/uWneMKNtM5IV18axLV6JzXwfFL+NjxShGxDU+hOOYb
RTk4LnIZn2cFbX0dZdE31lr71ZAXHYz3gGYOvca2Bt7ov3g1CaeiS44AAWsT86yVS6KT63imcvTT
z29M/nnatUh4oYccu3jB5rBYxA+pDF+G6bFUvewnDsvYdnt5xwqL8hki9KRHY7iE9kx+aKgBBFdZ
BbcieQutH4JbdYeggATjsohHYl/Eex1fzOrxwy1r0+IWiV4gPBKEYtAiWwZKu6mvBLq0VV6WOozC
yDjT3EO7tMMd1hJx/HJkP5nXE76Ih0eSacRA9wm0mm7y2GLDB300rquhb3i7BLCkKkGKdeOHnRbH
x5CBH5S8QO9o+ljqeoujZpbSkJPrIdULQNsBB34LhTpU/enphALaSRLBhFJd6kSJE2c7k7MhDzxs
wQ+odeDgqM0P2MaUBsuEuxOkpCGhHcE9I+tDYa3Uuv7XMt6KR2Zqj7QMVOj+CGW23wc5vf9e6RS3
ed8dA2ReJ5aNQS0KcvqPMeSp7TxN+Mk8FiBBVVXk4snB56+aNKR++lTLIghpq1+i6T4GwxGAzXuD
LPLTG8EMCLov3leMWVYrsW1FEg4ndK2vf9CE1pur/sGRIm40ZYenv71QYXfIsWIK6wdC3rTgBFP9
NIVpN8VdN/AT5RHpXg6ECd0a6usFf0uO2tUWGXDr3VC3EpnMK4xutz5vADVnCwYZ2elWs/725c9A
G7grdAMlfYOBIwM6ZR4YTs2+ak4DoMOrr36yu1c7/QB4XpW5m9OJP4UKf2yX0FcROxbG3/TD89MN
+rYKvRuePjktMGNis71IycOoZLI2VMdBStFQ3iSQj8I+qspzBk4i1IYbNh2u86rXBewaPaZwxr0o
0IufQMaiO8Jjs0Q1oFLMVLfBroIol4HWN0s0LbApJu10IHesFEnGlnUxCNDUNZAZkSyQm9680q6v
TsqEQb/oPeLOM7lPw0ZwqXvRRjWydH6dwwE90lI58ejC7o7Xwiijmh/Mk1jNBPj0wtJs2Fa74+yI
q7wBCddR/pys2lvrzHX3qBsd0H9rRm3x02TCcuSxagUskTccgjSlIAbKrAKQ8zOjNdy/Rh5FLVbT
190FI0wDl7yDbHc+3V+KQPkN3FDgfN/UCzqWMjYXk8pivFurVfzm5HhQenFxkrHBGUi0MMAoBmod
roceUHjmWD+fEyTP/Vqnp4hn/DJ3ODxv8Uzw/2zb1jb8XrE7mnp7qhUBD/YcIMMcL3xh6+z2j+OA
5j7isIGqqB7RuunxCfxcDjOieXvIr6Eg6gk37iqbnNKrgLWldaKZ6WmYuztUJT5uP6QPfxMob+tH
zunJfE/67OexIiNQfeqGlOx42t/zMXXrJxAqtHjaSi8IQRC5Pjn2T5JsK3sul499jjG2J6MEqPdG
7tK9EVJJELgBtXCX9SG3lozJTTjhhSpUnGcgVCQ3gsi1Jy2+EjSeAkN9o8Rgr8isqIY05BWeETYr
st6XaM7XZfAA38llWMxk1pwCtouO02X3e7w6NV4BweQVLxSzRJJfWupdnAERtqoisuCcQE+eWQKi
tAUXJ36D1DHy9wMQMuy99a97z2NI8t+jiTrCsdqRT8b5l5I3CM1stTd10+zM4SxVhZ8qYGk3fEQk
ciuNou44JFFQbqNaMfcaom/MoeBzDoXXEX+JZQBSDM3ePeTW0CMD2nkNDOLWAi7WrEfsOqLafviM
d7ciZ+x7E/jpoo7TRkscngr38UiNo77n63mon0Z+MLAL1dv9JyasuFbz5xTyB8BffDHHW+dqZc2a
ONwMqj5aiH8DZFrqbuNCVrBPJyo8pW6X1MNtEfzLBumg87Ma4WPmaKEeazHDaT6DNYXNhA/J6UBu
0wFZWSA8RF33kltOGt4SgR5qM08wa3wF7svA2WDRZAEfrxI0wIEBVJGYcWv+/z+QK3/63ehR/XZR
x0mgm56onQEOjQvw8bm8aO62qJbQzZgiTp9D4HcT7vMnK2bev+1H51rVGuMy59veOkatee9+uDz+
SiaQ/yc9p4EJbdaiUfRbvlI3vZnXvcu/dYPdugfVa4TcbNxW1VLt5FTz5esTLgeYwMp9GQqh1MnY
/IGkMk3v929uSGhHl4A9X0CBZkC1naFfThpvjHDb/wKtiQuAelSc4qsO+9g7n1TWEYrjLA/Di5wv
ULTwnWKtR1+iPAy66EOMzyHSOjUEKIrTnFnEcN76bigRdkYeettoMlPnlBrM6AXUUDAibz74u3lF
EWDMrmFDejX/GZ77Zr7arp1W2B5ixdowd5GT8s1Guux2JVURtw17GwfIccTAoGAZbRxMhm5A8AJW
OwiE28dNKqryzHdYefzeGN+uuzCZ0mZ/jgobzrmOtOYQTUtDQPNjr86CclMPpUbUOnxzwcl4Kj4I
1EvcX+6NFIVzOHE72LT6YgSY1bFXBpbo02dbNOizm3ZufNL9Rj9hnrulx2fW7NqhJL3CSNjuaQ2v
SRjUggUSCaiqvfeadiw82z7AQ3OGjakiRH3b3xa4FrtdIl4jZTJFa/LTqsYNfPT13QoDIONPrRL3
qToUA3h2yB80gPxn8jA9dSNIuFjRinsX0Q1KOBUkj2hHNLZ7ET7Yw6U50Wx1waxrsb6APn5egyP0
IaEovYi3Va7JK3w9eY5IMkqf4dw8R9PUHvGOG9avXdsKyXrpgkHS1KbNGzsNpu2L6dTq15FNID9U
ye2z4nVlMe3LqJ5P2X2Qs1XQo5caCJ4qpkgmW6ZI2hRQgPFmMYHSzNkykTjGC20lM626O67s4/ZK
aB7z7FcecLCPsFEPTFzZ/SfwjUCzfbR1Vf7SNn7zvt5JWLWsFTnDPFIbSSoYq5jPvorF2bUGQ3gZ
fwpvhMwxQ8He66q7ioB8eMggYl62qQWxD+x8EmXTXTOT9u+GPYNMsCQBverTr9wjK679mxBhrN+z
vLyFN4+OgjNA0leXTAfXEt6JbZfxuKl+hQ4YRxkENPSNHGqQ0sYpXZH/3JMhof+/xwHEgoBpot8v
tYC3MD2ITGy3w9R4rvFYFr3n8UVkvviy0qFUgi2JsfhH8YI7/Q4yzShSYshhZOMD6Ezx5OltncGf
n8+6+Fp246Gnlt1Uqvf0z1WiJm4fAh0X4m4cwec7Y/AzwrbwUcN63QNXjFkIYXaAYurbzJQc9Rhd
Qf0mymD8/LCRitxWczGfCBHVzgHqEtYTmoIRzFabIVmt0ecOe+B1pzzW4MVNohy2AEpwKcePbbbA
5ofIQOEu3qdMKWl2ttOc942B8rL3EqH2ycOtalByPOH/gEMEK5qXBNcfCLxPHM6q3X090JvnU0rc
GxRzwaR2qWf6VzowfdQbz1xIgN/e6YLHR8xZdtHoAH2IAm56dTgHwN4N65kUMCWfPoDxDg7r9MHx
KsUlUCXnwdOflykL2ncKjVkNZUqFQCuKSlrtkt5rXZpZYSNOcjWktxXHJD2JapxR5tNPWLrFdpTL
lfKVqsKqTBYwVVi0oYsl6DsANtbpxd7lYdTuN4tz7M2aIW2YbRmkaMu4iB7/8Uen6TKQvApZ3rAW
kk3Q5JeqtIUIsQsJW6D8JRmAkJoJPkqmjBoSEYMYzxHxR3Dg9KGKJLpLPcW0vqXJkEWpjsD/YH92
QVvhIN3oc6AtCtqvPeOl9Be7+ojR78yWahObJZF2IMirDWc0YBDNDPE0uzk8yKnqEiqcqDPzXnAN
QgDx7/AbG4qOTrIp2/4bsUQRFZ6E7cG7PjDSmxjbll3vFeeaxljXqeojjptXFS63Pkjdd9r9WNVR
iqL0EcY8dxOSDb6X2NwcH3R5Vrsz8zE6CzY3UVGw3iDTrfxVjiRHy832n4nuVlQ9yQEvK4foHLhk
yXtI7icWXSsrGltZb7lzycgYipf0BYwF0qYW+6dqAM0T0qZEUJplMI+VR9N+TDGMxTShQ+SwAAzi
BbkQmLS1iLRHOOhz5waXN6LjAw9bouPncOiIPy8elubRWYb4amFvvWnsgGBsEiLWLkw19enKxD3w
xzN8MjrRlFVXN4k9r5wj+PxDZmPjY6R7jjsjR+VROwS3X6zU80tIf/PNJ9+5AtVetvgxZ8GpiByn
s1Y3XXk1/XLVeyxUI0LbAEm0G0jkbXT7I2dj/Vpn18JePf1N3WypOG7BdewyJFeB8DxrDSbFo0Zo
aEsthXNbPoIQIUT/J4I/Vvxf3iSosI/rMJjySnZcQ5zMxageLjibqLaOBE5n9t5HLaHdn0Iz67vf
Lb4d4EXrkAHuXLpUx5SG/bvcJJDbois4n2VadYqgGIS4h8a4jqGnUsninjVNrzx3FQjRqEsiSOOr
YgvaInXKNDE9kjZcJZMaIV6EeVeDoT9k2jxFRwkXGHCDZ2hsxQbbpVD40iJ6lpdDOiT4Hpg6udQk
IvMDLUqsEfUEsBtW/Y5s2a8B1CLTbusqXMNOkwbrU6De7aSbMs0CYf+BoNRr2LrtjD1oG60Q3Nmz
RBT5hnSzaS3251xyMprGVYnPMgeHqJDBrHt34Ah5HXncyo+ReKXL6c/M/s5KODeA9p0xcn2FPHK+
qx6edTlFjIfKjDO2spunE07I4tqiG+dlZZvHvb+OATbge6HsDd6frpR4SuakFiWMlwhQtE2PioZZ
gl27oM4mqOPkqVjn4tOoG3gIUVaq8NxqTUFcq98N+o+sjJWsXvTe4G8eWpRbtgV9EIRzcxX3wDmy
ITPG1xpGQbUjJvjAk0w/W78dWxGQdX8ECUX3rDQGqZWd4WgZzAZsJv8dPqALtEoKq2+fK8BoNphJ
CkKMjqNwM44GuK+w214ZAiUJnueA82XMArouDTZypWFtUZlXxy48mvXOKo9rN6eOZJ3CzcgwsVF2
FbVq2N4jKxzBdmiG9R4Jm6CsLm+52RFPhIxUxsh5jaUQiwh+3bX7SIfZy4I5SsSToumVLNBBlY2l
h+3sgwEFQY/fIXxw2NqECMTnM/qIseBRiJaxKolSdHnl7w9CkyzhY0wChGJBthwSQ/3NkI0FJjBz
HfqTpjjXk3fbQ3WEPooqOshcXvTrVi0S0TjZzkW/XmHXv0jXOTCj9hSNrKtxotRXIaEXFnc26426
9jyDa8X8ISuxRF/k34WAs2GmSDb3/oN84HUIsWkWS9v5WDkQyGBt6cI3N+ZSmtWd930+MjKZ+R0B
0NSj9Z24zER76iwsyYykP534SwDdX5Lw+kf605M2ycSUgfOkNoH2LcnQuM7WphxzCG8rihgUj/k4
3tcmYI+pe2jUfN3W6cQt9/ItukxOxVhtnMR8ouCxuF76ujk/+mLB2r51vL4NnAOPDbRVV98rJQae
/ryUc1yJLKiKknajbR7j9BHYCcaaJXJzW+L7kxPOZhGmmKWAM6LaCAQd/6Cl59JMbkhgGww7fwpu
wTZ3kU+y04IseJhHriZRZTwPksJ++ZLAuy0IrB84ZWeDuGXmBCLiZZlsaoVYsSM1k+OoTQXIWo3V
PrMAcM9PH3hWDm0JjBOgVhqAceACTwc70EQWcCEtKqCFzFKPTbG3WnM+0c1CzDTgtoUXBYW/7LVG
zo7AD4SLScEbYFkpMeEvyvyZxhgiNY7bqmXU9etBc81DjAVOZ6vYNfxMiR0uThEnYDi1tJQweIf3
ZL0NanviDU3Y9X1BwjpfQ2M8zhIt1r4ksg0DPajerSnIY4hBLt5hYLXzBfjssXlUuM8GDHqvwaaa
vOJH/O7p9Q96XpURi+gI6V4CEvICANGMi+RPj8JYFxvV1UqYkDK62ROcN0WM5zfnfV1dsZd43eng
Y3d0qvK2CT2dBz9Fg2ljBAMCg3AxNCdSeYkfddMg5YM4CoKXDO6Z42oCjUF6+VXhXauhCz4Lfr7E
cX5v5Kzs4lOiPZozjTQ/DgoKNKL0QOqeqs2OnM6eij2ivx+9jdF4CBLNOyro/6dcqgCedLx60GKK
82lnvj7ICga2KX8pbyOMQUHpoDVTiq33TZtwpVDUAJaikJ0CnKQdOSTAa5AkFH0JdTAp3FF8D+QR
b8XGe0ZjJMTfPgRHMLw8kvTTmMEA0Y52j+Md21SCP2vHzXoU6YS2Z7aATYr905Yu65cz0jvmFHUx
FWi7gyRrts4/LPMIrsyM1Y5d6HgCrPrpBU7nCGS8DIuAIHuV0+FUxk/D9tpdvREWLRdn4sb6aGKW
27axxl8uS/cpEuF8mN1JbYlC6Sc7tqZKH91FZc+NTEK01YC4xfvFeIA01wrGhnzOSO3Te64LvA+S
jGXoLkq/1Kwp7QZgnkCExsKgJo5q9HmeyLfvQ+FC6Kzbe9FEgI3p0CzxDEajDDjjrEaUnz3FmkX1
ILh3TWL6DXqvkbJZw4Zl1AKQ7CmrR3x6g/QYbxWhwzRodW075YzxmuCd4CpH/hha/HezOHySCL6b
wPSDiJOd17yH8TYSktLLrOsLJMd8vO7lKLxdBfvm3L/B1ZwPiFI4hkVUz5bgDx+N/EEaZtmdXmQC
8vQcYZT1AZl++4nPObd1Ah0P/UYb5XmLGe+Hi2yIJve4WE5o71svtQ/EylXXOLP4nr9QT9hfgxGI
/+/6twN5rPunTx9LL5dFgSNagFZ3ytAJaHdx+naSzH8VbeHmvUHTfOCKkLUetV/XvMqEBt0c7X3C
RJ8mp19DWDB7EfjuQjTOpbWk64vNC4tReutKDYWzwi9sLmh6eRSets7/xMGUMLhqsFCul+n3UB4B
WyTvDiWRuWUUc87Wyqs2sQkg1suFmj7v2pnZpsncQDaZWGNee7MOmyFTPsg/2u8epWzH8P7o8+FC
F95VDiXWKGqBD8ZHLqWFUwEU5m9f0zZXQ+k8CL7fRUI4eRCdC3zxnvHmJIHH1TY1Vg5WMfqSbmhb
gWJiKiggaIONCM3cfZzcN+Ozjml5Ged8SDPxO33sRayYP3ClUnoJ+8ebRhKZFfQ/az2bq0mOXTkp
dZbnGEE3MfRLvrGW+aI7WBkIGu2qYLVG9Trxx/KbE6YRnTN21C9tMFulF6MVyZEfifjlgWRjxR+l
jP5he4U+EwgJt/M67oVMFpIMXldtBVP704GRe1t9MYGRHhmoiiCpDteNsuW1ggpx9t4mpyMXXzE1
SxGe8id7Eb1lmvzRLxjHwbr50cZDxpseXkxz/ai736HpFiIqtxsRcDAhZxV6y8hiXdvCWI+Td4Tp
bzNR6HuhTC2IwS8bwEtW+eAPmZnqqvWORr+7Cb7m4hwAxEFGpKbeUhlxW9h2+qrYuZSHpBSFzR7h
IE/sT6mhrhKDjf8iV8fqk/k4eRVuaSjIkugLJLzrn+hcD9i3Udu4yjIEzzFx/CrG0PQrH6IaqLg3
1j5DmcZzIWOc9D6WV42lp1Zk9wXREOHYEYnVVfNVcxM8vJ2TpuwNBdHZJdCh2xXSBQsn9X7bNkWz
590xxIkAx7Gb4sXbbxGbRjjXXnIjJ6czk4KQvDyH3i7uK88NdgrImJaKYT/qIgEQAil2gZly+WJi
xrW/niorn0Yu6FlyVuu+DXUUyzRgAB8/kFIhBZXLyGPS0m3XQUdxwMQRxbOi23L+JL9Hdkqar8Hf
jdfi2j5BkKl6vRQAs+LhFfhaD1h71x9Vs1pNFHDhg5PT9+qRQ7nnFQ4s2NoMCL0Fn6wFH8Cy4pfj
TqDh/kAI+MjvM+5ALen3PhM73ZSgB8mgFvKHdDR7LPnTijwSqvDphSZJJvVNdj8cqICXn5JBejZJ
EaRD1ZIVAWNg5fb6a32x2HZJkyt0jq+o/YeMukUG99CRnzJkXXqF1r+9bVnCcAUT4fm7HVMbVZ+w
YvQx0cpbivzWCU5NCESZWHAUOZ9XHJLgebWeZxQZ6Xp/i3N8IqvMeTHim2x4vYZ0Zb1wuZdJrMvd
qQWybmFu/jk99Be2GB0+ZeMEvi560Tv/Cjtx6ZiYdQMD9eNppO30J/fanwDgZqZf6z4FgRlEL3CC
uVxiJc+N4ka/8RM8FotiMMOk3cKjpqJI0I6QOXOF/ZvAGpeHLtz6mYw8gMLnuMLis3z9vnuK6Wdm
EwEqJH5j9ZFthKYZ3MXZebppVuiFnDOWjR56SAr6DOpOuTjwum+45VKGmHT7CJIC6ga8QUBzYORG
UrN0SyOaAjMK4MKwS1zNcaMsTLMB9ySd3wC+6PzgAz4+GxrrBj2JcCNJ2Irtmz1UOSo6YVRzbxUI
yfC79degvtQx1HIcX9gXFE7Q1NDe5j1gg5NBAc4fzy0lyKTkRMN/mJOFz446DMJr1TOsN3l8EPKO
pRHd1SLhwmfyakzudq72opPV3KUTTjhZZq+FmCGDxPPFGLuG04gERkyXJXab5ayZqcaAyG5Jhwni
eC6pbg55kVXwnUWlmR2aPXGLYDz7jF8i6hd2o70gt0z0nSJExPu5pSExyTspNZGEagDLE6VCsFGF
CRIfbACNIS2nG468qtKw4UGdDs/PSg9uIGVJTx2TQz3YTB/3ym/iMDhZyng2dHlPuzwxv5SsI74V
RmvIxQcAJAyipDtOdZhbftyAK/JCjgptdJshn41umW3GRI3FngqNNCqiX+wX+XVF8N23+9AB16uH
cXX1n0YMgPb/LS8hofnxSQZ6gWrpKNkG2FrFMg2jT4apIO2M0UFkVagJSJxnkyhGjNEk3Grs4l7/
f154gD1V5O/sbbNtHfDBYuoGHWfG8YwP4pcDawRzYv55r93OrZ9Pn4MyTS80PRLXcI1kys+gQ3xH
/Cp04OT4jclyasaVSOUDvrQ6cLv6HySxHRQ4qqe6R8rTPyWU6F6SdVoqIwSDu3IOp7sPshabQXGl
BjwLEzWL+/4KkPjQFSC8eOzWrs8/oDDtZcwAZKZliclmqg+VI0OBCNMfvmdUNU3DsxoYST5hCe1N
kmIe8lL73+YZOjoo+4+AAQiXnSVVI7HOzTRV/YBrRmy/iVHj25N4QEpVPrly8nFPtCFpszRC87Nv
Kxv/3x8gS3swzXt1XYdwgxI/kivBxW4dX9yBUKZ3ye5eO4PivOCJZ8PT+WsdgBWOu7qjo3RA0aSn
Othu4Y1+3tZrAbI/HydKJsK3QiSikWjzVLhpBoMWsLFiFuQjOt5UmbH/zrX43DGAml0VA1tXFEhP
Y9qtt0YfaD1xtdS0AZlwQAw3snOecKf4yaiwuDEHd/ERTdDSuDIU14ey0u1ev7+/vjBp/q+m+13I
tRUQ70jIS26u+fxrLmjpewnFpj26mcK/s2THmaGOYOd6ZBOg7h3+czcWez3FuGXrlNRu4ka97Ppw
fTci1ldjA9LJc4VS6D9Ksh1Kzw7lZ1yYcN/FPdaCwJIg+ts6GK/HFkq9YJi7hjKdwTnSVmlLooa9
3yFB70Y47v1U1Bpjpk1Z0PltC2ehe0qnEaxAXbEsN9wHOtbIwfT3xqk9Iixw1mg+caj7NeKn0YlY
lq0GNMsqywXIAMsfBvLB/4ksErY4QSDc2sJ3Q7KnWvj6fNohOzq6eXNdJqCJ3oEpJUZCBXBY7wPp
IXTqsTus5bx0OUA/XPXw/Ym3a6FEWPTfzfyPLf9ZTROpFc4xfe65n37VhW7KFOWIoOFNKXhzhaER
J3eFz009Um4OR5ugxQVk+dls/VoF+dtJ3GrIUnkR/5anJcxNU/28DrjXv7JpQvLxcvH7RxOIzPzc
6cR/PExkSHu+7KcP6Bx/E4nxsUdA/4Y1N5GJk3jrGEwIftR8OwYoDnxCliIfvib7DvbmiQmByai8
TwA4xEYVxiMdGh+ZusLHeVoIE+8+0c24rIrxomFaHP+IpjSX/1x1RN5Tw2vQpIDKUXVNrZGW5/OF
sEimz28ePz66DPKN7LMRjhIZQVI0zRsqhlb/LDCL0hpS4hE/uV8QQQxHI4RIlQPnH1I16KjqF4u1
ymCetSNZiNtOBhIecoYVSTk2kgOrn7ck1jPPndpb7GvWE2jwA6I2GjaNIBCQZ3inil4WZKYvuQG0
BSK7fTcAeKFzQVw7/aW5mcAvv1clZsgjiDCtdh/hYdAGdZyTvMx+GF20KFQwOOchI8agD3wnDWi0
Xo5ynBgcX5l50aubIyZMd3zVhrCdSWzTzIyG1TIC9KuDISw3I/0XHO+jlOPyy8QZTDAkIfP2JEH/
Wf/RoKEh0K3QatnWUHzk5fMSmr2BsU90IerObH8wVbeoQkGYZh5XtBndCCGGeBS5DcjHqmPUOr7l
bA7/aAHQrwlSuJqRhSDpvTgafzwGR3vpVzWV3FJ881G+Wq+wuxubQaq17pTcaRMshSfiGG/1u828
gEyhloWnr5Y2Y3LE8ISZpRVCXP7/Z2btGaTyrxJI8lj0BcH7Gz9LUJ79LhBsvX2WXkDWWvcAdAFi
7XQxOez91WPgrHObHQSv2OdiYeDNnxPo6J4Nqr1E6RstgLoqe8cujuKhQWMCFUM9IczKngB+rj3h
X/fwyBFZk21nSpuWYRFGT1d8uUgK+HVxJl6nCtUljTOhTiemdq2tARzTsB00bafmG+7LyDvkLwxC
P7x3qOuFk/SUrl5MRAvopBXiWT+IebOgO6tu2NNUjUnHvZQU3p3a/7gi0g2s3gZIohXEVzUCCx/o
aVSlTNcZduEUHznC9WJ0hwv0LIntr9hNnDAg5c6TQFwpVhkpi6Yqx008HyFP5lni2XqwJxiEdN78
IMR8TxQffQXWl761IkOTu+/fu7M/tiPQSEfOGPNnCxEJovcg9gxR1R07VK1Aw5ndU/0RMNl/q6d3
ixLGSe8kU+akfsYP+/mAFiL7r/+QL4v54f1TCzE96p1ewUbGiQNGjVp4leAZ32VRos8QnT3bs8Ns
s9VYy3IyUXjW+LdIM9oNW/dkri1pYsBho6DL+bfP3Nr1vmN5VkS7HmtVw/yEIlmgxumSISQOnxlY
Yynt5bmtNaW4Ypf5UYHDbabbuw2fwjEvBuSW5FPQjULGEKDaEnqd9se15xuU7p8HGPCwnDQwa5pL
A+aVB+gr9ukJtf9K0eA0W2/EnVwgKRcMXEpAOMRfXJbBpd/R5LcB60MHDlkvVoFrqULS0hpEWxuc
Ka7cM2bfi2YLAtsim2Eo1MmvymmFDj8AMvc+FVot5p+05tv0W2szXeDJGJQGRM7zg2QY218kpjlG
eP/usYBCHKcoWLWUjh8oL7ebt0fx8Xj02d47v52EAyLfTBEt/R9CShnioQOz4drh8CQzIp8ZP2rz
8DY40RBlXq80g3zbGGNFiC1+A3ETzCVgmD1lZllVDfxDWK01Lja37dK/gSGRa/zdEIEBAVz1vQx0
O3Fhphdp3kCd76UnacfwwqeEstZ9wXloWkbWLw/HHpaBbrYEyBzRTzjBjlrW76jvOFuibFo4Iqi2
aOSgSE6lbKEycXpdmKQrI/Ncj0+TtTnzRXbpOvmFv3lF/5r3eawIWE5+7x8Wjjiuk5VO58Gumk8B
mn0gIOvlfVBVZt1lYkxDrzJyjN/kKDR7Rf1R0rrpqpmMrr4PUrIGvPNPZV8cCqiO8C3dliD7DiOK
nxyPqfjsVBa2cIceF/rriR2V2it3OMEz2B0IcFECS4/tAAS0v6QekB317TGg2qI3PmVtMPqvP3di
AGfntgY9KlQYNM7s8KhnRXmEZgeHbeaP1uwwk27MUW+PussITe6U2oE0UdbsNGaeZI77LhnMCH7Y
Wn6zMXDbaKdK0XOyyjtfoX3HIKPtahEGxArR0JX9lXV1Cbz8ybHkFwBoYRJBQP0o0LjVUWueUqck
FOEISB3Qm3TIncR2V58cMHBwK7AQzvRMWcpXV5jiwyt+vyPwkcj/6N/jdhv9fLf8f2VweWlcYuqI
PwpRkgpyS6NUSBrVeEeouhRCbAf0qHUuU39uOU67SjRSU0CuvXpg5YX2mZbDLW0nN9YHSvKF5ySN
pLYdoRe9De/UZLGKClZOSz+VQupymD7QHfFB1JdpQ6fyurhodJ+FTOFKI19NFP9nHoPLv1qYghaT
fI7M7j63Fbvqck6uRO5Nf0lZinC+TLDyJ/En444v0sC7HCIkpNy6thrfZMjszY4BtGDQZq5L1CRZ
dPYgVSHLQbqFueZyDrKP77JIfH86/bUJXulJ8OVdEGETbRZOwPo8kXRQzoX7ba4TjaF646XSYzJa
+CcNxcUwe+7e5gTiHfkoAVaMyEaBsKDDtfBENlLZI9zSeYRLMxHktPugd3c2TMqDv5UXH2JftKc8
6YmMz6GAuU4dpV0ZgYa4Dx7DiEmodaykKq6AWP/X951TeWxVZZi/vXt/PPw6aofs2MJu4fNwK66k
u3znN2cqPrpUcrlkPUUgl/bK0Q9RfgBs5t4nDd3dQKH0mSOnFLv6R5oQC9Gxm226cH3eZ2o59WSK
Eod4YHk0jlwtcEH7yU7UxLhQPdFwE3lMO1fExoDxiqKkBrjCmpERSBu8LqTHRv/Z1Ak31SoI08ZR
wGF0H2V4IeRxGZDb6doy3F44UWATir7VWr5CwM/d7s//NXllnRHlsayg6f5HKf6pyvHGLo9wftL4
uNRk+DCr380xOlVBBrWHvPGbHbqYQfNqEIEz073XQx3ggnZ8EBqzVcyWrDy3XY0/lQq8g5na4ibV
uEBI9lwGzhj3XPRlVy8Oaibppt0qdKtjbEkY+aAR8pl1SLu/4qIjEk9wPX9MbS78rZiOSEzAN+tY
l4X3eYE5lJiZJCJwHjlIRCrVVAGtL5wQyAsQu/sNOGakBlpUGTWm1t35y3oQb64bXqIxnHfrdRoB
at271MIhOi88LEtgzVEe3cL49XzHdZm4YLbm3XUGt3UASKNMt07h9JDb50BYxg5BuIpcdn6Wd7r/
Yj/YlFofTiXNraNJfjDdIZaypTsq1ufcWsH9YWAqH65Lx+8MeC6I5R2ugoB7NsC1EEC8wkDWd3fO
9Iy3jSbk5w1nLQ0Sds7meUl9OldWY+CuU9ikSnKQ0WPjmGhBl/vR4VaxOVB/qXe/y3ZS/Z4OVG6h
QoEbBZqRHzGoDXpi3WgK/UqmGk/scZemtmhDqBj/5GtSxFTUKSb9YMPiYS4BV8+iQ6kU0DtA8Vzd
B1NjKdc06PVFjNNq3ILQDG4smx1QuGywKxg4PZJo/Vc2K7HFIf3vQFXwAOiC5Kcyw4FOW+quzU/5
uxSb7w/rll4LdxdJ0f1OVojy3uV3iUZVZFarIucfSQEGSrykW+BpVegNL3pzAn77IM88acZBFsPP
R9Oiz2xipPi5DXqUTmJKkvO6Y5fsSZjD+ZLNdYUkP7xbjX1ctf5P3NlNKBEE72DxmO0A+PWrxfo/
rNXw6k7OtsaPqMynHQLyhu+8jJ2jr110PpXUTAvCFfo/um8BdlpM+uZZIYNmZaZziL+5J5IaebVk
0sDhfqT0Y4JtyC2VYbLYas/9pYKpMGTAx0ngj0rIYD1wunsSGWYGGBevBDJROc2eHYUA8PoccggW
wo66pedGTSZBMu4I4ylacXjs/Lz5IkR/wqRmbxIpjL3pamcK5zSGJsAFa5E6RGDH5ky+yuXw2yw7
QIPRPMWH4ZfEBBuJQmNxAqmG7raSK8LmFJCCqXMT74rq32VlRc2H7VRmLhG6PetujB7Ea0UvYKkb
VgRww0RsZPr9xVXwBG9CI/RpKp34TpgeByj5GpzCDHlKcPViFdxxrelEoxN8JM87pWd+i7mlFPXq
1LURAxgJdDnXOhGW5XLig3zIdLOq3luWUh4XbK0fAPSaAmwGzsPV+MzOezaVs3hGj7mHSDVpjFNq
9Oe/OfruoqqiZZjO1YKjqXuGbXWw1QJMHkhTzKAGGW/K1bw3+iEO68BHg+JlKXl0CCWb+FAl2gU/
axNceOdxmNs0INRttIGek0xuXs5WFZZlK3DLVrobSE14vxi9snFQThTvwsCq4s1H8VoCJBDfZC8t
T+llN436IrVh/4nelRwvv873/CJROIQUJo7n19MsNZRlHOB0A3UoFTDo5ADjBaQZoLIWnqibwRG9
4SWV9Vk0RHkjlT78gUJptJareX8l0cTE2lrXCSR2+n4f/6F5nwDkGdCNETbB3QSvnfwhKnFM8DC9
b7MbXS8G1SkIN2Xx1d4sQRDZu2Ai9mtMxV8MDjncBpf/y8f2rKUvW4SADoLiKLekcGG8d/8/Y7xR
oaKi7wDlx0YcLymCkWJOcFKAFc2o//Y8x3+C4g8gUIcMeMnfRZln+7ohY12spjrkoGmMr3HpjKNS
ojMW37PUajQt9LQDYCSht8EWq6udxumstY+1ENFSZ7YTyjQQaUZ5uxJqT+yJspLsc38U/InncHAD
OwjAz95eEMbV5yNmVpW7bQ08IgMix8fv7kTYrfMKoAY2Ou6ED8SIJqnVzMDXya2ZBskC7I9CYtqX
w3Kofew82Bprl41b6xzX/WIv2EJHS6vgWJFyhqXoSXTMALHu1c4ZnfKOn6oFeUi1oMNb0SBp30fM
M/kONiIbt63jcpkxJPbMDgvDNjmIHGhMcqHa94SweSTS5TiYyjueP+zGCHjNYkuYUa2s2kArcQrV
uhV7Xv8M00Zc7GE4LFwYv20axzsWsRysxA01uODQAvhwwfA/KC+ErOJw/rh6r7a6n2MrMiCiueHE
Ni7LNCiNEM3EudJiHAqqI11WKUhlCZZZLZheLlfhC3Kqr1M+VO/usmV6gHoBLnb3LyPXNc1lIbJW
6up3v1dAdY5b7kwVdmK9EvgsK9oK7YUhAJ7lO9sTTrkvcEWdm1WynEN6Sr01wQCTb0QL4uTYs0EK
GkgccMwDU8SIOP2T9P5gme7aJTuvsnofV52dBAFNnnWY8sVVTDlEdJzumITLxQz9Z/2Acm7RULem
LqcOj2zVanQKn/ooVOoSGdUt8AlRrCqooTvdOL7wGqSF7w/kSGXLCplpguT0zeOHkpgE5tXS5uAw
6shNDxUwag5PR9dHDDZnzz+nboGixER0EbF5oosfH9BLKHWlpjRNK4dFpZAraSJo3lWGBW0aoAl7
Jp1CuH6em05cx1KsiMuwu3L1soljH+Pc0jN2JKbRNpJk/rakE5quwcnWA4VJTYYPkCM2hwdg6sp2
NlEIJidiubJ1+EY8RR6cLGzC0s8Gp1pjdTNjjMRi/oCvrT1wLIcJ4KAKCeQnVF7y3Dzk1oRoWVxt
keJwrVcpP2GtiN97UAHSc0VEqcUTIzMfEeKGDYSAIUuRxYdnsJB/1tweUI1nZzT8EErKaoXVogMC
1G3bps5Fx6JUxB1ce+4/aNxPuUV+ly80jQgHZ9Y54CDqeVTmTqvMqxUb33dC8U587kBaickbFs4Y
436XoKuoo9k9QvrNS1CiElS8t3mpb8+Hfme8PNTE/q/ktUOMhwA8k4VSI7iEANuG24B/zUtL/k+r
J+xwUkQrRTtnPYXsZnGQJU+2opJKK+DgmGK0uzEqR6t40YjtrE41DArjhJDE6vRpIwykry8sSJE+
V/B9mEMo4A/RW+39Bdz+Oqsjq8JWbvaopsul3GsZDpsVwzYhfTvd9eioHBtTa7WXP7SzBlVszJZF
aGDb7BPhvp+2aaHmJ6P/owYJAq5AKJas6fdFeyZcOWVMk3p+NNjXE990qnLrYF0ISdO+HWJ/UKVl
E3Iy91yq3u66FDr+fxN9uK+5pq2Rz4Yi4OrHdtSPhWy2C7xJOT2oAkV8BITPPQsh8h6kTNfgH6S3
mleo1jXfh8Fqi313WMLWe3rzcZ+eNQJmlpxy3eL2NLNYkePVKOmLuT7qIJRv4hRz/6cqVsY+pEnS
5B+4Z4TfzBUTintGgK1hg9prNtfCjGCJWUKEL5Pa7XorptnAy+hy43qWSxk/8EQ2srAOxEBZtdIV
cOgP88GAjCrXLm+WDoJSNFCuuO5ss4XXy7PbcYUQN1aQky/cE2/WnTNtnJ3ueDIOIZNdD3csmpdm
OfsNYVADZq7ut2oWBJNfFnngjfHK415oTT7k9KfTPg/n4Ln3PwEBMRS3MnM7o8v9fHc5o+LIzj9o
Iv9Q9G5gWMAexlXJRIZfIWVudviHlS9i0uD0cSO2k1z9Fg2HpKcNTGM8z8jaMmUUisjdKn+50RWG
knuwyyuPtkiYA6hYOr/JTvzZVALOm0qSViJY2K0b75WaZkOqHJQvLtdPH/y0KoqIrCReCpv3uhVx
2oL0d6eXoOVVekUv5T5PSQC8pwBA83h4NKiz15pOpDA6f3cA23pT2tEPUhLl7HCXQLjmFrs0or6D
AT93/vM/kawKwIKfIaQViDNoq20WkQzs/Gy33l+y6/dhAtTmHDjOo29Zp7QlNl8nB3IDu2ihrw2U
p0kprz7o4Wafh8V6i+22CEaxuXxXmGEogHTZN6icm/Pkd77qk2qAnRL3NZr/9hsYaHjQulE0UQrv
KIBXi9zQ2wWr5BxtV1r3Ovz9Ngb4arUKghJuBnarhXj73kpdnaJzpf29Wxbbd46caLf2ILzLL6TW
QevVolo9piQ/KLuBS3MQmqHZa7lLdI4jzGWxce4r9Xj6yjKgXIVyDtPuSeQxT+uUMnr7DAk2e8wQ
tQDKDI6Bme9Ir+YzP1PPM7GEa2gPGHktB90/bugqpmSn/g9isSQa1XEGlDAaJGDMgEBBzP5f4GvW
ZPd5vC62Yd5I6DkDXZ8kKtvzJ77pyE0cedgQUX6bOmpXC9J1TMHG44dKQo1qvkG37TFQijUkhkmn
O6lXPMR08xwdWTT1z4bXl3JGRVYr6EoZkpl13VFJrHFwIHqWzj0xxB+t6kZFVMYuY95FfjkVlFHY
ZwO0aSM3dX5vwhLDPZnb6mVYtNYmdT2tx7RGdrPrN2/AuVMj/+5PvzK16K5X5JgVxk8ocylNfFDe
3CZ/ZGct81LXAhONdEJuqpFqZ9z2I0Eg02IBWChYiY1sKw89h2m8tJe81UF2BO0aAYrzfabiPOi1
4oJtLRtHuw8xWstRny6eGFDFRKYE92qRpUoX46m36+SChKMnqnjDqvY3CeVNHICScrv2TrnPU2x2
5NGY6LJAHRf0fN9QhESgHLmT17lAHJiA91ngJQns1ULTO/YLlslz7ByOxbvWvYFqQwxVj1U8sodk
n9XdZAWo6/kOTNK3jiOXcS3HabSguPTs+4YP/xJoNZMPpJSRnVXyEV3ePNfslP+rwfl7nBUnlxrh
ZZc9SvOkRy2DZr2hMX2WIBzcJ4wWAJKpwU6qGrANscat2C5NbXWdlQqJ0cbU0qsZBKmi2eLwMjXr
W+lsjXY+6RaoPmrnUq/W3TCDyAtAkd1l0UPpyXe+642KizymgwRdu6C2I3+pqkOV+1nQQW6s4ViN
ExFbAD099U+4Cd6qmvpL2N5zHXANJjjoXF+3qarUH1hmyKEBm/h1KtSEpxiBaN2kRvTh6fd/RdWl
AlnbwJoP6QkOQsj54KjcJA09UTM4HxPs1qAhTKIXgKAuruO8gKRmx+CxMCJPglZwsYywdRQpg7DW
RMRjzuD0ndxyEzoww/wcP3uYRkRFJiDpJrCGrDZryoEiK95JfYppTsTW30BsOo4SVUpdHKNIKdlr
T3w7bG7iNf8yI9aKiNE3qH5NgqfemlmvSATSNLUv2/o3VBdsfe08mS8/U4gmRklBPULfz8yoRa6S
sOATqH5G23mtqOjZWOKCBywzNhM/+kbIyIb58LGnHy0ZAHTMyBh+HecckBC2VB7AHzjHeRfBXlgk
Lhxa2OscSpPjkQXlpCDKSLcpKBrzt7M5vs4jZsXxxQMrcvd+P3ITbsPH2nI9g9/Ud0lc7palgWMr
m3dgpS232JdIQKO09R6n96i9kro4N2iKlL6GU50tb5ZRrlnJ8zSwaDpRrvQ0+Ty/xRrskbh+XNO2
WV8mYOn3ZPBwFVfQZMnkLmZ2RHAHgjCsE8d4/YnJIhHE5hGETEtPoCNws/cXUPSqCQSZc97Jy6jU
umk5KeY/TOMie23TPT8nWNA/isSGVuQgUpEK5VsRqg1Nlgiw9VCBNq2vGoBG9mmU4qa1rP0HpyL0
CWG0cAl3+ld8ANl3WOFPN1CgCVXpiKiWSWvzPsQPqgD9BuXzZUeGrHRdb0BCYM4fUHc1xKFyml5F
z4zFh0kInvE5t7hw420qMLqC9+W0Vm868r8h3I6gzNdrd9aCdaDw9NKz2asKJxTivnH0XFm9Hecp
ZgPIKXymMuN6F4fiHLRNg8CalwUmPSdlHLmCsjtNosKpVMjgJm6fpZs7oBGTjM35nF/AFSV2H49F
5lZn7MyQOHpKzTZT/iuzZbafIqB3A9oaCYCM1Nx3hKdLMAxHHuRUzZ4fxNSNxXk1SUHTQ7aNn7x/
gAgvft5OGWe8/OLRabJ1VVLllV+XzE1ykGjA3ayOMqJ/BSiN4vIP4l9zEamVgqnWlLSG1gZN/K6j
pcoBgfQnqfXxdfrgowXG+oCf9+jLf4CMpdHanPpBkTGBl8Bkew2cn8NJ040jA6nrKS/ChapfKGla
lVo9MoKcR15aslZbIKCHtTSaqglQI67ymogqNNkUpVlnt8YzZwptJ6q9dSDHsYdsM+2x/e3KHOrk
CSa9XaTpQX6yRDbF2O37MCFeYvlO/w97SP6JFuLjflAebnUsmE4onMc+Kx2w5Fg9CzZ7UANDmzsw
mex79ZdCqcYF3Bn6QRJsEyOC3h7fYXAPrLfA4pBdpXzmyIHVBaabg4p67wxdNNVtm/iPDfnpDZOg
R2+yv69bWuhJWZAej24FQvwMmDL75SjXdhrtJ1r4X6k0+8VmZPFOGhbw/DuEbE06rIKmdleGSaPx
WYk/IHuzWnPCNRrpXL9NyZm46exwl+rGAlKOpm0yfZqIQPUcmTGWAFk1v0QLa0b9M32EV7iJXiIe
v0oMy4/G1KJyCyMPhFjhYJ7p6D1kxm8XJGt4F8r6Tk7C39n3dGoWTWtQTs+gxblpG4D/H2Q/3xbQ
vQyfALYL9Zvv/u9E9p7yZILJxsMPU6HB/uykF/84pux9dMtN0oGhFcdzRACiI3rmpVqlUryjTkOm
E4KdmCs1do3FnXvapEERDuAv/Qt0MLadqojLXLY0Bz7pooMOxG1M0rBlBqLs4/Hv6IeWiSJB/nMu
itWBGW/adLl3cyslt5nK0ff9RIh+DzveAW2TfFRufLxdVaS0nbIMp2fbcNR4v1pB3sqweh5So15v
yTp/VFG41fS+MjzaWobnMChSr1Q0QJzasNycusxH7gchU4CLNGY1cGzPbNis0LaubA98BRoQEBbk
jB2EsdWVYWi0FsTojPO1uaPfBbgkrmdM5Z7+6h5K9vYZZBomv6zedO7BznN7SIspNYdVrK3W+Gua
Sm4Sm8ctDzPl4sCUjzYD0MATeiEotucxqB1rf0xZt0Dfytf98vbepLIxUUTIfNOfgeN9COgqjytq
mmhow/WvmMWz9YCQNt5pERkanhog2nXiE9Xiz16VMeXTuKLGAMfvSJY6Mq7QQy5W36PXtdp1dXf2
7tGcfc1//vDLyiEBXnDSVIV3iWj0IBbXtHkDkPTeyRfMuFwhaZq0wVQrYEMiAKotqXT7V4dbXrgY
053RoMRJvtKMFmnu6c645sPI1oCQ0F71Jq8vaUl3Boy2ookntYPdDppI8OHHi/7+s+qVn+eOerO6
fBtwCZjGF+exZGIuMaDjdQW/PbL7/k9KYlF/7V2ks+kQDa+78PwgTScC+G1TnIxzkRijqqIlN/CL
YGy9CMiz3pEBYKyxLt7a67YDkabaiDAlado0/3zzPd6jeEQlu8Ok8pZTUWRWFq7RZqUOgoSbkfvP
I5wqvOcmOvo01d/Wq4B4wIsR+n9YBYU6zCXwOtjQtdleUWgHevoExhU44Vlk/Ae/u90QvYM4ij6G
mFB1yje8OSV+WnKYgkMKZJwrM6SVWviLZhlTN2eVsRGxpozNnnAsnxME8N+8z5FMAbRpgw6XIU9d
ndGoVWuLbAqvGAp+4eflYTzIwHtEpEkhhoYXUqJwBumsBA65jjKVY9PjDtcomNaMwr6xCe67U91v
Ttnjg+Y41ORaaWMalSeqBo65torgSCdgQv3PSSJQQm0vlQtUqeS6jyR/Ug2GIZjoD+vds/QamvQU
a8wkc9wuEq7QGXaBmwe8FNBcrBoa25uPlVXeiMAl4GcVDuGSqt9NQc0O+qlUbW7K+6jQGZK0QG4C
JTjbOP1Zv0itJRqHcBFcMAQbL8xE0HvLClVKhwOPqXio1o2j7UGJWn8YQd+/MEsXi1o81JOg3V27
DLP6NwMEsFaM1QvEoGAvts1HKTuRahRQPpf4DMV1/1vESRav7IFHTWSCAzoKmwYL8xQVd8hB/6lU
vRLlE0G6x71b1/VD10yjqiEjagLtBqULIWiYyx5o6TqozOMuF8yPEnvefCBjUHYmSPyDGY7Xb59X
hmgtoqEw/ozJ/zF3VbyAbiGiAMGYcR0AKtqgMQuN+zXwIVgwiCiwiJrpLH5Qsb4Wfdinqq+5krSn
2CEFsFqYp4/BolcVn/jp98R3L6woBk6MmOh3XAdveODj5rzfKyPswd35LMqPLVLABrrO9o+m6T7m
pbqTMiGSGXzx1r05jjpM7G8SJOKQFg2KyhVT02XT8KMVR4j3q1BYF+7Dty6FGkhEi98YvGBkkHTI
f/RvDeUKuaNBK/I3jSPr1ioFbfSSQvQ5syM3OaskfHmSzF/8qQjnYYSjdmwNIXUYJVxvT/TOk2S/
oqBpa0HL2fEKjJQ51xo9ad615wV0sV2iGAzU5wAtJA50eTzFb/PuI5jX9Vt7hURKQbxTE6IZGEjr
xaV6zWDXdxguOExWndQE4E5tuxDt0OW+IglUfCkEbuERSe+fGDc2V7ehjgZtrWXqEFqCR9HuD2um
M7U7iprOl/6n3us8BhTsHagDlmSSbydOZgVofj2YaXHfXpzT+djT+zfEarMOe+3qrEk8kchm+t2h
Bu/pW1fL+iiagOdLyvYbZbpYnYXCZ3bPxbbfLZlnQoIaeZrJzVqvuGZEBLntCzvpK1L9+OIttR8W
/ism6BFSDHgPIKcYt8dBA20R4upb8ES7vhuVJr4E5KWrJz+4phaAt1kcSYRlzEgabmmp7GOC6r+b
fGrCYcugcVaYAxVscShu4LKBDrbjOgnKkWoejlH4MK0axpZrd7J2c09rD7Cg/Qdc/7+RQx/irAtV
WVYXO+gxIpKlZg+vPvzoP/fPmt5YDhTrtbF8JMEI95y49qjQJb7dgeLgbUO7wLDq4o3tHPrkxdVe
3/RaRLEdjHYt1Lp5aYo6zta4uvwyOqs0u6zE6nfYM7dCrWnj80NGvZZOPI8TZj21tj7kff7F9kUn
EwLvh8JWWkfC0bUPUUNrK2n+mccCG6KpJ1cJaDfOS3Uxt9a/Gu4KI3Nz66R4WqX/2y+Rm5k/0OXb
69mLk8s3e/ZEegvHCaXpiGtMM86Wls9H1PdJrzRjG1Ze6fOiRpoYWDcRgjwOYO9HLQv32F8I5VGw
7qsnwVHFOUhIANobrdBx/3AZSspBz+GDlu72j5+s0tx62uIUgVL/zjkdNINTc+46OVqaWpraO9Cc
K49GqZwQjM7zbrXeepYNO0hxB3wcmvcINw9x88XvGXGfZVpOAE9xxSTb1tWYRrD/LtAFIVDEu/dS
uvegnuJV8EsShmseW94lmQEgO+8EVIQVv4eoPqva8LBJ7h4ikAqHHaHF/ZZYWfrCBOJKfWw/yCVV
+GDIfoW8KaygE3rrDHogZ2O3JXCpXrQlu3bkEanfdnUHuHh+cbKNzW5b3jbT8GgBdH2IaNMC9poD
d1IzPZvob/M7oWhG0lF6I5HE5CcT79P3LPh7ghimzFCova39zbw2MuaKwyxNtlDIIkpUn40G0sMB
QoYKoUJ4ayqUe8QGYfAHeo0FXlKXj7iii+svNQZK8XPmzdWT3i9eyIbu607HkGQ3W+fIc+KYSjxz
z5gJG+6d34T/JS6sC2gX86vP6zJYylo/9Efb7z7xkbeBYA4tMHUtoYCVGS/s1AJVtZ6njNAsR1VO
WV49ACgdGxyx8oZljY2gPvxtgVrUyH5sOt6DXjYQbvn6cXYg6uXeqny2CSD1QFlDBcjHiaAe0ezZ
qs1fC4Krl7I1NKTIRVHicnQvJ2BNbRXLGGCwxIOlvXrqcJETG1eYXaZhATWKp5DGuEFRG0TebPw2
wE+t4Q3lYymZZPYEKICHCnM2cP43pd6yzknBE3101g65TjK5DZjmnoXwsR7bXNnPAKLkgxRb9jW3
oQFyzIL/ApiLLbLB05kR8rrIx31cQ2QgsB9NTeMJ5gehM7daei70QiJ8Z1gbjhBkXlWof7vyiAv4
8L9J90+0eqQHPcFKk+0PxOZFti3a5huprTBkUk3YiZj9Sj6lczIKii3soOj7PzaHXD0vxZdvDQcD
5HDgRVqpF0TWlU6qWl7ssPTphr+3u5fJda2MJxEmWFUztsmc4O0CP0LR1Gf0RMRKjr5bRl2/mFnG
SJpr8MH0I1gyX1NTtMVnTXZj6jy3nzxT0dbYGfUenHXJ9WazmEl/2Uh2+mBWZ5XfCxHKf2A7rq47
zNW1wOc19Y9oL22teosjl7nwefNhRpIlgHYV8HTy7t/lMdpY9yR7Xcc9f/fzxxJFmY1WaysRyRcx
3weZVucNzWBNBw4v/unsaFkdzNS2PeFXiCtPGiIVoEIFcmIGtOzhtWMUjzhjFN4WLQH+9/7XYc1y
MQNHwfO+0o1096lLSirvQGdNQWkPHmrYvPKKyqFmFAOlmzpwa3sNLLwtf1BaC2G3C1bcwLQVb3P/
rWK+aUEMGhX5GDMk+xMJO5/OC5QoOrGa1fJknW6CVhRKRTmUdnjwLLaEe3bMuBebwgLac4kmS90J
n/iddDFALx214I/JASrFav61+YVLLlwizpYNITkYJ18c9Iw/EI2J6cIIQz1/+kFEHlY/yBdJuMxc
4K+LLrcTrSTUP0Hm5avBuEo9OQ+LiVzjZ9MTmAPBjw0r3OUH+CPS523T4b2/loVQw1I38Dz/eI6+
val6ljuFU1hOYtfF9+kJHgXaV2w02/ZC4xPFNP5Eo62rDakNtUNGi71T4BrI/QYnF03n7/FdXB72
/uBcm2e46uRXXLPujhtzFX2ob6u7RyeOKRHqE8lHV0sBltAtCfsJc/0A3KJLfhPEuEe65Z7SLM18
0OKQWq44QsvcWE3tEbcEqJrqMq3YOi6LpyUlbVf6a2fhdbCpUah6oy7xreAyqOAVHarwgF2nVh3n
hqdIqT94hAsDPhbk/u5DOo/Y8338D69FuRIeHxnHvJ8juRgNJ0i6C2nHikzsThn6DEb4nTXpNTyy
WoCxeooLj9xb+7nPZNVsguLXsHo9p7SW1S25rxbFiRt7qJlWE3z6j1rHAAuOICNQ/AlyCyAav9wO
vEEgVfi2PemD3wlHz8Zx+qSlOj+5fY4BURk91MGSzs6/RE1Cks1WoXe+6lveJF2PpRzj8MhVjnCt
axcV+JsGqDdrm1Co4JatLB4Nx3BWNNvb6mxtju3fIvsiiiGMDB3wDVSixiC3jbUrSG4nAd+BeYvi
1T/3q72sSxvWL8u/0HYPaiU7atYpGfUNX4DA5xadBIZJOyJaP8r+FPbcOhEQSqyQHH1xZXkTSrAb
wud3+slm5MmGxcKZYToQZzyXKpRxcj6kBW/OCJ7EMgMKiGhuBlTdJGqGo+HRlIuoVpOfQwKo4AeD
X20uZRpaR729izvOhuBOJi+jLLbFWcNREFjuhOZQ6BnpPigfaTOZIHE6b8beom/xYCK0Tu2GKYa+
z4fDz4sOoMV0wdCouTtpMlVsCAozmT1zTy6ttDoXT0N20E5paLhztEZ4mYncgcWcCXNthkfBaavG
4v0hVaRX6rzv/H9bM/Urz9l1iv2UPOziXbr6RXKUyHJA4nHRVL4KGTOghapDrHEoCJKF9IaZWIPY
sHyVKJZ1GayxrVyVv/uns6gGabuPLU9qUWw05DN4Th9Pb+HAGrxxxrSOv1Q8GD82m3gbNjRwMAE0
daU7NnbcZ/BgltJxur8Yvr94ItUaQIdHfcvdVUzw/HfCTs1hlEmd2VEYHlI0tCWBd+HhtelQZjL1
QmbB6A7QqBq8t9ru0W7R6ZQ45VZOaM8731rkHj2BU3yKueYuVdjX5mowPKeZY3B5ONKdqsRGv0ot
1kj8SV3GdxEQy3RJqjAGz3j9YX0LGAJMAyMh3rRP4bqTFgnDRvVYyt4G834STitHFqfluJWTwzWK
8niOkRYwfYtR5hBs/BbfYcTwlS38cTIZMfkfq4ocsDqnex0gbXwEDxNPLRhGFUwhAbfJpzoju9JX
e94Rh91c116X9ICp8zCY2hSGTENxmo7bgqiNPFqL/4PTMx34QN3URXmVqiJkzzQnLQseSyLml3bD
bUHYD8mVUKGIhiXbfC888GR2pHrYvSmKLDaJm6wwU+S7aOmDkXPst+JTbDD0Wd8XU1naq8X7AZHn
wZiASgg1e5m3iC3jSyDDk7vu6ZL5r4osw0GybvC2lT8aTTAaO6Qta06ecThFl+MPGsYJlY03I2ix
t8Zm7G3Gb+HI1gs2XLkOn+Iffw53UNhdJWN8G0mQO5HKEK9ulRpqou5X/vjqtX9fsZ3au1w6O21Z
gB2qTvp3YEn9RXUF8x8wWnW6NR9m7CVMAJG9OZH1ZoH5QFrTC7//4SUxpx5A0BQOp6UND79IalcS
S8ebsvsLvC52tO362alQbcPU8emFdjvU9jjwMZp9rwhbRQVUdo0aNR+r6W1LWP+73UXtKosDqa29
zS6XTC99xYxji7ssIlQMmcZPjzq9l70p60+xg2yEP48/slDzTbCj209J75uRyhpaYFltlTV4Ejjh
yaepeDh44d1yJ5+HE1di47Dvv8gpeuNVSfRbwhh7Nl5tteOfxuq64l6IwgYqOXUQ0dbDC9nOMyr0
NkFkAdPI1y5o9txgOucYnQ4fGTsn6G8FG3bUTn7PEeiiSSFAVkU6ZvRKtkFDCui7Ed3auhwIie8h
83FCAyHMPDj36gFMG7iE1yy3QCA6KN3xKMv8PWrssw0Xm/TK8eP/nlY98AiPc0k5Tgyhfx+NEv1O
9wytyDKkltfWvr+TQ71yKlHOhby/0VkdQ8mOAWD+nkW1pXDaCaYFIK967zkEQFPs7joLnsi1QhVs
xKPy1j0fmjfNDXUEdusyIooXDaTy01+wo0QCb9CVqdyqdoUBHeQTAKsA1xHdoLaeF+DmYR4DfNCR
4utvyWj0fzm/x/Z0B8JNKugoub7Rj+Ve+aEgIpxfzOyHVg9nILAr611EotT+7o/As9KsLM3Tl8gb
/y7V5YgJM/h/MirusCgoGb+YKzR1DEBtAuzGjO7ynp2SwrjoD7e0KPotFumvyPTx9oGg1IklVL32
SEcTyemIrgRmZsKz2TrpkUEZ2r3aN02hpgbc+TVDcAHQUez3pTOm0pG8HXk9Meg6Q5Ol+JkEJdU2
rg+OuKomRUzYqwOGWAl8ry9zvKagU/iAEPHA6oIQhJGmBYiVQ9mBKyZHIVyeZbOc0WwDROyc4ZfP
xEZR16YvTLRmkMnqNbYDYmUwh1CymnwA5xCC46pqQ6J2wCnBPOwuCGEkCW7HUWok6DtyFx9yTb0f
bWeMjDLWVd7cD+4kM9XPoCAdydAcLdpSAVx+f62NaPX4cNnE52097YkvaG/ggZVIMnljcOFRY9WC
MlNh/Yc+eRbm6WCCvqLaQpj2RDAINcycCH1ZpRnIVTGJyKjfBU1kRpQfC3qSLNNV9WjkiOE1uVwN
YgHbSKiVZmz25/DJPlqBCQtOj4tmVb+FgvrIOAyBFYp4Q9Yzw/UoqAK18thRzpnXxR2uNyzZ0ZFY
+j+vpltTdJ+N+YwTLiTjLfw1q7vmYPywL9nxFTqQmUgECYM9vpGOyDjkHjVGDxGfCS9O0MLqoU9a
vTYp6hd95pZnlgvGAg0Ge/LKhdVWFmcWfrQEo8VTsmsiz9uOD1JoPXCZdHChHqLNLtXPIwtNvhJs
ApuwX9D4yq9kKXNle7QEfZDMkNbRtJrIKoS5V8G6G+sC4Oo4XOzASvHBL+rvkgiuRGgj1g4JdHnO
/mTMDSEBEn3iQoehMS8RzTqYr/GSSJ//1JjezCdYSXIwBZvUyM3nxjl8aMurABTEPbEuQ0LMqtkw
2Xpur1pQ0mCkn/mLLLUdwI5CsctmGiR3FyjKuWElxW3mk9xVbeIEvcPF71yrtpw20IZjNzXidd9m
7AhJJFqs1rO5ov2IkjJ0VaMYHT3fBBDc/JSRf8q3g8doo8vMsyitbyA6wFroar7CJIMqU1FSkgKE
z58J8sCYLY7NW0myDNtuiaJdVYQX5Hd2ScYyShpAvhaNnHmngQOp6bROF+W6F+GtK9MCe6TzlNfs
bkW2508gBXHVB3n1K8A5xh36gF3dgKwNLCVuBn4Q0LGP5Fgy2l/FYveOehFH9mLYEMElNBvwpj0k
WId00X/Go1gPOpK3PiqHqa4vFxRrdukbzLqGjctgSdmkJ6A2oy0SPI+eUz4FvN3mXXrqHZUUMo31
dlfBKxsKz/WZ+oMX9+dPdg0scdVZN3CNOgyPZWMSwnsEU6IAumYS2pJzGsNAag6sVJ+S27JYzocY
nqiZ4M82XYt7EwNOE/Pj/SE0/VJekitNGczeqdYHZU29JVn1VcGoeTywAatcxVewqVQVRK0WwSSF
Ya8kKxqHEATFsI2cx8H0F4btKIegLEWTL725T6yWoj0xGwrFZ+Itzr4o+Po7r04hd55zFBlfeme1
UlGjbrjRawB1OOrbJ2IaNgp2D+1xGu7lM0nBSDZ2RzhjbO53mO9rB1nOzYeUS1gPJtRQf3ZFg9X3
r0uSxVwaCGwdBbuHQHoIIIAlK7SRCwxiJvhNzrXS6JUV6Xy5o/a1ND4nBqd2mnC2bFtEwT8eXb/B
lKdzNH+jeaOt7H/coaYlbepbgvm8XO1caXvmqqfQPqm2R5mM6pmgHbL8PskrJAjIqCFaHF1rJO+Y
ckc7iZUz4QDOnLlszwWOtl7cxv0NqutVSBJsOIG9TK0cQF1dck03KYc3npVxR2Manm3zYAb7sAd+
e4msJnyMVpdD+Gx7f/8C7l5JaN75EzBDqEOuAOW5R7zcDTKLrlXo2cmVMSaUCU+ORRyJRozfXc7k
/8xOAHuTNsmfTQh1tGv8CDBIQe9qS5hpEbodTcsoO60qvIJKkT336gncNcE+59assBB3f1p+5Ldt
QxqL6IHJ7pjJhJj41iNzwW7GoieEWsWgaaT0Dkldscr8XxR5PtHOz/feSA5RfOWsPUJkBpgtXD4u
Kw0ys1Yb2KlMuW2GluwxQ4a0x2HIrsBgVhn6xlae5d8a2BR8d95ibNGEWrrOGpVtQUKFNq1Gkhj7
PXTq9NslUWSQAuo9/P7WLMZzx8ItRveEy0DeM/gH4rERmPReL+ACirUlX3IjwL6v7abW6DQnAmES
IMEODSTnWudfMtgd7dQvMX5EyBYFikTCGzZwI6fu+uztNGptVIQ8mP0mZ0hN7wQab4uWOj/I0Hr7
SRCJ0RG1u8xjAPfRdly09J0FC0MKTLPeE4yt4oUiETemS5DGXDQmhMj7aREAl4SPpPon2WjxUHMP
JRs7wmaEUZlEd9w/rwq/Kb/TtjGG/G3zBScJ3It0O2yka0bNiVRXND44rydXl10CuqIrPhJAWruY
nCEMA7XKZKR0Ps4d1X2pv2GgiAE/1y7472yyHWvNHqYg/0Kg4BXxl7Ely+aMt1rUMd82eSQoPsE4
Tin+aJYC+Ov8Mfstyhm0/dd2P+eASLKQ9XG4p1QcorEjzYtR1rdxU/byuadcl0xLXqcmXNRxAlOf
xsPaDCFVF9FZp0ZO0rOvmG9KfcMstySyVdLYi0LXcfSuWem2KfBzmHtUlPeP2EFx87keoBbFzGYe
CMPs+UcJAvBHBH/85CCQT03WaGyirKQuLyZrXaZayNUQSzl9xszWzdVyEmWBwkvrOFedV1YGi+gU
5ENoB6x0BRLqeMVy8tmeUWqfkk7ekBxtNKZeXjeexGtiSEdw9igwiUHYlkTZV3Ua+839oTfm/Ecz
mr/yb/A/G8dPHa5zpDgebO7TdMT/tYz2wxl9P2m1EqShshopHZNoVOc48dfoUClpn19obPk1kJk0
tFFDwJ1vabIZq5FXTph4ECKVHGyAqoy4ag3qo0wC/3T9JdHifkFgHelSgk3i50v2lk5J9/R8Fj3k
Y/so6YG35xi66+4tSG7rwb53tqxxUU0qADOi0D3Px8GGHjvbfSEYgEYOaM1yRWhnrR0qE1ypH+4B
nShqj6xd7Fm4j0oj9WB+qi9KrkCXJMNf6c0Q9O8zxlBwg7ZfKZZ4E1P0pClUJuGTIir4N3FAdG4c
I7jg2qucZ1gpE3LG/fSgMr3jgp/4eRhYhRPWow6rq6Mh7EzPa0KL9sMXIljj1bDhZwp5Jhp9yQk2
sNU46z9IMHM6sgRsDS6ECBqfVt02Y6qwQEbHgFGQ5GmVC4qOP7dwCFoTpceSS+QUFDYMl/LPMhp4
4xRlGbeTtNvHNTSnLXlkzuod1f9DSmLemeC6LxTosgyjYn7Xf7DnrLnwXjjamCd7cIaksQUaGepB
bq9//nLEI4M1nXVGXyasZsovnZALc0i6cIglnAebo3C995SWlIFpHebs10bvvKN8UQ2xSR7oWoim
H8sf/xdEWMDX+FhuijUAOC1ZJu7gODU9iPLgePwanoAeFX/IsyypuOLx5fkaCs6udQs5aufLnOTN
2TTja0jJQz2ZuZ2+nbLSstg2ZSAeFsIQJrEjevHb9F1qv6zqUuyWGk6qiu/oFkp/QmCeI75e4wiS
B8mujPzMICX8svIrr4liAsYdybR+a4R0GNcpxpYYP1PvPF0IEA/s1JsUirvUVKiYn3HAI5BYWpDQ
rwn+SftESb78/DWLfnrPi6Ao6nvwAyJGf1ROmeh5lw9nAWAeVNXKyZhZX3FSGY+C36o6V0PtVyM8
6UDmF85s5QOYKLCh93/0LQJ2QiXWgi8iuLklOlVZqiZMITQHy/9mGXc/zjOyLGhn+NHzCEEIm26Q
CVVp5+M/yMFbjpYQFcwJvlbO++cTjqgZVDODqRSqGlYpwvgv8tnBe2yHtCFU3W6RRiD1gsamOjMR
iZtbd4vvE9CujnMhvIgK6fvj1pVpStfYNiKaZQksXB06Y2UGtVTl2C1K1rSYdDtxzK0R9G65R5YY
QpbQBU74ZLF7kUBC450PLGi8fLQK9evxGzsXqU0trfKr2MJE1aMhPR9uKO8bekPErbG/FE9OsjOc
GTzFkoe8VMKUYhmPTjQ2PVeKPZLK9TMDHbF66K7wpyc+wm3UBvWYPOTbpH4YF3ZqfiBN8EsD5Oga
920SnRizV8hb10yvso9x/1hob8qh2D8yxqvPPOkccPFHgtWAOWIHHJOeeMT9I9GXumLgHXACBpGZ
y1uT3hm/16hUKSxEo8uMteJNbddnjBNTeEoRKDCVhjBwwW1a4uHHZ7m91zUCQsEjmcawXopt/gXE
W79J0/0Sg8AfZGtR1b3DDsyWBTKbz9zBh4kch7I38L7n4aGc2MA+XHhKjlAPz4aQJff2mujc2svL
Yamt/VLkerzt7obogNkCLHH4057zmqjEg3jZhRyd9CKALv4HLo4kYec75F8Axd/GdOh4bUsbJ5ya
Jd4VPRpBImbF60dnpCDasxvNsxMxYP6Iwpx+oN8PV4yGX0hHK1rEft16G4QyjpOTOYIUPcGLep+R
pVgoXoMqfm6zkF+JzZatY0+O3hGbdZirMKv8bHtOu5oTfc/iSjYWxB74/iJ1sp1bdic3nehjtQLI
xT/KOX2Ydlh8xEsQniqtbpyaTV6wKvXsu6xgS0K+vx4igjE791hgOv1stfI5Zm+q7eHdteGlll8F
I4xstoRZOD3ZI3wfjrhYNHJ+Q0RXUraeZJzqq8RvdvPGtR1zGdT5kEPLoOWlC52IfKzDnmaqeHZR
vgqLLSkXrMvqLST2OhQ2eR+JWvfjX7rhAO5LbECpo1a+xvH99+yR2BEz7eHx1uDVgyw7F+BXB93i
W1mVDSVIBPDfGmafgELvrfcGvPdjz++9cjZQcJDUm2jzFCrNwuAUwHeMZu3/oBf5XVJCKp5eSfCq
BHqnKreVY6slKSBCyeFcJmQtSfM3BJy2g5RURFuHxrXaBoomwIg+ajq0aZtPFYWQACdwUhJ6Svd8
eDuJQ4nsMTvm4yMGh2AsVMZQlQ6otmeRkjhUiTa52qwT4OKS8mirx6sbSSnAta5hDhEApoDZKH4r
pzuX4chZMw7VF6YKH29BiA2tXHUcpkwxbgR5fG2pn4DXSTg1j7JEw0+NOmS7Icvy3IlZNTSNpiqk
b1Dasq1ToHdf0zdgC/Ad9nzUnej01U1KVfOV6taVgMpfGP3mb8CIFGx/sBtbltYBpIrpjHes3FtA
CqScgf+MhUGmMxCo2uWq03C2qrAbgj0iYW+Xq2mhMlI6jF3bZUP7nN9LP9DmF4JOcBhh0NkeZ26t
MYEhnECPimwCQfglLFQMKVKFBEnA51iiDhtQu3CRmIeX6TzVuHP27rpmDBcsOHHpjOg9iPEmgEqx
9ceNztj0hYT1Rv9h1Yp9D+LmeLNh/q7x/dcJe+5/orkHsZ+WpE03ZByYwuEcLx8TUuHdOhLHRoDU
kgGNLUnYIBRBL34lSOKy5KNUAZjNSqzftB9VniECAT+v36Z2NOh0Azaki6Hov0KhyTSt/2YkKjxl
qFIz5/jhvf9WuHfaiFQszDR+iPFaX9H/XIEWpA+KqI85gLUqCj1qzYsAGwoEDSc2o4OI/snskdL5
21FZjnV6g6dOxBHbRcfC0caGf9ZzBtkAc0O/2kqgz+W7XAk8ymrRRvQe/uc4Gk3OXTMzlDgI9qCY
TgdYQMtUcJIzEYu9GQrfEbB5brImfttlGSJReJR3js4ZWGyZ09RQdM3apnj2XOdpPoKIMObkhNw3
kBVz6c2AyA3arL8LLLYQzNh2XdfBwYnz52YTed9XoLHVpU0kaLqWIN8N71km9UnvAivPGLjNK512
hAyakrEkSc4NosZSaxP1oY1E5AOIqOMpmIA7IbRz5pwR6hiee87TazFrZZucxRlrt96BrGI8wqeh
QHRQ8zk75BlCE7QAThjzIZ8f7eDRIsqR+bGhEjGb2euoGT1RA07hjgxvJRqbAmIe6HxhGYSP4f76
rsTsDpWSECkFAw1flhrppNNRhY13se5FOz7xaWz7rZIUGffqh62c+lFda0MfxD8SVCaF6mOuyFzo
yBNKf1UlSrA295fEb2mbfjqnK9oYSznwXeOXNDM0JzD6N7MKdrNIYkplbSl2Aly+lZ6Y24zjn7ei
2SG1f2NTF6VSq48a3rRl4jF/B+027IFVDXEFO+skVAZBa86XKEGm/Ca9Tar2hOu4x0++utsdn8ek
V/00L/qnnZNRDwwZYZgPxeOGYF6avy09uUwhTOds8SlBLYwEeFMRCvGKV5g1zPBF01Py71CoE8Tg
9vX58Ld5cfDfAVuz/1vsnXWDzTI+69c7VmUoqY8rAbJbfkbTqMobT9FFidG4pnTlV15/V3c4RAHb
SvXjTCc3GyrP3PeOooU2FGoMmG0Qhm1ARmo/5FKyQ6TTEfU4k9w7a3sE8WeqL4xMysDphiZKp1ed
aT4vx80APSmZxzIRgDPp0wSgF2X9T6dP7kwfCQo2APkmz7X7FDM10kHxlodVDOAbVgG5JOBxsJiM
DFAi4T59DpOGMP+wa5zan0pJ5VCEKvgGebYYW9yJXwku3upVztmkDiU5oz/L091MVls1H67iUvrY
2JUvd1By21yVer/ZrAwwfpTIo4ud0nKNTtpbHeY+XmnXeODZ9FXu+bZZ0QTcSwNdI1qRZAe9uyle
o0W61Zgm/xH963wp8OyQrpVKqFXR6tP+mM4sH6E5/dvPflEeV1jFQq64amJMHKuDdGOA+0kY0IA7
TctLpksg+FprWLytviuApT4Jv1rSgsQX1mNyvMYIvQKKD3p5xP6nu8btXF/Q/BKenbxqafNfiAor
IujkPqAa9rcUy8Y4XCSbUdBZwbOkShUXEommoCasnzmAsWG3Uz1ynxI17M1PKXn2PlvaoHdH9gNk
ENpUsHyBSFGemeGKqVcAifUjpENVf4c1krAe4XTQCVpiDGAsT01Tx9vaJR1Hj6PVqq0pN4owtjxK
Z9yNuEvlZpua+K4rzjI/Gcc6KHW0e2LBpFn70xI4XaV9C7gGLFOrSoh4M9P5VwQssvvhXjZeTjXE
gq7BmTbEOSDsl88DYrtPh8Ms38HO7pPT2wthTZ9Iu1HOYMbSQwcy4qYwvzTph5PyflgIOEWDAdG2
x7gtSFtbHJ+n0tMTl1WkqZnMAWDwsOVpTGH3afGifvRWuEw2I2k2gTIcKlBKDk3jgBl+KfMnWtGM
YBVu/mjej8ZgSCp0w2yN7dY1QVguBPU+dzISVCYd/0g1k/egcj8DaeamN+KHGVd0bMmuI3/eJn8H
e2XVgQUm6iI9djUitN8aJYJSjuJvzZyIr6mXWzUa0VQgw9PgzqL+d7p2hzxCew1axuhhPkrBqFTE
H2WdGZLinwU+0lQLUUsrCq2hr0p9kq0FWDp1jt4njzB8yPpxk0HexQhBs+Pvg1dVwn48VvLbo6/3
jwTPkrLMRboIh5m8jb78OtDtjLWuw/dB9rCdHnIdqyxRnQ3UVhhSLhPEKj58/q5La12jGRy2zy0W
tye95OxP5JuTkNKajMcF4dH2XZcw+BPb7LShpVmN6Ox22HmiatPeBgVc0Jy8YISseGAc/C6aPoJ5
YDOolQjtpc5ixnk9oWw1v1HM1yElIOBIys3gLd8IqFXBbT6x0xM6b04OF4czAh4AXPBm/aJ+Uiz1
xx+D+pYgpQfrbzOhzT5gGm/TD/JTQbXCEnkuNtDGAnir/lfdmK4bIY7PJqyrwJjBkr8MQ+BZQmL+
E6Pn5vI/AclMj5X57NQ4dkeQ3cjKr9n90iMaCR5E5otFTQYaa2GeCE6YTwXWtQAXeYPdmYtE5T5m
GqruN0UckpjN2QX5jDYEHVafeI2ZO4mHMtqkemJCtGNYzM9b+qT5f+wqX9YU+uWdobr+XrZ/9nDg
PaGMl1byYxMKgF9hMJgbmsvr7N1oEEgBlRve5ygA+XvI9XvSwBc8F00I/wuHHzloWdBYcJcQYtV8
86hKt+oAqlF1cJQcf5pzToEVQj6NBFy/VQACPlTPR7Xz6b2XyNKec5rNUeyZMxf8CYfExtoJfs3D
AQdEJhHNWUcURMg6zjvbpG1ju1p0gKGFIpqU30b+RcsjlDvfArZRLfQrKBMGNqGEBpBxjthYKSoC
QEMEdc++dc6ukjV/s3VlmoJekh3LECw+efDZsNVCT/uVdjzbsuq8VUR/JrnHdY9HdhdLQidzlQ87
k5s46rxOmwY3ShjkTa0gBUhiWTAf+pnODrP8IXY+ZhLZH0n/BnxHst8Qlg+8BTpZliwTCuSPOIZd
Qb1nHoBBx/N+IKmpWP/G1wyQB+nioQQufCBfkyHmdRk+3OypBdROMG6NpgAoPOYLsPTOvbmBGtmS
xFuByCQj/GGsJEaoalinHGCRBZlaWnmSsIasEfQ/+JwFRBB4f/VuqHAimAfoBPOhO7DgnAtVcYa5
moaXdzj9jKkX5pjMW3unkLNTP/5A7Pz+HxpKbZwgMZXWEi+meQY4DrUoQEyZ8wMuj4XbkNkepvrN
x8OmhcbGBPUKXRvmkkP2WXpTTR+KFicIwTrXWrSUDt39BjTKavhuVaK3iuyeGBRxwZ7ANGMJ0FVl
ws1+bYoe4SK9F492XDYoYFXtHs8D2uH6DnapNAucUzu8/xHr6iXg7L3cFJmR1JkHjpbSEP9PSKlA
8Tz7T43tLO9/D5/Ket+H8F0ihNo5FMegOi/Z1m6+x+FUaJpaM3uYAVKlV9NXo3nHrj6CpqNNmj+R
r8Vjb6kfNj9uxSejucp6LeVNVP85zKV6xCK+qKEnfog03237QHMTwcBrBu1sCiF57rZvjkzy0XBj
j8bUCJg9bHRmjpPgo3P0JHGyi/5XZYWgvt7re4VBIoLMGkCwYoiwBY2BQKByc12gwUBTYA/6MKpN
JJ32G9wTScBGUmAZle9YYFXiITaysocalGEpUt5RDzql4ASdqdMn2bQYiubtPofFVqEIsZhYWTJw
cw1rvpnpJS20eAwPNjNXK0y7jbibKonUCDaptors4RTyjropbDZFmX73jhzFyU6u6SkWKSIb+xDr
NDC+cEQzJqKZDgiYO6TgpICZxUvoXKRWB+MlF0bkoGSGcUvG3kfMcMZ88SUxAS3dNM9RKUGi+vJy
vYohhtJK0lNqvX9ijknbfMbqH9jlz4dMI9Y0glNcw1CXpYHo9BXE2bfVla5nwq+oD+7/slGwMym7
ZGy6+lU+njbPq7LoL41fIvIL5FAPZFGQKMxVZkFpF61TMv4+XscEccn5IMBPMvHO/b4hMPTES4LB
deqTvOMK4ZmL6I+DwFe/uFxNOnunLEeN7SyN4NDu7GtpXFadtGpGsBKq7kx7bKWPph4aVSBgpY5K
kn93tS0pR707KgZMYT1Li3VpJgXNDSnclg4Z7uf54QsbqlFRMcdhZh6Imh71GI3BO2sMqaTQUnUZ
A8Mx8989Qh+HZxFTbH4rcBgsOK0Re+xaakgjr9UtGYaLfBHaammF0J91vSFmQd8Dpi33ujXr3AbJ
x6IZnpuDWIt68bA/ER3RXk7pO5tzskB5XokpEkzTarJeWwtitAYOIiG/WLeP5GzNXWkQEJG3usjx
MDKcp72Fisbe2SJ0GFk0sXVdXMBpmbGORI237Qa4/Bd9/Vc2aicdYnpRI0iW6/StLXr+XBbvE4pB
VwRY3lzMy79naM5PaL08KqcQJfCMuJ4DIBqDA3CotFgxzeYiAba6Oa4RnlyJj8/QSXaXadnrMCCY
aFlYctFi+EHtCe5dgcX4lGzbJiHlrWbEEPpzCgQz6l8evhksCf+ZHLTvf9hwhKVHOZz3j6t42Pdk
2ZQUr6EBfJ+IW/5KI3PL/NpE8NLl7PW/xes9eZiRXLhJ1u4HRNa3Wlpl+Z3nZdflO2H3w5DUs+dh
+Vo9JbaJ1aM0K+lDckW9QsIXHfK0CmLKa5rqgV9cxwkgvkWoVYZx9/mf2hob4V68kKKk1y6gvfgj
/B0c3jGFyfp2gu07w6rBQZDIUAM/X3FtW9OZWHWJxrzGEYfbtCWKJfE5BFswt6oimNjJ/QA3/1TA
bqmTnbF7K4XD9kJC/Xg0XG4FZReGik4KPzVCn24IT4tUL5JS/YyuQ1D8z20EN3cRxmasDIca5mrn
ZeKY7xQf9VQ+We8C9tHf7ZShELpS+uyO2qY0utjTjUc2S/JgRUa0lc5XlHrwr4bzldecCbDBDh9z
QzL6km0+O6tHNaPe3qaAPKrhEXy2pyDimVAiNKttp5wnvZ7z/VruUU/o44uaNBE3YL2Q6AngM/q2
dl545xtyhxTIJ+uQF/8rIyQNdyaGk0HJ7Snj8VtVpeG/gQ0Lcp9F++CYyAJNKe2nHSMZF3H7Kbx4
L+pw8HRpKNqwjj5ov6J6vBIIxp1pEAeDMhHqTc1oFb0m21h3ijaPvA5ug8dK4o3auvWgGInmoa6t
+EHkB67syHPYpnyT0us5TMxOHA1Xz0Do2mDB7wbaJfY3zUpldDTEArNZxwxyFbx1uKFGsliygpqT
8gkL3zHtbU74tpAU6CXgLLNv2a9ICHy7gQcRtQZzwHtneqblNxpShcJcastGeNDcxc9SxyaEO86+
xeQF1wmitQdpQYTzqjNE5FOmM9hFIoIIy1ucLnDVxtGayw10qZLKLHo1TsBCqLkUkvUqObu/3Ds4
7VTm4yv0gb9a+LB+qlGNfauwiI1IA+digsRMlnD37mng59wuhI9aeFMvxPBJitfjpY0URFLCB8us
eyV15PMNpX3+zZzsSXzm+KEJqxMd+dP0e12F6DsiAxXaOgIyo1YeMCiIpobdAGaN1pLuDooJHRT/
G3/kna2prlWsRx6dG9RXq2I36YWPvBQPVfMBkfp9yWdwJ3ocUTZaAwEXdFtMyNSjdFdXjR+91Dr3
4m9N9eyxMneGye5QpSZfl0lJrg1UZOEpk6e01ut1ZEIeaTBUpOfKEjyaUjdt0pqnnEcL+pbpPnhy
s1jdo6ad+q9sN/tTgV2tFaxsja4d37DCHf6UlPPPSMoGEXK89ekEMpjdp0emArW6Bbl1JWjCZG7i
fCINsM8HEimhT6n99UnmgebvjJddY7jIeuBSG/EbjJzf260Yc9QqCjdpV/WZMOfy0dKh9yyqZX8K
xh0VakiHXsYX7IQydw+Z63dw8C5pBw8rC12OL4D4HReGcObTZbI1YCkRNDPX/Eua7M2DZfM5vF3h
6tzxSjNQfnoxqPOJtN6bAeYyXLc2Y55ocjOXbbJUOCha3IN35C1eFQvh2x5Ou2eirbltctAmImxa
/SXHI7uHU28OoLh/PYWPQStd944pqhoXTLjz6vMNWhJ8kX5s5Fao1vgC/5AvurTKXzeedSjjXAaw
li41Dz+pN5qxvFbbf+E0ycaEhYvyX6fPbNAOOKw+TMCE8yWtGMlD+3Iv59EQeEN0329mSdy8ls6K
6xEF/FP3OBGeCdF8GPhjmOjl1hvyUWqEnqwvoiYWPqOnFdj//EaII5BnkDK8NZxpzk9m5KCvT8EC
iPPD11ew4WDGwFFa6i0dk7661yv52J9zAfkVW5DvmeBEEzyteCkpzlFCE6WlI+L7O4dNG3arqbyq
r6mLDj3i0VDa+iIvNGAV7iALrk3gVyjtlVqNOj1mWXOqcHEuhetC59/vfRXNlnUmH2k5Mw1Q7d3p
KR5ZI6wNIKueChS/i98wdv8WWGKT2UcJgyVFBNTl6O/odZQkrcU+RE1HdWVxdtEuGQ6sa17I9eZc
CkOH23FDShyRDkOdPuu8zwEpt4UiiLc3Cj/fmfE5RvOY9p2cOZA1cZ1vwyfmATGrMbR/u/9qKqUu
NQjX9ueeGE9Ms/AVHpEaS4RmXp1g6cXAgzsDDK1rKtJqB28fD0RO28UbI/wKvgqKQApuUdYg8ENP
XA8d5aRYrYY9oXlemRrGGP2Xxi2s+k+TgLRtJ3Ju+6rjpDpHhZAWTLwfNOTtEjD21Myqu0T4/vPQ
pMP5huaOyQKj8TMe+CS9vLl3YqSOrbyPsgK8a+SAqSbKCJhtIlsq8ABrmeEhlz/kE5kERW909HwB
b90Wr8/Dpu3+mZhx3nNKlstCB5KCnAKsPZpomZvTS9p+4Ci3ZBHqbqoWGeqWevqyo69D7q6U5Dfa
CcckLKhC1Md203ZDDLGyuB3LKvHa+VMyMgG1YscX/nYXlca2pLBAG6KkO7I92dm3SCwpLqDEy7Lz
/4CeHUA4+fN4ypCuuc7gHDPNcAAToczqdobyKBxV9SoijgypZnW4c4PiEioeTlDDrYa9EAHTSQZW
gL1c21v2pEiJFgDJGEmV71LrJtpRm10jIoruoA/41puEu37r68gc8o4KzRa54iZSGPuPbuSJDjqY
wOHYL1fhzU46qyMNKeb4aAboyIFmygK0PfJU8uQKZeLw9/OIVA+mYvLwTyumSUOnOkbtc9Mn4Rsv
p9WVCKs31KHSR5rrmUwKfTRAvdjStU08DkOqtdE2iAnDPG6frGrC6+PcB2m1Ub54u8YWgCQTYOoJ
eC0DahiNFHH58md3j+gSUV/D95OfIov4jKTIbw4TPttX8C3soMkpCSN7839X5JQU1bil5hxNvlZg
cVGhDjW2nb/R5zMFX8gu3Xc3OjIzSpTlNNTlawkfCQFm0HNkyl+JvYmWs1kGhKN6U6mZaeQhpK8K
Oh61J3Al4cNxreeV/xIwddH0t6fPkeL2sB96iB4WTDNkafNBWAfHqKyDRskjX4Psa0g2ZpdatKAh
nwZ/zIoAAgMMwvx/ufCHOOKHNOkCekCVp627LCIjrLvmlSGD+DIpUD7FL/gvgm1oli+GLH18MPJy
HbW3uL1pzJ/7gq0cQ76WDc+wmNMLxxM6KOdYHPOk5leyXWmbnxCI7TTKpKUEIYQrRCpd/5fLMrnz
60DKlzBvaYH6Yzb5RFd12LszUwbGY2/KzirV0XX/P466oq2sJe/+ve65zm/E7XTUtI+TC8fB280Q
/g04cR/JDIF+bEb5oaN8PXQ9d/eUuA/+P35x6ZwsB6YhWuq7g1HmR8azlYWKHbpCLoreiKwZsDdV
XzhVd5PTwjuIYlceuU9hG1E1zm4Lfoxi1cnyp0OlM6JvclKSGSidnA7PI76ccKlV+CNNroKmzT1P
B2c/9f8VZ1A1LlnvpK/9gqxsblO5pJdnhlA1KyFnJ5HsIyLQo6yBFtS9jN448WM10YQDN8iHkSO1
NJn3A3F+wzbpV1avPfzgQOZCPyWhccNNBRRYAdzZcsf9JyxB1a9iqYR5tSVNyUtUGzN2h1N/nrT2
f3nokeHG+u0Col7jKkEooKG4jNFAJ+QpxpGX/9WH8zO3cVjCV6mHV2m/VUztj0MLhCaCdAijFuBy
GildHKgmFPaX/ubWTQNf4F04D+IeRURcZIAkEEBhm2WO2JyO8ALf9wJz6BYoMfmIRh7pl5/3O6x6
EwItynOkxhMFIGuEXu76cFotlJUO5xvdDQ5JowUzY1ehv8llkqQulZ+YN8USZiDbVi1dkLYRMG7K
jVUD9W3pkoOR6UC7vJwcuCDBnJXCmvSRB2RYV0TVtmed2OnodTHNVYMIxAEvMoz1oGlnainMfuJn
kUqFqbzX700mv4ImqX4soECWNzmW63wKmST+meHH4NffpIQcy1Dv50spW2/7QzGhYyGolcMQuMq/
vN4IAa6Q0wOvrkvt6kr7i0jybAQ5ao9NLdCpMz9JuobIy97ZzlbaV4pmlmI3Gm4v5vf6o5twDWB6
rTlaNMk3rLHEN+3A9jZFr9n/wIa0WW7VGJUKg/P7/+Sy4Zd1vco4NjjN+SjBGogf/qeNWue8aJZr
3tPVpOqNWosLs1hGOUZ2fGdM0NjcPcvPG9rP9g5UGGtVUt7MlJ71WMcqXGZmv7vt6t8NS5X1LWtk
DlAIUO2VHaAg88OFYD40SkjaGG5hVDEsvu0V83YO6TzpNSLazr1ksmCqyuY27OUCH0JW+k5ruNQO
xZy/j5IU0UIfE4SYxua0yYZ2xHzztqaxMqyiHj4steL8FRLBXF3glcFp7HzhX8GkNOJYsE25jdV1
2b5tbsDAvwChnzFGfCtN+enoHiSNo0ehL12Za7MDpOXwI6mcnjrxUCv3QpfyWwLaJh/rxLQBjV3Y
vaqENBuoH9SFXCeQZxCAeDm78e+NoJlbyqwd/U3qVhe0fYZgEhF4xJjWeMTv0qJXkyIJnqPxARwz
LkoyuJg7ClA65k3TBDOmXT9MEI64OSaFH+tXXnAfxQXPnrlzqzTP/WQF1+/NABqSvCWGg699p+KV
T0zE6gQ8LJUlc2B7DyyTEUa8/3R0cfbJ6SyCatPMOvGjmKWydfs968ThgVi0iZF5BNcJet2yUjbW
HmQkUTvDKvtc9FCHMdoxbD8nwYJAxany8gDfI+hAhvE5RjVhgI/CnAiqfqm6qQkbLmeMv0SINgh9
P+uULI6GecDolUWV488WW/TCHGX69ngII2Wg8XSQdEC3R3aUDRiLAotxSkZY3fyX5pbVkmcAbzv5
uBcyZBdpYIWqC0+5xC3eH3SyKxW50LcsVpdWc4tLXcKDon1vp6vDGGVCi8mGCAbOovxJXgzFAajS
/+w9aC+gtqhwurUq3cz1wvwTX/qLl9lFL0wyrIMPadnuhQkm2dof0bWRii8GXBvBoNvxc6FEGj/2
S1fngh/nnAK/gbig+Gsf6SUe32r7XDE3+tCutbFBcRK3PMvslhECU/OKEOIF8oku/4/vBEJl/7l5
VEYR/kh6iQOhBcP7QjHJxrkPXZHkyEt1edMQx8zZp2LAR2m9mfSMTK0KkVfj6G5WpJGMb/2kBf3s
mU+3uq1dyRaIIljdt3Yhhqf7c5Y29D7B8px5h50KcHF8L23CNvdSFdC0G8dlE3DzWq8gKA5GE/8D
ELqRH+jvj4QEhBpBRsMovY6zpdS+DT/r56eBhvnd6Tm3oP97oowBbHZr28RWh5Pw1JuMJvRXX8pa
Si7mgOPSGBTBHCVGGS+wMIc9e2lQoheVDhsZ71fR66TuwR4f3CErJjSTf6IZZVG879y61XfFpLNa
BQmwJvXTFWSXrsqUAcqsWFrCQtsCUOwxJXUFHIo+774T3zAeRbY6C/6Rbs1sQbTes9WwNpBvZi1s
SE2d/SY/Jjk1dM8zaRzybZ9dAR2vTBfT/WABxE2AafTqldzv4K3sljZGhGqtrBGELk8bCwOMYz+p
YbU27hcxqLtuY8iZwhjbpreffu2H5UywJ/m4RedJ9FaaVtQaUuDQuG55WulEuZC/2b1RyIlmj9pd
x+D1Jt94lausqcb76BDtHjppnxrrkmAZRYGgK+Xg/GAQ3WnG6ExQ/6kh4JPDOM/1q+xt/B8OvxR0
Rf148oW7S2dIdufRCz52JJk0OIUgDLZ3BvCE5CrvllRhRYBve4dnp/0YZY4tR5TGuwJJ7ozx0pYx
xMB8LkhxBRqcVypF36t0TSK30wzpk645tf1tprO7TyVO8vUbxA0uWeVxkUUL2FISpbT4D6LADXz+
CQWSDZkdCWwMVQzPdu4GV5j0H7+bCgkgcBfZzhcpW/oqHPly26v9/QU9dUWtNFspJmaI7BHWnsEq
dtZ6TAvvtG0cr8wZlKVqf4xc5TI4O3hoNNuXzuRFunWCfFioq2cdMbJ1glQSsK2o1UF0M7b+ie/O
3MaTXA9YwzZBgcTadzsXKU21DNShAVpTFQ6KOnt0aE25Z7myEh+DNoSAohOAfh1rN4CjlcwJdPNx
YMXw8IA3y5wf5RSLI6nO8/U4eaUC6AYhMxF6c11+LINAo0PuSOKKTppxzEFq6mZm8I7IH94rL0n+
BuPbDpejdexrjnFN9k5CvC8Dd6R4xocC3EaKCRBU9U3UV/V1gU9RaQ2v/7+xXhT0+0lbiBQfsALY
CdybQvrj1FQCAFAkC+muKUOOxSIR+hRnNUI6Az2B8aL2YeQ2AvqPk/2OEtMmT4krBhbF3dly6HXW
Z2LilLLKY9tT2Fr1wiJic8M4M9X1VWgZIj1sd3n+I9Tl3Vz2BCTVcN0yREyQQTckor53O9Z6tW+H
d3e3Q9Q1acEw8gxbO40a0/qdqafvuoPVWzL4rI7qET+sH4sRI7RmUboRCWq0jrsD9gVYM2DdxGoK
f9dpjWMQPw5rcEl9LOaduUD8vIkQoHVDu2mbgZwHPRedmqrEqHXAtyL+Yf/Rq/GXBnSVs/K4xcuS
q+QgiIyM3Er1pW/Uz7dypePdgyQ7K+tgK/ReTE0w0jOr8sr0PHMvdG74iLeqRYclKszjz0Anexmy
uRvGtTS5jMcflS4Fb+5ntF5JCKObn5pjy2dElO+jcpUAnjd7Ihdi3TuY/c+nWqFKMHVrTKue6BTH
4PNramJPG6fT9msS/uNnkeCJLmAMgWNWlq3Wf+Z4XfqOOA1Xq0DR5T+EFvj55zN3oF7XAKvGGCZn
H3TMogO/TnFcbaBtouaYw09FV42GCdn5VERmK+U08yjdzqKJ3GN6QbGSxWa1I3asgfhBnharI8WI
uRUg4HtcoeznbdJVby9CDe+qzNzLfJS9y97hexwfJ3tqq5flquANszC5WWjJDygHyKXi8+17Asqy
q0My7uRfsmEvQnSjzXPM4D0a7r71QxHbkjazDPHpnAxipejSI38UJQ3qwH1XAcvqIt5V0B7K6sRl
Hq/HF1b0OVg44Xpn9r90VQoqia9UuqoP2n2uL6baDldulz9bdGxwxpNfRUC/v7tzH0P3H5LdoeZH
prgkED+fhJO16bMJAIFVqgJORoblvDC+tpUc4Zmm7uaPlAHHKaaNOCxSC1dxTpBLokX3KAIRk+gx
ENm42IKC+bR59aN5CkdijumO0NHZIrOp/pMPjFfFVGEHEpxrA8QrTROllc6OzuLu5R2pnhnkb7za
e8r5r33cuBedG0qqeUpjbE536oZBGQaRCieVCsMO9ZqMwKNOs6Fpu8pFSweW3carTsOv1Ag4mkSo
MHVgOdbeKZNMsVj/MbYQnEzYTyJ63byPo4aiCseQhImm5zzVruWKAWTGWV5OkddUflBBynsmjOb7
ILucHIMv54/Ms0LvLehk7JGC7cBJQejkBgz0Z4RZi8xHVKcG4CMTp/01vtewpC9a+oFppGthWrLl
4Cm6gg2tGpimpyWmvdCv7Blt85rIyD6xu/iDlqYagDEQRP3tG21jPEBI1A27cqjEYGZrxZNX/UV1
4PTXmssngIvmTYlbgQD1Xl00jiAQ72kN2HkT0TKz+mvQQUXdS/Xp33XS7Js9Bf0d3vVP0gDfmkSz
oRz4wTIGDONpntwCNmSHXPYCqSoTxOOIudhyyuxJDVvMSce2nQJHhQSjz/5pzaLlEAlEA/uNmpsh
Z6f+UEJtRR1EaGopQAiOq21FWHgmhcmtPwtrrZxGDuGhLY2zqnSnAhqO0y40jTC3JxqiUSHayK8G
82eF/+NPgcEJ/Fk+njO/Uh/SNv9/uisbXIa/3ibpp9udhFYSW1PLslitUrbjet0EkUxM43GPwhDs
fHmqe7O9k/01ZM18xjX3+SkBd1f5ae8MM8URZbxdN3vauBI7KfO8+SEdJHHCReBAGpdV9rFtlBOm
8SFy8C3w2gy0mK9LCavQqJxe/xKcRF7Qe1oQHaLuyw+ZTjLUkc5TMPhbOg8IUtBCp6/jr1etKRV+
w4yAGjc3vIYHp7p5aI/7CMeRRUbrqAIHpGAK5lRo3Xtu/F8wTmZglUmC3VuomCWGMvAGQBCbe/ki
JeabMZLgW+muXFNSd6jmcudFdN4Ny4woLWev33Zen7AyGshLBuvBLq958PTsi2+lSYZGT35yiSl0
Rcw6VcbEhV4dFK9HxGZCI704llpcCj3qaJRMuyqhmv+v++itdPt2y/TQUVUUV3QE/0fdkfiWChbw
N4/O95gDjCLy5H+cYtzNDiCcEWq36SpS3r4ShgCR99NDfCX4D8maXjDWlr3bEp8/x4qtBImagSNa
FSNVXc/sDQ6wQJy0jjxZFUH+r+XP0hQM34UpsKChv2yStEMZrsxt8wHUUVeglEssjFkTaGwuuhZN
n5gNy86dphXFIR8rVdPaAfDjcflml9qSIM7sxA9edEGg/KKFHpO5+TN0bhziplwNF1uTHuDpQhlz
eF1GauKED0AtdEQxX/IcYioliNy/MFq1nnXEtKCUkpNS9eqOpMMLvtTJpCceCzfM8W+P2M1Z7JPU
8wj4udiFbuMVfuF5PU+vr/NsfY8+h2u2ClntrbBx8nGEGudwifSDaUVtBnMx/vWTo4YL2ISspVGG
+BVAewP08871GbfzevNvaiOnHmS87gtzI7/9bNSpHvMj/P3aKJyfCfss3VAe7tk4hzKyhAUFRyyk
z7P7cbChaMhWo7UeIEayxlW1I+v1Lb5B4EYiOTilyyhfEhPBmqxSPTOQ/ysiJCB0vY7zOpvtOj+h
uRYKI7pRP7/4U0Y2RqpVaYSJDfzfo90Ly+UcYVVxAOJwcR2A2iQ226XmFeY4+QwfSiOwZX1CJBju
bvLyWFaQpuajTrbm/XMdcKG7HDMO02IrzJiM3TLlj7FHPG9I+n1YiAoa3p+Zn1kRHALPmVyLdRI4
c90kLUu/4KQHeqUQUTldghw+SzhYEvw5LAeEfxd6ztOLXTG7HGy4HNFotCtgaMHe81IYWD1Ywrl+
9eLM6+jwKcQiMsVHjCdi0eWaTOsY89H4VMbzUYJYEh8kUvwSzfbj4TQ1BELMoZoVKygWDEz+H6FP
wcICC3w6xTaHILNhlCFsbQduBC2nbzRYs+O4AvtCy2CwVMQCo7DNxH7UqCHKCw+oXyKjRxdaSjxc
hcW5UESYACzNcWoxBWVzrOK179zaN8Jna9jyA88VQ1mAfj+mCBT78Z9/+A4zNTS40XzKramk+/Jd
pcOjlnP9utc7/F9eae6pMsFln5Ug2Fkj89pAQr+D6L/5LvWQAur7vhUvI5o1Ej0Ay59dFeh7/McN
AAh0BQoxz9Uya/iqQ1GFNpCE9a2H1IcM82KnFVBaU9G3nlP5TYFbwpbmhSPq4y2ykCJDZWttkgSw
aCoVzVfpTBEm/2NForvrwiWh/UnpMaN6zWl8yMGsWEAj9WixNCXJUATsFqyAA9UZ6MRODiGkWGl4
KxOj4waSV6aelEEcojgkTWpJpusaXXx60qHhLRqxUwILMM99X499K4FWhEBFJDHDo8aVnyTb7Jv4
rbiB5ghJboBoz0jNRik5CVUFNy/wG9fn1mllehaUVOtXTIXv82uLWpLtvTGDsdqNkWyziR1yi0sG
73CUz30HuimzQoPfzeFnpVFUqFIphHbFU2j2JeaQHbpubj8v81tTULGUxpGVcZQVlx7k7DKEZ0O/
7NwZH4Ez3AvQKriQWh2AnNxXELap4wcf2rbM1nAWtBjm79ws2v5+ZQPCvdE0R8Qu/OWGYfS6dU4h
X9CjXqsojArNLgRvlVGn9kY3iEL7qBeArysepDYgg8Gx7jEvM3oP2WNCnnVToIdeix2cDLsh4IB2
yZ/zfDuTlI88Z0fl18c5gFHRqTPFmlQuRAO+kiMX/Gkho5IN/j9hH4VDs/n/i2j/krohkU6gPj/o
kNv1pQeVRh79gTzYFvfHwr3hFemS1VIFhnBaD5MiuxXJziHyzIRYOLYSzI3a8lmlyZgJbmv34Kvf
mHJ4B+x0wjFYH3SkMgwfVr9Ch+wdP9oQ/c27alSCzof91UaBuXSd9zir6htcxVEvY8iQFPpWeKCv
7XrPJZrGEJ+b2LR/l/jXwbInfsMV4GFUYXbqkKcJCpmxTi5HAkCV5J/2lDgbXILXYq6TreBIswTc
53sqrpZRtm0zMFFT9XicqNipmKzwuEejlBf5IfAQ3X7SYelN2IkIBAcV+vCLswg4oyPChOpruZT5
T6nHd8xi2012CLMRlIn/hx/KvWmvNazXIywohEjLCDuKugKPXIHR+Rz9wl0XH1FsFhh6biONWcjV
1H0LJQQ+OgcLJOA8FOubvrNKOmUQwCFbuqwJwVTMQSKhgn8lVN/j2B3xmbiJ7pNRhCyAsuTqii75
K2yOlGyvBRrh+/v+WT5UAkZOIn/EwgG5MJ86B3aO8IiY4oIORbf9pbO6WVa71NkiMJklvRvWU/oe
BaQfeUBjf5sQK0CJSj22HuTQNGc75as1mRKHZvuwVro5fFV+1/f7piJlw/3YNnOaYzKVD/qNHzMA
QJuWde+FMvUD+hEkHTcXw+3NS6pCrOo6aDU31njZZPbQCklJHRDziEaokYouvlXlkv0YLH/C2f3C
dMVtNmwWqhTG5Bw+DPBI96hhoDdNBHGNXleuDSRg/b0As64ArVpZYvhZnNwOS51wEgFzqXWUwyps
FoKI3NGJIWrM8bTV4kd1L/gQMOlBMFmGLjqZlFynSVkv5yk+3ysEP3JotVitstXrOy+94Nx/rrbL
/QCv+XEa63k3u1ll1unRtRfyE8oWeqxnxPM6Lo6xqMT9pGl5As3rGAx4Wf6Zp9K/mjraR+ZPim4D
urKSkdWIuGP8SUee4HfQazx0YMeO2GsSX1702jlcsSRLRCGYRxH+FvxbHhGpkgAm1GqdHMvcqBaw
8ZVdJILkwgcrXHf7PhZUyDMYWVhzSfhQsz123xJlgW2kexSkkA6g+E03AgnEqO1KAJqX1i8SuYqp
3J3huTJXQ8G/19HCSixCZTRJTYqmcVyHp2c2Ch9hpCXdbRprhS/Ng+j1oCsXIvbubY2BL6cBqTMu
nhZIpPFqnVl2fm7IMOQWNBKBiU9Vdstjmxz3ttKvwCDN2iSTz4Le7a/m9keGmJ6SdePYJkRbK7AD
IPehEWLXDFN1TRxY/MdzlAh8u+z9t8EcyycSNUIFZ8NoHPIZraRNgg+dUFRXwzThCIxrJhb56+ge
re4wO4Jl9m2rTEGKB83r2tOw+1shXtL/aUvjiG/Ju6hwDqXILFSHCgDZSBmp3/TjEu+RuOcpe7Gg
7tfwoMolC7F1xhv1CXwsMVWPyD83JagxDpsqE84SoG7HKZyHmOEkff9G9seyEc95+0Ouib7u78B9
7qI53OqtbOwNuzlhq9a598ZQuN4EeYARRfkhNd8jWw7uMQ30zsZ0DUmfnMQEH7w5Si1azYMrSRcy
Yj4K0+8EHR4zYq9W1HP0HcxBmR9x4oqi7r7eKClfholuyTSAwXTe69h5R7U5Z8+HJmn5yc225xrm
hfRvx9hnzdISPNu58Lh+3t3TTOCy9VUBoDXWvIe0Xzy0sRp/Ahyi4DNOauS+XCmCMvIhBe3qzViC
ubaYisVF/tjGZ3HHV5yGIpcxwKUnuLNQOH6hxNKfIPs0OphCSpiGxZad6k+Ch/SCX75envFHCS/T
kZsZsINXBDVnDdJ2lkxcRUcoiwi8WQzk4CvS6act4wQ+ZWOTQy0Gs4yq9D7ekoo9435Pwp0Ruxu7
BEWwxLNKfPj0PF2nfwH/wdmUMXdAS4pTlRBLYkK0TWjGBbspzU01VC72Vo+Sm0VWsUb1ZT8AwoSs
HR+Xkz/0huLK28n21ciRy/Qmg/VOmf06s7/HzmWaZJZ6SJ3WtH/lPF9LJrF8T1gRu37/1y8FZGr0
CJIWtlGAo9uvD60sBj8lrGM0e6AUQCvl+eeqfsdgwQcEu4X8hAyWl2j9tYpolZLvdu6xj/+fx8GL
7cC2MS1ec390FPl9iSX6n7x6rr3ds9C3tedRiQXIocAF4RU5R9uxj0iNHtokD41kkyW+3bGiu/LY
dlWVWcAE1ebkPt6vGty0HvmPmOC9tGwRgGFVtoei2YjnYGZUEt6ugVAYRcIHTGWyMuInxWDAf53l
Ivd97FE4eGCOCLFSjHkCCecCsx75Xzp5vTn4VgwFlx20nJlfQAx/2II986nH8FM0FTjNv5LuGvTk
EnvMr3TiZFu62dLvQtXE6yA6zuZCkNlILGkJ51X5hXAZ03mq/J3H2L2nfaokr0rKOmeB/i8Y41qp
NjqCdBbrjoD4djrxtdqkBx0LYqeF5Gha6A9v0DhLW4TOrNbNQBr2pNAlqlVy91bDiWpcePPBuwos
GgEVoSN9e9vg0KUZybCTve1ZMN0YszLmlKg6Lq5jKzO6APJ/QMnzjXaVoki/Nwr9RBs3k8TIuiKf
xFIU2H+vWnNESs6Dix6QLNx5QjjMgLOJAOM5HWrdgB5cEBo+ydX7WTWF1LXxD7nDViCip8B68hyo
0w0X6/pkAdzJQEYWZWLnd5DXXFI7hMrDVeq9jF2JJ2rpWEdoHQNL1B+kaRhEx1pVJ30s/0l6te9g
hP2eD/OXFWElKIqS86b3TtRPOdQRPLVyVN/Gh4K6/jbp5q5/Bmo1DkxntAEfKft/dwdCy2x5TN8J
XLodE1x8zxVrKHLcw1JzYB7sCCVQoW3Taz48pVIsvsA7VCT8ePwFFgytBvacdZjfY3Lr4pGUG+wT
Qc+O3x92vbgzGgr4VvhYcrnG2R0ImHPeQfZgPlQfCfa60CKw+690jGljpltDsREZ3Bzkjb9Gm5ty
EpcPTrvuzfJ08RCRRpyliBLTT1GCgBZ7i69MOxQ7gXPl/HRQCoV43iCjqsR1XYrUSqc+8dzTXaVw
EpHWstzJBFMKgkytA2zZn59/e8DzWEpUzKn02Rlx10y+5VGEQrQbUBHutRMBQvehKdPnaa1ADsxK
8gxa5TYBORMb+BMGo9/ogOMiBj5rLXUkGJ15GZYlinvJCvLXOEEKVupgmxrQ7yfAvLXS8gPXarqS
E7zdgTvbHyy60dYhCzcwypY+7YivsCut5FH81S2M1MyVBfCUnhSgw4wrd/Lbl73cbMcmr1T/02qm
Q6rAuzwMVrXaDLA8D3fhJsW2XLKAMTm6jYP8tozmTgJbnqO8PEFLD6m0ruuHAr7AMfp9a8HVTPdR
U4cV1tQQq9oo3ShOOpadtNYeqNj8z3yS7KFxeZPTDyzjikTcX3A3K/j+GBFTgOAUzb7f4cjoJ2zy
qTRYry53gBSi1zV9YXxPj81mLHRUcmkDkwq9++Qht9OmXXM644N3gOI76TftAiSPiprwlkcMRP3x
4TVUHFtteQhXtbmVuR9DirAWyaAkP5i5x9GimNfo+qtsFdpq4RbDLbSLgIJHzXrrq+Lhs1CBvqYy
AK2eSOmWrR4RfXH9tegkDYUsXBO7oZCSijIUTYS9s1MLyZIFZZ3/iEpey1SppWODDCIie9To2q+i
xq2hTS9qPxj1GWxOr1lOP89RGsIuFZyvQvK6yFjbvWBsb7NYCjE8zAy2KqCUy1uP1fsALjcjjkEe
vPPeRbkyVwSSaHFEulsioA7vYFh4uyDBsMuKNHuEViqt2zTCOz6bbkSvdca0hswEX6fvdL9An6Eg
N64SrsH/h213UQVrOyZoJtWtxiubkE3ZTIuO5kDfMF4+3BT1UtedkAf2BqZpwDdy60ocogyHHpRG
cZ3PsIy5I2O390QbzGSFj1/CLvCe4LoQZKd5Ly397bQs+ho8Qtk7hWP+qThCt3c2HNtBBVPd6D6V
HiqTsh7+VHk44CVOPI4T8DfWeSO0Yw/Kvq2XIEiBH2CsCbW1PcQPJHz3jXCkpAF4cBrT5cKu41AW
V2MrmxXFOWvwttoQWbtZ0MpMtqUb9rmLo5ErKEndmNUveul4FSr2mVbbqfLejVajDz0TMrBIwwPm
fc9pks/a8ByuNrACjk0A1v/o0c4VwRzPpCiLHN5csXtLEf/3DZApCgmXCADg1CADL5S6MoOlc4N5
070+mMr7TVXefi77fwm7WjnD4igvJXzyogCpbHfH46lk+/hf1HD5BKWfBIE4/8ks30481VHQXktK
p+jaCqhuAWEa5Duj1T/LBJhL2U6B7WoAX+jI8UNCPDmztndiFTGHu+9omRO67xOSiDnaNUcmEME/
kKYW/K19HCGEDC2GU0aUsFsb7j8nh1pjQvjHeRwz6qXywtvTF5TgiovWkdT/Q32vaTPIn+OPpZda
J/xv+UrDc9uUXOP6pAmCRxayIYHp23MHck0qLuBa6ly1wqEU4x0h9Zis3LZ+Z7VCPgMFIMtVqkgb
YlGG837dbWhPGL5VIjwpoTM0s4l+LUzEtQXOfJ7DGnRVyU+hMV1+KAAq0BGGlKC5bSc4VMTQMTkz
T4ZMko9DxII+bFDy6tOvDwjj5jop3ArbZB1cRdiICJSkPWEI+Q1pD6wXthzV7qA19A/4IR74FprM
WvbjaWAitMG1g6ErT6z98/EIrtCJW1kjWfj3qCdRMOhokN1UqoxpS/5eiZM2MkZ1QORh6+Gubnl2
tQn7ttMQHl/4dJ/Auw0DekKE1PSwSwWFVD6AxnikARymDCofz1rXT58Ea6wjbmLI+SLAZzpWkrEX
tBFddWEo5UU9PYicg7Pl0wZauCgclR+0Yjss0CtNLEg3gEJ+MbQKdW5ePXb7ig1u0YAJ48xHqqKy
rtjsw4/F/oZ6jqsf/2X7Z6zyoxtCrndIuES2OqK8LBgVdO8BqWhppX9SQR5wx/IdUWLMJGrjCYvk
n0bkO5I4BWPA7943J2yzcFnX5rBu3wLlqTKJfm/ZG1odirsmgrWgksFzMLEvOzxcHr4Z1A4KLjZp
47rpjkhtggUXxZEcxSvPLDtUl7KzH0ayQfuQqX5OIgIFLjTu/RWdx2/lqsDFn/Sw2ZE3WU4puA1G
sK8X1XysqjHR+67MoLfoCKAtG65ALekdmW8IvJCSuBsHuNrMq+r0hE3Jvqzwn+0UB0Qzb67SQvwL
D6xK9998WyhGMjpYYF1hhxI01aQy/d5dbsRh+I0HSGWAei0kmr64Qf8FduT7LZ4Ym2u/Bobv9zkj
4Cn3YO51SxciBZbi7gDEHoD4y1QiYBwDFsag/3o0Z3DVVP5gMY+fnB3yCQ2A2odotYZHB2fyXDpW
5CpccE3YN+ZpByqXwY3tnStWnPgl0YY0pDxU1O9/wlVwMGxi+Ck+OF3lgmlDMnX3xwnobmAqCECv
uNkMYFqcmiJVDwmI5/k/PSSHd4pw51JCrrMdke6pf0DFAIMwvhKnLwFLiQPWl7mVzpBP2GAG6rYP
Yd/xjMFKzNRumxOR7QkYw2T1+8D6OyaVSNdOXS70Cuow9fu4KkMY/SBvkADEzGHwEMT9itTPQ41x
ZM/k4XWOT6iMXKis2s/GVnuakvmlB13vU3PceaoujWaIokN2QY5J0Vx2Dsgi+ToTSqv3AOQTuLnH
MXzI5pOCtNesDMpK+7q89nhTKhc+OKuzdsTsAtWg+9e/ff68zo/OcIUpRMSngoUm2C4zPLCCWP87
mu3DsJDwfw1S6KdweCW+DFDwJ0xHn26k7hBCG/Ayk/M2nR+5bObJ2LJ3Octo1A9sMPGGYqj4X8iI
PIorlYPTmlTh6QnMwy/0QzmcQypfG1YEOWdrtmVLaXjudS1wYnV9nccnXgeoVLrIc59JGuJaZyyg
Y5LHAq1SFpUcPQf0RiCu6fvjabBvd8l8MDpMflEH+CQwnB9wmGBzJlXOyXwWmH6nSfBWGBZiWRtQ
bm7+kJmmxsnWEAM4j6cm7+B3Sx7dIYc/srdTKfoh7f4hMChorYRZh76gGxp2W1xJBFTKcYCS/LNB
DzDKXr5ApKzRPX+FRcQiomP07kBeGTfJA3O536zcQec3OunNkQT3tA/ZK+H6YUmIQH0ZXdRqSRFO
knotJaFgNgiisGpd4lmHKlcHaTKOgVmgY4cabIpi4Lsc9H9p5gJVKr/qo49ICNtt5/snIFoNW+qm
epA3umuiKFnAg2WC1LuMfaiA0jTfCfK4MF+4wQHBAZ9PMNlyKkfbkwAO24oiSTvKPa+9sp+t3rRP
vSazU13Ogc+8kl476JPm7zsyCBLcoJhGaU9s037aahkd7bYH7eTEs0Bydwn7i5sRxOZH4Dtn5Z7n
dJYx+ou8jwyciW2GOWVjUiwHxteFQp2jWYi12TYzV4hLcjSM/HOPgd0vXSdFt/tUswe4W6ccM6Oe
O4d0+EoVMUoOyEPNGLfNHkDJ0WAWvBr0V/3bTOZz1DcQRNh4N/BPCCnz9CslLwE1oAu4yFyXHpOn
POHkyaVOBayqSqUYGox1MJTbC3Svz3wmNqLjEwvQg7reS7oRr2fjI/SSAmigp3mrVz9xaayqbV7L
GEIhwic2MA8QSx72X7i+iIT9qmbF3h9ZAeC3JQCqSpb3I2i4gNJ13FsHwtVFWkI2WnfLAjI4lsa7
CgFXYFLil1rjOaC77v9jgqWKYDbu+Ewpx8EgmOBWBrFvcEGWsE5Np0m7py6S8Mdef4rRLycLsf7q
ofvvH6a5IOwYz8am0eXk3PgbC4FSospiFglIiSLiHrf1hcbxt2nohb5vlQXFonsONAYhTtzPGTt1
ZKAQxcd4Pq58cQgM1jE+P9xi0+HMdsMCAe8Oert3mkCB9PDYEHQN3nYB/ZupPD9ZIYDwaNH4D0cp
3GmG4crP7Ea3cJv0kbkWRsID115fhVnWCPvYZLZ2y9mKlSCKY0ro/+27pN3gxcpQLxUOvIhr6ZVT
jhMLNY1rWF/NJTy/3F4dcLVEUXu+fxFp1IjqEznNQBkq+qMYbKsdqt9zk5JGKqcvukywSfMvUWrt
KbSbwsFvTd8T4SR3S7HYZ6hcqw7LBJswRPwzt+fuicdJ7ETRc8zvOb8NlI3O7kUKQQQ9PhpsL/5K
fXBpKsmqj77Z2ZzrtMeX5/LxbTktQG53HZZZRB1lxbFHgYkX2eb/kDOoMbgE2y9xp2dhkifrtPNA
ThH3Tl3UZGudsApXDmXjJDKFIkUiT6wINEhMEb5IIkx/nb0C4yu9QrLkU5GSW445/sDd5PoeAY6d
a3HRLPEW/GNKzkEr55W9L5nrm8FHot0S4FujrLuaWcIHGP1vgOAZPFJYXaw0tla8EUvCn7/wDZvL
mbiAuNT6he+NcqWoHEpj7xOzfzgr+JY6tyI5b8ul2fUX9l+7ODcQ9mQCzbIHh9Ncr6t9VSHsUP4e
XY3NgNdB+uNWg+vnwce0UnCYLZ1lDDBB/vajXo8hNleH2gm0j6ZMTwiMyZo/s777lovTS5vuBTn7
nAPKlw3ihKET+uEv4d01vtWntgNc1ORXHRm8yW42TrsU/dJHUU+gvMZrz+nB4uC81j6reBdkiepX
o1fyrGPWTrpXDX4+1eAfM9EkY9h1pAmql2swofvBPK61VIJtx+L/AiCPku2M5kkqnpy/7sueQFdt
Gm9Yu39IkIzCR9ZpSLyiABB7ONKAeX+dKH2cOopzBv2p4ve8zDr+zvolGZccnmncuSevVnuK//yL
uBug3HlL4rPML0Xfy7Xll6V/l2mqa6Xrne3Sc1B71WB91M/PjNZ78l9OtgU2WDjSd7PhMHSixuDY
+Y3vyJrxnVQbt6ryumS3AWpfKdaO8jdMVXmCaYvCl5lcwXO2ZZxWcibc9SS/PL5Nb+nLX8AEPfcr
kud+7jQttjiedl5FYebFD0422MELTjPZHoI9zohzOL+6nA4VTPpL4c+76XQM3d23DCIVuRnqMz8E
5uYvlnItbJRnTboDejz1wIUemgdiVuFtJqHWx4Cizo0ZtaXjMnNpMhZGQJbkLDzMIqSGzmkhJvuL
DlLWplbdLj2fUAd4mESRWIuWWw2Ta5WDyUmkxmkHkwcRfDE0cDuKDhzSvqjvfQ8opIBc8J8cvViN
naG5HFXm6RupTg1ur6Bc6W8M/IQn2p4aTvLY+KOjdLOEa0i5upQhYHagPhS6urfffjEbHZDgeCaH
PIVFe4bljCNVUSRQeznyKHrTNKq7UNWtnNTqsT7aU94Ei6bfc9Ez79fe7p0q1lpo+6KCoG+feT6I
91q5rzrLdI27QM/p4sIm7/cn3nFTlEzNtEfw+DPbYiOqGfQAgkETZalItAT6yFMwBi0GMtU30lea
JAY2GC4klxx3xgxPme8hTzmJreOemJF9KHt/lgcju/DK9yuGyTYQbA/2lMfffnouFZDRpxYnC9+u
aI2iVzpUgUv5/k7ZXGveMgWjjzyS/ZfAACAo9JPEuRnELsHNRwp3WBVBATYkjMcf15jIA7Z+gnsc
tlsNJwlI6CtwG1ZDGqYb69pr/R8hxms9Z0bnUtMYMWf4AibWP4/aMneaDZM/NWW94BFjTmY0FAJQ
VoNGZxnKT1feLmue6Lk0PYVqByec9V3pjEfUdZaZV+9sq5e9D/BJJljck3s1p5IWVwO3DxuJW9ot
JUKM3HDK64uNDELYDAc9wgd8kF4wAmrrL+sd4MH+/v0yYYmkdFsa3p1ZkSdv22fx1K4orp3XquTR
Gxzks2PbFmNwBY6OQTkuUiRqbZe373DXndYvwn5N49M4AZ6hKO/MuIUOYfz+irYqI+ijdVjs/3Oc
6sSZOBgMO1uxmyzrb/kBADoVV79R/1fAvjXctQEX1UdY/a3H06HgBo0+NgvtdgsUpg8gSnRIbd1d
tWEzu5ydOCRgDHYSdHC89ZLuqZ2pU5U0RKbdafUXjbk9b41OWB+bToyYNgnt2SNLVhRYg4YW4uRD
LmVyZnw32XnRM11i+b1tuC2Ggj6iEnA5ciom6wTzLy8qk38my1YV7gxxeOEG05hzjMyy9JzI6tZL
1exLZgSqVemXEqn+sORG5Oduxavu+gmhPitzgx3ZBt3+SGj2OjDq0dwLLJ+J3YR/b17QZj2SBdEp
y576F5E4I+cCoATd71xZqLJqIsRYt+ojyxgHUO97QeAMY0q02BafwXHZ0kmXJxKwxazBagxSghML
I7Rx6vXXZwjNXHT2IVKgpIA2VOdgACeAv7JTUUfaCf6RpAI3yGSc1lC/xINm4vH0/NmaJ1m2ErA4
hSX9Lun+NrE6vJwuuEy+Nyc/68bExpYUvrECtRX2SoYbAkmIx2abw+np0fn6uHVELWE51TNBdaMJ
b/Ra9QMmhuk65nxIWrfNB6UvlXZgY8zxTbv9CgMAlziPQjMkTE1mDmd6CkMSCR7Ex+dryRPT/3GA
5sUSdSqchRNjrh8maYTRBkWIqquzKlVB5n/ZDs0qezuliTlrS4n8AWALwPiDTfDCtC5kBnxB+txL
UTuX/SikxnsFyIrmGqKln8SsZy2gaaO0RAY+UbROUi3MHdbeq3fYjPVImUIwLAxqB1kOxpGaCxVe
jdnQ45pWjvS7JFkz0FtRyZHv71nBgVvTSFYCUyB1FFN1j3BCMtmjhQtg/bTs9UNENtsx7HIfW33L
mbM/X5DJc/IEi+cblEKnyaIRgfAfc6Y1YOWB/F3NOz0GV/1LkNe1QH0YBPrNztP4IOE4nbz1B2w6
pzTGyPqsLv/6pddWl4dnmGjOe7QFOX8udwo4Ri1PKiM47JSwf7OHIzZrfWjen6m3/UZtG54pIMuj
AVVuZi6CrEyVjSizw2doNVe4EIVWvsV50L7zsdleQ1kCbMF8heIfipCVB0vbfl4i9oxKOhjGmPhP
HluRA0iucMi/RdPcRM/RiEFUCg1UlciGXTQLGqq3lU0aA2ZXY2Bzsod+MWRdxdrvdjoI0vMyQiOY
oRo8NoC9ID9TmdwR3yoW9eW+UsB58h2c5X2W1Ky0v7Yw34KW5URIfXoDFaZthXwJMfvgrDrxlSmW
DA6AENhdqL0Q2rpyqMTB1MoB9gvJsksKh7CGX8Qlm9C7hgRYbmuF23rSzqjcSzXfm6klCRtxSuv9
nr3PiLxqp+CN1asTjAnQxFL3uZ/Y7yG037GMr42EYMdBkPZy3VKkr/ny3CS04BrygjYyiu63E7Od
xRz143bNI0gbQiiVkbbHrWjXIG7LepUzKfb5ZuEyliVYmv8OJD+0dOvsyPDYiG+EUehNV9MW10eO
WX6rlBX+Bx7o3x9WA0oDZaV2l5H2OKe5TswLeg+QF1ZaNbX5gaK2sWFwt+LJXu8GqbaWk8x1BTmS
Cj1klCVH6Wze6HQ373tEVIhpVrGgPbDOPP1DZoyXkHSFLLJi8pMvzfhU3UX+L7Euh7MgnvLHvW6z
yTBhifGytumojKC2ETTduWrLSkayutN7sPRip0eG0TI0s+CKt1iRCo7tJMXfYoSC48VsSsKqK3l+
3Ys2asH2r0xTlRiJDhg3PpDAEvUr0+86CCaymX2JfyYcG6O8i3muTmA3KtxBDl7CQP0WRkMajhtJ
ZKjmja2wYexb6aWc967HIdx6cbYWULWjgKRTwKW5XnvNhxxAZp2Ui+ukD/ubtvMshOcCO3js2+pW
9IYO4awvifj1gRo7g6azFCSscqceIYEUHbVLFGjN3AzCrpXw4+eRe+EMhpbj5m88D99sCEw2ZN57
fC3U6lDGKcAdHUxXjPOjnTL6y4+VAWKhHufQU7XJlk1b7d1iPjOe1Jn6AlVLBgWIZGbzJ7ZP6e0d
nZ9BwxmJkDKV8tOxQliMqdcSl0ufRs8KVjGZM49KgiVfDjANa+ke4LSvOja1l5wAIBOYJ3LGl9hS
ux1ifDgdyPwIP62yLO2UiHESjHPOLlyOeelW9in3jb86CmEc82JJAelGShqWJVvmhbaPyDSWP1lR
TMW6DMJyaOpuaVqx+iiQqUUNbKtDWhlT0CRtiBmfX3TcBblxzKhrp0MlBB72Cf+5MYCmPPD3qamG
42w1UbswMuY2yvGK0zdBL7pXPJ5bmiKav8TAPsGFPgjy+QQQUSjJ1e7Xg9I0//VD4efB2ZXNaXX6
ll/m4BTZQKiiuvUBntXU+DBIAhzfHFZNb1rCMiW7M2kJ16w+Jlu3TaBoKSG0tQtvIqqP8R3Id5aQ
hpFCJqHYYo+8R8mglQsEheT+PSk+huiTOiZ6z3/YGqpeGjQfuMImJgfgZtwrk9ecosIrKodiSAgK
q2a9OIM7DyNVSYoXDYdBJA6oDYI0UhXAz96RO5ljLglnvObsqjYVply3lYW+t099KTab3BTCjHgc
T53DelNaHTEtwNpI/zWKNK7309K3jmCAx5NX4P96Z2sRYD4dKYiXUy18kQbMFs2z/QvuGOJICEb8
4DTJgLxqx6hV25byjfHH94W4SePCup2YfwpYADrilv+WYWCUA4n/LnD7Vt2Kpmi9vwUcV8AcFBgq
o1sv+5pLPt2u9aoDoBOVx5R9KlhAUxqoarip/ELwI6/anEv29uF08eiFypQ774KaODPyNO+SA36R
YXcJkBxNHVWqNBn8A4yKCA+bhF2Fa+4Ff7YlYJT3htk+J3bEpR20+8aY+ldPTiHYiimiRqFAC/3a
ek3uzMbYxKOR803gc8x4m5HrgdBSpgF6RLFUtSCUQkia7zF382l/yo+JvvAedg4IIeu/aqFOYRYQ
B52dN8hdKapP2Qwx/EdrKHAOB8UfWQRbl6HQbY5ROfLwqtrJ3RtmEQidBxJTSB7+zDHksdAPaWPg
Rx9UgeWfWWhJFr9ZQYEFwVxCMwdDDxlhJunedq1ox+TDfP2AdNfkkY3CxFY8Ke3zYQqY5WrCavVg
4zmal6no0FpCQXwTRrG5eOs8JTmdFsA/cEJrBvlS2A4GPhW72aSG0m37ZKfCwj7B/YpY9MJ0U4Jp
lBo+zLBC1yirDR54RQLrwQ6vh50c/T+FSuwGw2bJqxA0oIp8lofkLYfyn0EED+vNvdkuHIuo9GrJ
XucD7zgDiK4nvn8LGtw3s4et6gVZmiQrmKcH+8LzXKg0BHbHHK5fW2LQ1t5wKrnKvN3m1OEN+YmD
EuhT+MC0GFhCDFcj98y3qwwRgJVP00cfmaWoUaWh3Yu5tPP0ByrlXiIvJSDcU1V+fNHrZGJACDlL
f10BB3HzFjis1btvVShQu6OpTuxbsawxF9epvWj/w+1gbDUssNO16/yHtQ6Dq4tWZZtX1fKAPYPI
eNyaS71rRxwC7JMjVZhEFagcVSIpPJP1OQpxIWnc+grz1rzl+aivVGnESD6ietO3OdljOFS+CZvj
SxVIg0Xn8bJEpYoc2z9yxHD3DNRPvf6rN8WO2do0VugDOeYoA0CuxScCi0WoxFqrZZr42mKdbAg+
PhGoc86GgQhbLaSp5vVo8wZtAvxHpnT2Kl/FXBuUlbERExQhQJwEFxElnwaR9hAHqQBu8rW4OgY9
0BGyPCxFxX0/yv7bAZm5nMsHWE/52EFYf9ms/xn2F7k+jejSdnINvh+FXoXUTRPlo79O8iOP9Xgw
/BA/5dyIpKrLD3U2JvZHjCREVTucAPSU/2QTO6nj2B6x2/+g1UFqbWN/NJ5fuAT9Vs9zezPEEUGw
ZoRRAs5CcssrlPr6gFBdPkOYN8TbOwz1PAm/krs6tCmRJ/E8YuBDakHCw9/5Q/FwJx9XC9jwLxT2
WqhcmFNAn/qBiIH+/Jl90YgGLpNI7kKlyVGxfwT3MaNEpX6grFoOxVtLPsxPeeM2nSr7CP/kba+T
ZzQcMPNgRuC/3G7cOGEd7tQ4N/lxxff0/7PBcGVmeNdJrgp9WM+angGekSNvjkoq4yeHUOlOdX7o
e2mspOZnClCrSMLey8wz8IZDkB4f6B497pqh00imdbAUQysIrg3WUkgj7PkQEzz+hnODseAZ6emZ
xch6XLtWy7PeNqVdpUTwpL3tgB3PGvMMqhSj8EobBWc+mXlmO3baQpkty4H3SrEtACNTE7RA8YRS
iQFYCcGlFo+dNNaJ/bMcNhq9jZ41E3v3pLEQKK8DbXio9lp/T8BlSNvtlPnwDV0K1i7Iim0wh25q
ydup9bprLU1QJRloIuTJjwLnBUG+mlhXOyoIQ9hBDupOjPNd28caY0wSC3C3/+OK/CyoUcSkWOof
QOCyVUTwkSVvs1d99Q9X+p9cve8V+luz1zXoWtDlrhC/ToSfYtE+jEmakBbXxyTzpV0pRVCQx3/Y
e+eiAqA5AnqC+fX60quJ6sb1SILl8G69QFcNLCMCHqQGJfR2tR/dVJt8X+r/qIDNWa0HR0ECG5Kb
19UxuKpulQc0di4YEW6QdoKqnWAdQmS3TH5itqxnRVh0QVbG9wIApIYuw8LgN7DVelFGGu02WwZg
KzwtEijO0U2yMbSDXeAozc8GAb7pnX/3S6kQwOOsTY0QK6LDOnNaRaeR45Z1yCWAdNqX7Y6lJRRH
WS2Vw3OwQh6Wqyk8r/7u2AyGNmV+oWV0OgmGuI/8WYj0+Myb3n9HRuOxKhmQncnD/7eodaEd4vj0
A/puygGWyecBmmFFxqTyu7XBmxd3c4R34n5gFYmkAw3WMBG0sIh9+EZ2wNkjMg+xe9u95Eaj67s6
GY1PdxvPxHfk4pFfbuYamPLXTG3RCoAEK2YrmOh1pNI28th2Ku8PTE9w6Ry3POMlPulZnrdG24dx
RMbW3Kt0Hk5zI7IRQwGGbUD2jWetcsAx5zXI6K8LrihTtkgohea/P5a/lo9PlFfZ0vVcOz3M+VhT
0jfjxN9CG6UuZl9nwNwGpvWyMK5LZrOi3CX5X/zBITZei+eV1OnDHUtfh6SmvM2+90669O1H408K
nSscX0d05T9TBkiuy6AJeJ/IG2T+g4oRqBGZmqB5lIeDyzOEfUV41hW0afBwbwC9ZcpPYavaY8ow
v0EUimFieVmnd3W9iNiIdLpOExjlS8ev4SKeJ/Ev3SjsZzX1UaBYspo73IMaSnXISNUu6dg2aUEl
GPvfV5QiYAxGjdEEveGqn9+gG4S2GAliv3pHCOW4m0MpOx9HE9rCYwTVjpdQ+l0ROSbMGjS+9HL/
yr7l+Nwl4l9Lu/Sk2oWUv4q++sdMWvpe9U+6P4THNhRM6WjD/qdlR0nAGyDeBpa0gm7D2lMGILQU
i6r3vs7jpR1sDPJ0+grFHCSzcO/fqFH2eQgIKT2+WOFkFOrQxgTpPWqUXfepD3q8P6Bx5cLV4hW+
AFDm6LDYmbxlKgmbNoHupemihh8NnHcD2uiRnzR90PPdR70rQvsIN8ErlgrE1Q6Ys7eFKopzNPt9
YVteS/5nm+5qWmQ2d/Vx7KFmSC7wztwOYB2SJyNjxZq9vLwodtJScb78o3hB3VjOS5/Ga/UDbto6
gId/C4uracZj7pLg9vWQVBo8+DjhzPBY0i5DNOAwWvihZ3iNJGD2QCySrL7F0Y7HfYjBbFSFORtW
19Fc8bcNSin44RMnj453GCnubWijr3f37wdS1CIq9KjJscJGGRHQvDrZoy7KpgBEbhITsyHauFeP
CexwdHItXZTtJhxG3axR9+FRVaSpI1KvlGyqDOboyB1i9ax2kMGaDyYOUmXTM+T49KSTjDugnxGo
p3OmeRNCjrZkGCk49qhmGakD7aLIcVaZY4XcJTC5d0mC/zcLR+kxhPTLLzZYptfUn4Rz/TegsycP
/AO/6L5eu4eNYQaUboGupYq3+l9jkAALPgYpg6H7ac5Qelh7EBYZf8zEasIbQ2GcssPhhKVIiAqi
K9PykmDEileUzpoRgnNcqCUg6MMFG6qAFmaym/5/6nrvOQI/PrFh3CH7yM46F4s8K+AVT2yUWeBR
WG7Z2MCiSdYSxJQov7GlUKpvlW5dluxMOG0ZkMWXI875T3hTrBZ3ZBkZkDCTt/n956cgyUJbQZE4
/Xp/sHBSYPDU6CT6igLisSbehghFk/+4E/M7HpVlE8ECGnJnUCRKBVmfT3xT1+AR5FbguDhSGCvq
NsfhxvLgpAPRHUQGoUoSIheE9UU29rz52DhOvoqgOnel7Siez7B6fNNjaOid4rkcJVWPX5ih8H3x
FaddFfL49hu2IXAV8zIfuPx5iLWDjIDONXNJJmotMY9EgXg4OohVnwDygORXu1+kIgJsbc9T6/H4
xNnWD8UobALXFhSK3GwjS7yGalo4zmUlLcR3r1/yCbQDk0EcNNHqdNzeZQx6dyn3xuuov8ytPnfw
dectMESQKpELulfb36rMo0KmKdrFRya/8//6S8Q4yyhzzmNyvT2Wtyyn7gY0CauGmlxfVAY2aa4d
NgGZWZiX67gVXU2Rc8KZDHe5uRTXyAPceA9tM3huo0srhB6Mt9jJr/09AEnUMn+7NtYF3FlGmr2p
5Ji39s8wZ2oC23e7GDxy6Ez4dKenqPzwyppcKZFMChQ6MgLx51Gnb7+QogXpKqs14GaULHAP6bGX
fXUdqPvqIpRqSgC7yhnriKPWt1R6V2Dm3NQMgcbwQbY6ud8kAzjWOGvMzqFvDcbUT3Begob+PCs1
XfLeAbw1+MAv4AOlPxwbDx61ZBdTwx/eqT7fAhhoLWMcTo4uMDe31CpRj/bNMjylErfnAJ/yyGaI
y5x6Ajju9Oet8nj+b7kKGuICxf5qxQ00Dt34pEqvdkzA8nPx7EZeDNfRpU0u/yknb+4GSxJegMiF
dzzCtrrCZMAaoxknvuWpZjp1w9SABWex92k8eSyNLfKKcLzO6x0JdFhzC1hegjvq7hQ9+mA4aAkm
ukePNKSkvFhL8c3/hGGXUhHKa7XXEda6fRpknV3gVsg3e7mkX3brOt38uhutfKore6uK7IkN9WP2
L+zc3W2zgYg9gG6ojOtA7WkV2e9zYqp2vqCnAMKupQ+z1uBV9gGlZxk/HA3aTmi80D7W4HEdv7Lw
ezFF+HwnZJ4zYHkAVXr8Pr6gOJi1evwr2ZN7hSj8qGUP3iyRq7uMV4YTeS3VwqV6dgY86YhvZnRY
eYFCu/qo3KX8lyS+Xt2WAWxUk8KCVvkv6zdPRI7K3So2EBBealM/D3P5KpXPXbJr56HtMKvSfc8I
SvjCZPCh31sX7F0LHIE9E2VF8h/N97FVpcVI2Z09zlFF6BdXPIh5Pl9ZoPXjFp9mAxLvjYSLS/Uu
qDUPopbGzVjvFppBinB7XIQX8Fde7v0imrQwOzbHWEptQGR6YNnQixewfhS/yDsS5vN5hGj1vKjK
xtSKwa7Re+YT234+OZdHggsEGbPbRhczc6gYA+n51m/X+7xmiH1uvidIjO5LvrXLrd4qEIU6rfkw
PDLdsNaUk8KAAokjkfLWuzY/j518mqb0MPKMxqFgkuV8YqoFLxFCaOzn+2o84rixn6y3DVdKfuHK
+LLzsALiOuSLLJnv3X0LzD0FmjSgXs3yhWG/2CS909246sWwFlkS+5jvB5G9AQx2USCbSk7tLJwJ
j9ufhnVXvKWCrgXBkpFGV+/XbdTqcZYi1bu5SANmbN/ObD9QZ34ZTufM2ugrtVvvZXZvNZNK7nxK
+SdcT5cghK4SaI7YwwQ/EcAGKHo7UWn7BhCTqt38JfVfzTCuVWHBftdQTtqlZUKTjUG8bfgmXsJz
JxdpZzEue/PTussn+TTtLz23ahSBDIg/JiVW0Tp94RnryyDv/QW2Q2bicaLhRTB5/DOSgTzBwduK
y5b2jCLyorOm7xFQlz6SQZaXntJfwm1n096tOV64E3iGjvgHR40yN39IIeYnW5gCmnnJg93VYUs0
RW/s/OWndaVhFS2u7hrsPJtGrzyBns/RJPl9LQ09gbetdCedaKVcy3xdrt+VLy3gfbFstAKShh66
sEDR3+K1YPLpPfVY/bIFa7h2svbCttT4WABRY0aBXbqxZI68AVj2ECprbCe5uZGPHkMgqCG3ZHC9
GdvvRBPrW4h+DYId/YSAMZFYBgPyYP0qyAnNgXuxkk6cWrl2BPZp8O0+XKNV8IxyNfP4EJc9cAt5
VDK2awMgNXvFVN/04sYA7pfHx4EquJgHuLniP92J1zgFcuKGF8l9XHCVPhHfv/MocWYoOkz5LzqT
gTE+hGIct9qSYfYt0J76edlAcvzLJHW4eBhCIoHOKaFwRafKVwcMGc1r31Ty7C1FgxJxEcx4+AXi
QG1asx4vv9f2xT5EfpzqfxbPt62VJ86UGELsoIBaHfvHB7pcJmGjKRZmbp9d2E6qW95YaIH74I17
3MGXVOIeY4FvLEDNuhpuybuNogPwSig7rDmUMOhSqRzd9VK5tnrghIMnHsDbLTQ7JYiU7eF5RfVH
5bDfwblZvT+lt8TuZexub4TO8g68+s1ZwXhJHakCZP88lCpXoF359Yzhv+rmHdLSwyMBqtdnN1E+
VbpEis5zootVVQLD+ds4htXQupLLaNFWS2oexG1Drd+7dyJY2BGFKGzZ2jmqauKBWVpFdextip/k
RJ/mPX6mTB+xgxoyoelzrDVSvZB4VPBQeOlGMsw1NQ6+VakvbVegz075dmHKT2WgcXQkpWcM/lRZ
X8ODw+JecPJC2zej6ygF1Kxt0AFRt3OTm+I1Cg+WjBa1MQiqCnQ59+Ma+udU4z63cu+RR/+Iwxnh
iZbggg7LSs7bvtB8EHDiUGYvlymivXw0OZ/RE/kBvYIWa1lJbee8i2NPOPwDmwju9lpDTA4vsYnH
Qx4bpt5FYUXoPJ+DQSPlVwraxN5nLi11Z0m6cL3qqxESwXGfR/AyQ8byOCMvALAm3OIEnuWBL97m
xwHjllKv+UpQETexuOHeuGSQQFSAcTB7xGeSTeNGVVCCjgNPzVl5w/PMKBsVxAhqhazIMvlKwUFk
bDpCdHZb4MDfkKB0SFFR0XJs57lvlrCRjhYfoLQ3g9G/0vBPLckUQQbK7+0FvyOzb10aBiK0S54E
+qjYC8eLsBvJ+shHPfCml6c4DmOB+DdS/iA2MVgKS+OBBY4fURIRDQQYe1bNo3tKX1AMQxthLNVH
KsSaq0LrlI3NSL0zEsmtNR2mFiob7b/tdrEmLX5AX2oa0MKODzio9utpazGuey8B1V+kiIURKlHX
aGrsFH8LoEor6D5pJk3LN1BbNM/w3qhSUtOkb7lZf5g8cNGgAbGl3foYFe1eoVQAtblPsmpzgBZa
2xch+jLI/DMnQIARZSvqNtrdLYrs9BUnldb3Opv/CTrbWhOqph7oSFrb6j72AXYFq+nbnyx3gWYB
5ATVfPpZFmD+jfkNOlMs4smTEQdyYNOOMsaeeZ76DCaQI4iUmBYq9XsnbH/tEUf6gxt2+Ca2S4R4
mDQTr2DthDUsAn2WWZzwHTfFcnqfu23cl0IWGYl7u0wF3l9mrtTPbktvzXRrpyDtsRhxW63qVr4Z
SQQseBxnOdOhnzaFgsCggsLKB00xD7q1es4djPwNFDHP+yGjfJZgvlI7hghFTFgx2c3xpVHHqqHW
/EYqd9jeEylLBYkC+QcMGU2jbD7vYs0NF0XhB7OkC46Apn4+ilfJ4Vi/N24VM+HE+LtsS8mfw87D
GFdTsVARZP30BHui54rUCB8eggFMOG1QEkIysolpcUvPHYtA/fFIf/FYetlkcwFDtUWmHC9RPZXs
7oCTL8NJ8XkJTpHgNTnf9u6EqnTmi1n4tM+CxpzMMBb2XOohhDGCVJUAiV+pe2tXq7xv+2FojNmk
0DkooqH/zP36pMhtQvZ1bOPC+Glc+bQu1U+wYFBtej5HAoMqQ1tQ8+5ywF6aTcMuuyH+NgQxNx12
PBDF3B99r+tV7JWIbDqDVHrBEPMdMHZU/ZXYWzHxvZ4n2J++ViK66cuV90My2BJM11UwSHUzSayE
WEbRZdLsh97gcPYo5FMRxWHgLnYP5Y6SULaJUqEA7/HuY9rvVWgZe/4mt9Z1DtO2acNefvoHxamF
iR9Jz9uVukBfZZX6Ke4cicOeH9FzjFg0kyT60S0S67kZ1D+/Ne4A4qb61KaSr3j159oKKxAB1t2k
bxxA4kBlpRXcm4eBAvuQguLqvbIykC7rqUBJss/kvuzVW0tMzPiZHoKOUXItjTORQjl5/OyAjrBi
DY6n0kmsDqV5+OiWiQQ01nUIPlGMzu7c3MyjGOzE0WypP28r7t81OwXz0vHZNXlgd55z3OpItbuD
Eu8AkP1WXYE3Ceh7RRsnFiYT5mLPZ31mzYtEacIluSosblwpiDNkQuBl32cqiQSNRk9EC0EIYUxb
xdBazj6JRmv1Dh504NXSZVdF4H0o+e2eEKQ6SA0UAyrzX1ETx0K+tfL5f9OUFuuQ1/g5J3Z2ZnLk
Y16WGtb92EnelJ4jS0BDIxzsj0AgQUaXvLYzHXSKR7ZmrdoE7n4uImt/hZFJuw+2IFuYkpj9UAH1
SkmCJtSJFg7hg5vOV/S/hRZsBpUP8z8M+2N8N9A1rQErHBvyvKrOW+52GtH7GJgBcMBplRsMckSv
eHz/AumUbnchAL9owfxKt18edwyWFMeK0JFSVuLU/h3WXu2Z/XO3NuDBb0koKfGWQO617GhcP1t3
I8yAKpqOU0maMdbKGzj6lDJAbdOlSMcn82eP+LAOsugEkHy2BBqO9If6Mwtx4ZaFAINEuUD66HxC
C2YqPGvMFxXf+xS77/p/UHXOzEoCQxj5bwYY3y6EQWERRYJ7sU2/nTC9tYq59mfNckHe/5Raerx4
zvimT2wtm9eVJalt7BgCPMRC2wIcUhzUJyS6kXrxsHMqgmie6KmBV/8HTm6mPz/JUcGaVqi6BVbR
6Cvh3x4YM0Zlr0IYkfqdVW+NS3abe468tgiSGoH90y9wmXk0SPwNHLUzm44YXwUyJBKQema8oK7d
0ohnS9LuH2LCy6IMPU1HnV6Qos/dD3wAkMCOhhev/A8PCHzTHkXsc46342t2oJVOLWnGwvjOnPC4
viAwJY9m+fcQBQ2fMrJzUTtg4vkb8lgZczBW33bUcusicxFNOtCQnCTzcDUT3tedPvZBwkzg8qIK
zqfEgr2Jn50s1zoxPt1lvsgLkEfBb33IFf3vM4w/80OKJ+JDgFtbhhaRGMXp12dMO66fOxlHxi8e
zZpqMnvW2QEG3qFnLnmGbzNd82YRDovL89t5fZqiFikd5xIvf0BO59qMgHB6i0V8M3iVt26DsITB
kQ1qfORoKW+S7oyAVXsh78egcR0PshY8swjmS5fhMKr2e+sjp6Ru0g9JBKxB7gUCrQhhnY/+/ive
k9JSWPHrI305h+/xzUZ5kRVoLBhVaFnDInDbVn3lFXIESn8yyOtm/i52gYWtyuEjUs9qibvgiOqz
zwXv655fkkji9hG8ldQJdN5RN6aPiiGQ3T7Wm6l5mJ6uIjPBQHd6wx6PoI/9Ev+SUoXWypOdiJok
b44Haay7aaonxd0lRKx0WTd7WYH+pxjKd/SVCvhi/2sqBthY6iNDjT/lIVqnyyVpqoOZJ/sSBBzx
bAUlMHzXiOhCmkV21r8jmoOu385cYTNQOYT5TDu7u92QPLEj6/8Qo/qWcATd/6Y2lc5GkkagcZYK
jkIxXrIhqeC3IZ5Mdsxi5mOMpVEmJAA+zRo3OFzHpSXDYS7j5ZkEh7tTot/0BkZ2tLnPgCRO0PKu
jWX2EKK4FzEdK16ti/rerpJcd0TVYfqR1TI/53Afo4T4jKQ0j7v18SkPw7/gKn1LGd2SYDFk9P56
pArJdxHQzdcxEVfPp44Y04ny7UIeSR4T8SyaTzqHXg7wSj8X+RSG2a1xTSXJNRDyq1u9hNcg5Cm+
M7k0Hictb7r33v7R2STw01y0WNir7p/2Rdz9o3MHJjYHXy2xKlsd9QvBZSd+ks+BOyO5lEithBUq
o4NPY3JWGznxBYldXEiMEpAi1A8I3gM4kk+e+hDKgBi6D/qyGygkWkNa/woC51N04CPCGo0TkpG3
mWP3C3R8k5NItwLnyHpCezgMs/BeAFjkDquEtsUXTLA9WMtWXTv7UvqUyWg8PcaFSoHa8SccIAyE
0ncXwpNbcA/dpHlgqTFXI8+4YDno1i4ul9/Zryw0SZ6Yt9jnjoJHpFzhHKMaTcXnsqyzljmGErP1
oiHv1+0Q7qkkbxBGDizrQFGD/7ilZQZiaY4xPFg0TsgRKq+ltAF2WLAuwMoFeLGYWYp74ItPzt7D
2ApwtBrIjE8wq51pdpLmgFGDm9trmDLN73rSmP3Z/YnINE5bUW6UPSC1lufFBuQWvCzhCSfSRcMo
R9awCKf7SgbNGP/bCOVK2IO/ZbPzRZpgRYqg62Y7gHqt2BmdOWZIVszGNWkySw4XR7w6DI3Fj74T
Su9bnpujBh2AuZPp56WZm9ZmsTN6fF/V3KZq0lmwG+VNti76q+k6asmKfAE6+Pl3byuqf2+IC4Cl
zz9sZNbB2EwKYAG4RbGRnU4innuQ4y1UQgzVPVnPa0FJ5vx5OmPkf+cqMhBYetFFhmPsQT/jCLMG
S4QkS16h/F8yLGatrQP63uj0J7pl6Ve8F0I2XtPIVu8+xtO6NBuW/D4udcUJmwLjibNbOiJWFHa9
1V1PgHbs6u2OzXey1zMAgEfH2DgK2zoqI4L6LRTeMZoZRfAo711f6JEDf0hg0y+ojYsZKo7uDM26
aBRr86YaC7rhBrcQmcqsvVeDfAyx0NcpTv3js+5AFNgyEzljTx/E2EuRvzAFpeRuQzlK8+sDhoVM
4P5P/CvcMkBG/bA1pZrtOmeJxmzPK5XaamoSfkntcj/SHKW05CnULtcFx7fZoSf8ePWOxgjF0AoY
0jWHCAAZTh8+m73Y4miUpIE74ZKrC3tDEQ6aTtRPTMpA8+DwhK7aG2efU5a6JVESgsO+IR1WUbvJ
QH9uVVo2/R01IIl8jiBdQN3vcw30Pumwfu0WOIry2+v6dn31D5dANg1cxmq6pWdQT4FqMz7ojtOS
lW9cZwndFf96l2TI6FnIuNr9otbj3PksB4StzuTm2+Pz31acDpPyi7VBW2qqTo4djUPfS7EgA1cz
1Z63G+sgBHb+fy3ysfggTH2rOtHkV94fSrJQ6u6sXwSJdd3WgAid77YILAF7qXlBYdAXfYT/hDpJ
BFJzioGSDZcMI4IyRPNm+h8P/pvyCdsQZa8D7VbzRJsCubSHu39U+RCqp+hRKCfrKNOwzv6YR1XP
AgZY6AbhhAwcFfx9DwUSwnz1pAqmLSp5OC2aJO26cKXui8aBk2LLGAmC2iHPW4Q58ao6u4DxXiZ3
mz+2JR4gHl5QZxIS6NCEpu3kslFQnjP63pG6pfoyaUJ1IMH1ISxVu80mqm0ROBhZ3DkLwQKSKBXa
E1fNgiKcZV8qN/z1DQHZZo71pukGReK4vichxHkjzg++SR333cbTa0ZnnwUFaj7Ic4kPWv8BQR7/
nqKgxRMozavCHH3WuSvFHu6bCey1p76RpSFmyy4I9vhnSSkI5+0hEZRK9n1nxLlIyvGdE3us4Pkq
KGscxMxG0648oxhpqlxAonuP6JpSew1DWSiZzfcfc/Rm5PxE4mzRS3MfmX5pHIJVAbZeREAEMDtx
hXmoseZc33XGsUfI0pxQNbOuv9OdSr0i7eWCyLjCC80AZv4rRqtypprdQzz4Nim7EtGYpWFkSQ1s
TwapjtKyCB30/JpvVoNWY/Dwy7YzSfJuev8iGIYkARnDRSLgVSQchs2cWQhTcRdicPfyl5ofo8vt
djPu9RXFhaffAZ7krXeIx/sBT1nxG73VAZO02RN3y/LFmTmEP5VSDcfymXdQmepbc5BHpYPZC829
8OCDF1drSeU3T2ko6pAdWGFkW+nbh9w+NXcpE1imf2J9yl+/xnAv9RScdVXGE3yZ5/shPU23FGZQ
VSxN0YJRN3ambkMyWhghWmO0wxSFFBBFyNQnvvA/DdDixzGNvkcqmLy6ym1z5NOlzQoHWPqAXyNQ
ghw6aVkD0l3CVNdB1aYyUmqvE9GYV2TXn0qkMdrpkU/VOEpC3dAzbxQtWDynxtdIqmwYWj4FV6Y/
uKaGA8r/MMlPESFFTo2woC1pbJ2MZxwup12kKhCnEEEF9KRj8aql9YLA9rZbEUyIcPFIQjYV9+us
MHifQ7vIBxPnVPC5UCE78gKzkDSLf+jvAUUZs22ac2LKPkCVo3UuJQkg+P/fk5knbsfWX6h5iZvt
hNB/xcBWfMimae8Ljl9a92OYvCejjRiaxHGEkMnRdXc88ljnWNFte0ECGceUspWlL2Voqen+BZVc
X/YvfGUGeDKUcVM7n+IU7cu9xb7OAwx2oOCfzshxyODzPKqUsi1WIY8lOTWfzhr6B25QQikoB1Vi
/yB2vBaKKzk7aztkqH7T4XaSSP2p0bRI+YM+xqWK1Kin0lPwYGYWHks4ztWNchDAYCHNdt4XUR8z
IaKBu9cCFkKcDxtAB9SScvrz2ZgROTXX9TKdzvNf7tLmcDll9aUVNGPDfi4IEokySUMzQLjFCBPU
6jQG3j7TTBYHc69aOHjG4bUYZmcNaVirm73wG7bK6C0AfppQRqVvTLvMuDkBlGUuVIviGB3hSeHs
XB2JNY11d311wfx8T1l9Pdcd9/juaRGBzK4zh+Kl9EN9SYe8j7uZOUwa4X0HVF0gx0yS6inuG5NI
Nq1EcBRsuAtTU5jtUOjqmIFAcGkz5DSyT0M5yAF/c8WIz1WNlFxrh/dq6pamel3lPnTLGrZlzdQe
bsYtToHCU1rCpae2BnRUg3Hk1C72e4Qo+1GashpUKaJ1Q+xYMuGnt1Pr5hROdWVDnbILTds6X0Sk
f6O3cILTYxs668xgIBUt5Y25qDSBOFZxxqRgCeDge5WVhdX1fLvM0c4PKQmwQfNtrdReXPPv8Kbm
X5lJS+JfqpMKmaomlyYJ6P6gK5xGBHVS+WZz8YBRVP1OE3Vzsjs/ilAaYgpNl4bxsZYwc5yhyjaM
T8VhrGsEg0jO01AUMVz0q4QvPnb021rGlqPb6x1eTAubKm6OIDK7pVz7vRpfmlD5THiWQ5jGUsV0
jyeYrisDm7V7o8oulaHdLxGLve+9IXCqCEyY36aa+gNMFntOZ7jeeT0cANtUlx2ewfMdQol9boqm
FS3nEv1Vbi8dB9wzp+ii7++f1CO6rTpCR1mUYzO+5CtHX+6tGFkh5ex2XTSkKnMUThaeKszS3Q6v
X4d6kWOtDSWxVK8khMeRXrNu0e3C4SJV3mB0CwnW15lXBLbdWdVJ9dh/0wKcLycJVzvOd2fW/kMe
otjmjugv0GTWusXurdJr3wqQ0PNZ6VQ7zk996n47t0ogZYq1Gck7cSbxCgaOoQ3R6ykMk/moqWn5
1SpXbmoBIMrtmnEOWaWJfg+jHzes4zpOIz1rJYdyQYktBHuEDdMtUikJfzjRHEw1WrMDopmVzzyT
/YU1fsER6Org2OPKCuwOnidkjygFM9ycFwzbZE0CPzLu2ZiMYCBIm26P+4489TJBzxwZJ0FZ0QJD
JacxipIQ8xKWo/Hrjv/X1HtLg1RsqKMD91bzYrMH1ZWPf1x+/VlsHY1z/mcmXNuFWvxcEjbGspI5
+8M2Tt+aAEQ7/LlC+p24R9KlyyUp8tc9Cs7OrDvHZ+sb8+pVhwB+gbrmrVgmGJy2AbRVrZjTFbr8
SR22unhXA08UYrDPP0j/nsoLtjrJYocPM0RsZZEpIKTz6NstY6o0P1n0JTh8YaL1oRpmO1p8xa1V
cFAD+qJr5KKQiq0sGF4FNcGFE1sBdRntuebh3GqTLRhCtklGXJq+8enblwICRb1FuuP0HKFkG9VN
cpwdExn5H9DSlDblyMkUJgX0biFh+QPx8UHQ603x01EVp6nSBWhWQTMdpYAD3dPLisGYgKbUAD+N
tFhjMdaA4+GNb5ycJh2L3CMbgMCgfWe7meeBjqIrEgE0agLz4MtVxbZqWbGlPe6OqFTA6wgedsAJ
gG80cJTzvu5zCajrzABwUkeW6kNbhaHJ+ZW1ZSf9PL7J0hARPk5aJRuFzxEBXCj5MnuBhKQRfPPC
ArXiR9NUbnZ2IIP3MwDEP7VHslbjNnOFp4vl27yMyDTrppaPfYSun79V6YDfNoswi8LuP/ItmmLj
SwAxkOTeOohsMrYU0fEDG4dl1XIiE9QbL3VnCZtryeIzX51L7zsxExpAyD0CMEWVME8HPfkovlhB
AGXJV6KvRDLhzarMVsDdTPeb1+ZoDPdM+B8ZgJOM/yKSkJQ+GlEmvNoyUuQYWDXg0Qvrqa0q4wGt
KgCEbkS5lTUAYwxO0B+vEI+rT0gaxhq6bVm4+O/qUxcn00Djf/P5RXXkTX3Eg7LHieLwh/crl5vi
Y16WFGcwtG3docXo08XIPezuloW6hc0S4yOTNuHxOSjKN4qyWLh/IDcy8BOURbjWqgipWJwk9nnE
+BCIypD67WmI+GygI7IhblCKL8PH0CvkwfA9XjNjkSXkE08sEH14aozk3c9h42U39pCDzN3xa4V5
uYZKI8FvbgHEwojRCzM3pbizUDcPD64Whkw7yZPAz1IolsymHUxwYrfiK7ob+4ZSGVAL+XUsas0V
BvQqJ7trcX9O+mJNoCyf3Rrg6aI6QimJiQNfxxdxaZ7rQuyqlPdH85DaTdQ5RMF7fRrSYxP/sd3A
lBiwT7Zm+TfS8PxWxiFxMlKBHCfrfLfU78IgOeF7fyaEHH0M6G8qSoosIye8Zyqf+4iL3RzWst+x
mX8SjyMfORwn5Bjxx4qLZO72nRJrCYFAFJ8WpqViWBvu3o9AmOjhsuyBu3UQOAsW28cV+ZOgoUt0
1pMFKC3zCMWLS/J1Wp6Nd8mPWLsK+383KFiTwl+E1dk3kTvKZNOYVftzIxS1XzKzmKo/Z7/xxxbV
gXPUouPB2hByVp3h8GC6ZbcxDyDb6tQyDB4ZS7fZVhvUMJPvcBiebEgzQqbRIyFC7oA7Jzn4Xt5t
m8/WSqt9u02HEoX6yNhTAMgCMObHLpWXtESqPA/R7wJ71NbG5DwYqKDDhmr/kwNsiiQDfBqWQKcX
SsGAN5k1krfmVS+hfgX+h1CYaf9kJbw3rpxWzaifU8af/Vgi9fR/FN7LlKgJsm3DS5JMixEy3eF3
COEO2BVufOF4H5wUYxyGOLoYEKPx7C8yyQ5hCYJdxYFHpqeThTs5VMtzRw25+Au4WS0LvWkx2FZg
/HGVltVzdtgj3fP/zoyiGSSr886ECHafKerVRUl7ebDHnbHIJ7HeDDjtB4M5jKFn+oJohea+NhjV
iRoL5x2MGSYmcWhZMZnQ54xsVEuQwWeg53AKSQLJlUcz/JCMfYCSwF5hECrkE6F7QoLmKwogikgT
o5yHjYObVMlPEhEXXBvyKIjLUH6L+pWS+L7+hIlzLAZ0Uv/x9OhjcsW25MHnube0DXp/NuNXp6J2
dkgehFsx3ugaHfIdLg6Y9LOCOh7eI4HE4IdJvUID8KZUxYX/NC4vf8xSCtd3PqbkvVlD9nh55kW8
o86HkKraumpzOo2HPxqzuJhJkGqB6hStRqTdaamQlcSU2aIMchmzJ0kot7iPLmJ/K0JGB7v1nSLp
qFxmpg5DPOeUEhBtaISe3XwffUr9ISFDxLrTxgaE/vZVaVe4hBdRt/Ghnzyoj/XHXH8mbcsm7+1m
Ab6FGaAKFtATRctto81WVwbcN+phuf+ei4HqM+VicRpNjzo+NQX1FNSIohICvyneynjHnyjnpOiV
jXJSGSSA3M1ZTIzqknqhQLt+UUqaZ/lf9ZyTF46+Q8dzgcTlML5InMHP8nX59zaf+ar9mUJ81Gbl
OcxD1Tfg8TNQmBQBGQMgBg1CGfRITm1ACn/P8mboIXxF3GNmD3k7VzfC4Wk88cqxoAwrQAj/NLst
VPfquNWDJO+lfxWvTiqCeaJdpfA6ABGp83CCpsuxYafLoF2AmCr0/qn/b3ipDE0GEFsK3fwf9f0E
hsqZVx8y5v+8nTRcxDF4mEnyGLEr8ZjHA8O4nEqdQGStBLMHKTP88OvaKVdX+W6Mn368wk0tNN89
bbICSLXAPba6OCLcFxhOQvJAeRr0CCgAKYYCc7WFreue30it/9MOKiB2MtTdt8qQ+EBQUixc7CmT
lrDJBlf/ex+HBzqfFqE1ZmC9Vk7tglHk8+YjMFG2CRHAw3APiRrmN1ygE3VGEmQoCrE73+dCQKN3
ZH1J1RHLd6/EyFZvlWois4TJlb2pqp5p7s5XbpfXfl3YitBhP4oxt+/6guanpPew4y7+TbrTQisi
0yenbRE0rrA07sVUGKo69NJ3VL5nvXqUzME+iOs+zBn1g3CC9km9Vh5wj+J0B4CXBf+5h8zeIVO1
DiiE5wPn0rxr9/aCBjCMOVZIJGuiG7Fr0fmtVXjnqECnAR25uqxdLjkG6kpCipPb8nrD+7YtZmIw
eyGLJKm2x7qZDcnawdndCPZOY6qpQOGCoVmPsukjGaCb0rl/WfFhIGQEpASwKPejQ7Bdiaz3Y4Bi
SMq8dUz7ke4u5Ok56PMsKNBcckFVPxP5SwKq4d3f/bQHdj8Pt71QPnk+Hbc18DmxBrBw4LVH6mXw
W36kX5JvgPIteEUwZjPciFF+jRqca4LovgqZPOIDAEwWoGDXLGuhcdCklplmDkCXTIPvMLqHr/NY
Z7sShp13cmaZndlxKAfge6fN3i1z6KL/tybH2+dY0m7Daf62A4WKy2BY1eo6sZ6Zts2TaFpL3RbJ
JLS6LOrNWS7F93rvNwondb+iS90OyNankWna0sVNmibrz1Uih+BVBjgsLuQ1L8S/fRgDGZ7FkcSV
8pVMkrkfpre+Nlvr9HbiIeQR17lcYwLzye4ckjR42QK1H0mCSOol7Z5l833PK6oYf4biz7DcxQIg
Bb7MBRef/URfysld50jvR3G4HdtgjQFk82Z3xuJhbHJQpIth8agDInnoLp+656C1C+u5/6XDcyM/
lVEKcselhKTdMLL0F762cAfiY59W9snAL+N7r+kVXKXr3AyVZj87gCeBj63A2vnfNauP/yTTVFJn
L4RaQr0cgWnAe7EDfKllaLG4tAF0+JUwL1ixaHqj5TcMpLQwtcgWIeyAXFisoeA2pC0xyQJsty3b
4y6xg4izT+cOtW8IbVNm7gXBjWXgNSDhZNraPPT64YRstReS4FtqNBENPqOI4aZ1Ao8GSotDusdN
udTcTFYS826Hv9KFYX2eOgYdpJnDYIoEW6r+7aebqvPThnsFQzpNJ0OGlOrIdiOBpN6OCnNhPGGp
S+dXctPssTAQc3TYgDU1SVC+X8i6tmM/G/XmV/6s5d7quh2ybSIHqNWuGDDRmS5Ag/oH52oZ9RPA
8ZS3h1r6qtvyLzjB4/g70Od5CcrWZYKjjZ0roe7fY223xVh1CJNc5iG2DR0dzuCikwQRw2+JpPf0
Yhm+Oc02dvgzN8D9lOhddAlCLJDTZTQnor6lid1Bgi8Nbe4W11Oxyxwf+CPVsYJuLucLbcoDz3oP
WVN4kpFCs/rnmU3UoJrgRZ3OT5ZWj4d9ruWIC3oG+LWI40tDzWw75pOzqB51KeHxiWQEcZ+fIlYk
NPEcEYtMLddbdjDf00jLBKmCKb/lsy2qvuSQRSg9G0rszAN6bH6cW2yL3LuYZRZg1dv9Rp34sA+U
tdBh0dXAUw4fiCadC8tVa3w5NWb+IIROAvyOX1WDgYhcs0ZZwFZcc2OTNDA7Zzusd1Ur/nloMQz5
ENNde41yuNC6yhFYXURMWyzRYhjoUWUYf1Qy6W5f0HgN9Y9ejJEPW1axtgEKE+Sch0k8j2qWd/Nq
wrWdp1p7OyaUbNcvhgFI8ZutfhFE1ZzXF1YTcG0pvtevOgtJvzaCqvPKN9UF92jYFNLcqMlryend
bym9BcYe7GsQgmZk+sNFGMY8RrU86dMNE9Lm/lNV5Wv8VA8ZfRRfIIOt6uEumtyvJjbItLtjEWc9
Ns86VPLfVLIyFw8AVYLh/p+yWiZkljiLF1hftlW5g0EH7j/4GDH2B865k5FSE1L7yzOLj4rxb0DA
pYr3Fa1uGOwqfmYoB3gVpJg9hRy67O8QJrIVTemJ2oFNVgLjrFHWfSYD6+euzjpr/+q8xa0+EzWP
HSAbuG7iU4G3TZ5E/gTjUEsPfaZT3ZMzZc+EJh7pyqIPOayh9bGbo8DQW2qq9Xcsjd2msKR3heU3
3jQ5WwgqgV26rFHyDwyugL3yVDic660npJWWJ1/+1iOFhlwk+Gh5cdKlU3XSOS3eArtd0Zk5dGca
nyQTzXPDXItKLYyygcY9xP2Zr9n2JSZ8ZHVSLJQyVG3ITHfqnh4cUCbiWXGXWlKuoeM1Mp2ZoPhO
TPo+a/ZCZop/afiT3Ht2QIZBLAUN2xflCdfFTOKC1bYhxuZMbudFMUnPemQLbEFQg+BqDKyhKlyU
1nMnTZ+1gjWaFCXJF7hoZBtOue7zmyCytQbjkh4zTA6nLfQ4USqkU+JPdP5J6OW7XM8ibVN0YrEU
TXB39dXBAd8WGkNtf2O5ZuSRofxO2FpPtbo/V06kt3HAzQW3yrSx+6CMJ3ogbhuo03e5/SAdvRCD
yN3cL4DVEWwi2poxe9P06TwFRckp3hn61JUlcMpFyNS7pDZeqGvZ/bVGDT8urzukjFhiE4MU+kv4
soR3XsRyWcmKK7If91onRao0us2Rqx0XUuv8tcAHcwnQBYxH/sSuGdvNqMuUc4rHx03NEYZveCX3
7Q3lZA6RCBQboqI4zva4IPgOLsyVl97jzGVZ6LDa/MKlnfc08kdYVJdhri2Z3NzVBy4CSnPdagga
GI2+jzMeZaQe11se5idBLGbyqtL1K79oceq4XTqTJfQavYPmFn6pZrAvRjMgRGOnePGOXA/X4S9C
RDg5pRnDZQXx7y7QL2WVTA1+08E5zYbo8FP9wHtITx/2x9vXPBAvIYK9d62leAvj5cE39GgXQnfz
iS8goj/dEds0N0YQizL/hMhVEgX7SAc1JVH+oiQpZzTjr2tgf44udzszl1trflZIy5zQ42keiQjM
VpANHa1+PyPPfMbHWyMKWOU+tpg5+OobP/7MuvBhBf38hknBp38NUm/L6TWpXeCYADRoIOgNfcUH
TAtnEj/dFCs8jm1act0tacwEJa2s0K9mtKKIqJjArXXns62UoDxaTF5Abx63wbNYY8Kmg4uqsLoU
pWCnuiaAE4O04TrfxhNjHovyNoerScGdLMFeS0ONjfFhk/itLOzYm8hmDTH62O0j0yyJtuB3URN2
JaqJVSF4buZCi1PhnVbZlTMd6TXnFcH9A5W8x9bqs1QjnOV44mZaXNz8BpCTiTlITFjiQfeLMiWs
GOR90NbbfYgvWEkLxnMK/MeikCnaUeIHFmvHVjAnPl9gR/qdChBhcTSYd7kvygwD5AQUUrL2ogvm
eChmOCMxp7j9PBdmGwL2FzVfbTiFh4JiJF5aqwt4m1HxsIQoGyQDrKyWzjS7MY+3vq8b8eqq28jt
MOOJkXceo0vNMej83lpT5zDMY0/TfIfAd13Pt7riz3v2iz0MsfOt613x1XvcsbBSFVbJuG7rPfXh
mmpujyQFD+jjh+33v0zrV6Lz2YmHulzHp3LIOCvSoW0YrOWnOqdO314CfaReBVRl6W+FQaWUZkWg
REJKpV0znKNFkc047k68eqDMU/ysgw2jwm14+DjaAjY1hAc0YRY0BfPINIdr4IwubUFs9ZOAA/CF
AYlxmI4z/k0xgn3xPybEGa76qm98aI9lv2dSKqcRmhFRRd9ZZOWg4/KrJXylTo7EGnnE0cooEuFc
bsHf+R7aK0r9i0ZsziR6gp6+cvzSSqP0ZmiIZp/17CDHKVQwOtEQsQXoWsu4q9IjMJyjxtZGjv8g
G+mvba7rqe80q77hqo4NpEoON/mVZhuRg8+RnPvtbL9kQ3Q/gsOcEaNprR4QQMbzPbrxxBCUYShY
x0mauNqPIv6Zk0ys4+bGmPoQIR2LrrjvYHU7YO5iR5qGKbZyZRoQkIg/2zIaA+vabjzAp03CBxfT
GODWNNPUWeEizTGfan5B4fSxmgUXAl51DzMx7qcwZO8Rojc61VU6Fkg25Kn31ASakdiAkahOIkLN
c74pwGJj5GpKkqlzQrolTYlhKsaRVCjVUpvs1O8XmXtItmQ0t/POUNY3ocuSvlwKSIVUHy86ZiDd
li2nSiJDvL+RV/7uxmUFFKExZ0Em1LJhknTjqTzG4YpeR7Jzqakdnn3nAw/fE7npt2vk7WOfmnA/
g2kxlB2LKm4sl1WUqbN4jJA5po2gohoEgKs8KI6NPaytACBC9NAGlkznFPXEDZ5uUWiZR0PGeU1u
eD1h4WjnoI9gHr9PnsJMeEPoqAb0QkLzVQPr2qLoMIbUT/suHBIq3nsJHes0Q3MsKStJwtGvYO9j
Cd/iZSTjDdrHAh0GCmIfx8hNoW/5NONaG38JKx5fi7EXT/yD5OIjhHE6Q6FqFLZc6z247YBFadsl
E4DL6s8xaZ4/vNHWLtqEI0ukYHGULOFPRCvaPJup0TdBfjjW9IV2bSSB9PO3mYiw9RTKEssD4/gH
gz3In3MHodLMEizh7rW+VDIPUokSxq41xEDtg0X82ox5OBDraxAyKs918AdezPvKBLskdOY7/yfx
BwPHUhyrbucajqXsiMQVg+QPFtu05XKv4rcV0fgmMi34ttHhWYnE1FgT9byMV6g5C3g8L/wFej+f
Tk4ccRDh7YYOg88SKEDu8YFJyyj0MOsEWbNWqYEPhj/kQ8pRqIcGa6aGLGUmfIOtL28J6MooKRq4
ZyvDNQgLquq1S+VXF7fNhN8/20Hm5KcglHky6228QGZeUDgiu+epARuE9S7m6SHSR2Ir8ChK31bS
XdwX3Oq3ZbJdtGl5n2bWxzG70+P7XgWnOSzIjwkUKzGLGBiPRCnWhUB1m83xaLaYkYyQNvZbAVeG
u4vtokRPzZCAZCJGlr5I0AeK8Fe69nbvvSiwJIXeCgGto1yBgrzLBF8gYEeWOW64Hh6A90UhHVKH
hjyGIO6hyhBW9WHzUcSYgcJqnpchcmzK/i6Y9ve+Orqhb23N5Mu4m7dDyV87xfICcJ1S22Fi8sWz
lru7Mk3Z/bTaO3ANsII+FODWoC+beYJkpDBylOlNvjyuwxRx3T8E0d9JAahUs4F/bTLZtKqC6Nqb
txn1CwieQzrDiYNyK93DjMqFwvspKPwd7sekxmdwJeEYQgywejb96gfAqEUzt1JzUJvW+itqPZdM
zcfc+wD4Zc60WqfN2Ol20Mkn7w9VpsBHupDT6GoKzc4mtF/En8NRNGyhik6C40YhKzRFojCXwcfW
MzukLZckYPlMQLn564jzjmvYkucidBpSv7ar75jBiwQl+GLQdriRk9R0FWcc+VLJhByCl61s29sr
VMQJ3PDxR3Ow84uRNcKyXWqlsPdo9A71LFah8jsrY0S6YFAdeERw7+Apnquqdibn7xoz6Imq2lWU
hzPxFpgfix8cqYQPIIpttARzVycEq12KrDuelyASQuObhjmDYMSLq/8v/SVOmCwQxMSOsGmsREwy
pgjCtmtY9FtU7WLoQ3MtWyBLJsCnjWnqm13xyD7wb58fo4XMutnZhmhZMh3ehZOOp1FRAIzqLmRi
qy78IPQFSnp7/KPy2DaJcq42JIzdLONKk8sybRUK3eLVIQSZS/w5yUBmSe17UCWa4xBfJ4TXt3n3
fRJOxV9GCG0DkV2MEJH37AcudAtKeHXXSazbuVUlEBCYzGPZK6A3IMAxMd0vSFnxKOWCSlRdBIG/
BqIMKBCbveZGtJhRGes3DPMOHPj76MqQrXG/c5XIiXr54cal72ErHKDcEcJFqdoPJCdq2PsEI/5q
svousLiclhmQ/kGHhcYkzrfU5Qyb3ebBHHdd4OjVlF1dD9hlBkcXq/493L/3q6vJgWw8biwKqCgR
Mn+KwcrVLqydzKm3Tpd949HspLrblFHSy/UrjUMHa9dWywVj1quEf1776E6LgUeaCjt/OH8+jId3
GnEPVw5NAai2sCOigPT2/LAX5sl7imu6fALL95F/YRVi3RKgZJGLCNv0yTDuXhpXvITMQPDvEqIH
U9kIAQYNbIomdTkHVC/zbUZ4Auga0MNx8MqH+uea7Jbye5PK+eeEleXCYtDEwKy4cdZrba/Ogyjg
fk59VdNw9e2LKdikTRJtufdJI+nMIJ/ad6Ndm1GOB88K0kEIL/jmwvT0DlAzuqkBJY9sqadVEgNu
/q7UIrO0+P/ZyxMyT8f98BGr88D6HOHeKEUlKU2/Nu5pY+eeJurgZGLnTTUW2auYsYM8dtiEFXEr
vRLyyQfL6SYB52/zfm7qtaRo/LWrfZEi3bVOBgPyCAJh+YtgktsLVrkDVt3JkQX2OIUES5Q1tERI
1zPygb790m8TPojqF5Apy2Kft8rKR/+bsGCTeD+d9lxpdNCaeqjv9SYBwR01xV6KiUvXJlh39zT9
ytsfaqdicxURzFqWaN0JGzyZ+WP5+gcmGiIJbLBMmIvUf/w2V3RI/uJpMvDmpGheqo4+aisvRba/
He6uRKzzAQA48BelK+zbwW8WvpHWuNNDShQquOHb70HhAEYCfxtiz85+CAij5wT0QE6Kl3WNXnLB
6zcTRcBIiRNQ1y5+jYsBDRoSqJGy2uOumc+rPN2BN1qdKeOyWS7rn9LaxpmcugS5mceorUsdeo0X
TPXltxMybs1Gj0rqu5dJiyj0W3Dvkq6+1P4uQVQytUVTVXwkmTHLXZrU0W1EED2rx1SUHLE+yvDe
ifk8wbLOkGgMfljK9KnXhsdq1nSiMGkNrGo8+pIJg4sY6+E7BIGZRis4usQ9xoZiXY21EgqloKBR
IiHJiNvzOxLfVjCRlIKjfwFpCQS9nTU4LcwMdQfRVL8ECFFCJ9mP8MijwXM/zJXQTnFB5oHkTRjP
jaxCUMAEcxm20b8yyxOafiXHQJ/XpR6iX0vxLam231a4/T8zNf50p9W+i0nmRnyDPCT3CWXUk8dE
jcKHh1CyR5satK77zvwNp1L9Gi1nHthEmgimL0Cmt6dRRfgU2nuiiKNjZWc3MqWN/qAJJ+rn2PK8
bwhuqCM0b6RcLI4MFDRfDpNRTQvJq+jyZUPbLxqq8DR/2fvtmIjJsUGKqFVelW2a+1MbI3tj8WlD
mhlNhCUKneGZ1oDfgX6i9MhNOcYHONIX1A9c7t+C2i6ZvOjTNfnLFnIRo3fjce8GMTpXYO/gPMXY
W7xi4oqcbE6mxEV7HySyPfr7t3ynA+eQfK9BszjuJ9ImEW4TzebUVWnv9VEsKJoPDaPALNKKyFj0
PFMXgl+7AYF8ia2O8Ov3xt6VS5bVi9VBt5/39OLL7uNwejN1ALYy0rmaMqpfWopRX3W8MVAa1hNg
vi9no2qFUyb9JmQGv8b//bN2mtizvf22UOSnmnvlAB4YvAsMwcKRgffGp68Ws7f1fNXytuHl/KsY
YU7E22aeaur8Fl0hgZedbbznp4SFOEVjO0Hz1UcIP314wmG+g6m1lwK9fzoiEmliPXMEQ1I/3JbD
CpBJ5VxkGr1IcSA7rnlm/uozVrwnrKfSJoLheLRJTvjVhnXrbubWj8HTKTeT+Si1gr/weEMIGqvP
WDlWpVzzqiU1CBSa9qXzQkte6L10G42ZnWXC7V+NcnT714GdX/891WQB9PmapoD+NTpWJa3CXgiV
4b5JxnAiEA4UR2HjnzJDjiRWy8MYhw2uCjtlC81KyLUhjBJHsTGvOxa/VQ7B5TZ6Z60m2JEpgeGw
VvCREK+whHLXEfcU3g2VJc/B9xaPqdpM57EHDWKQv4y9SWsefjfQDLza3P920QZrGAGH5l+ltUi2
95J8dOqWZmGymxhKPhjHfPOQ1DCEJ5htIJ1In9bTRPtpBjmaJiDBRsE3IveRPle2b0Wb2sihO+vd
djj10jgXUxP0JCDJ4hHjQgVDMjTJqEgBMkXDj8j2sD8GvGZ3lmFa4uXdcOrABB8YAK0iEG2sl8b5
J9jecJurTc+JbcYVKfG49nuV1zeaIA5qQIp+T3GUT9cCorURWhn3K3LL4/Lba0FPPmCBC8AbMSF/
ueAyblmS9h+s4aKhbkXDqJD1jWzn0Pfu8Qh2HXdBZYaF/tr9caKuFG9ir5wJoHLVCN6gnE1ZVNao
nh9SwPKc1AJ4QP8gHTf7tsKSSdkZINq316y1xrMrmg7R3lVG/hrNDEl9ZES/vUhKdNRpUXJx2Vav
dU0UuOZ+qoNP5hE1VvbyGgMVR7RjLKAIjU/jYNGEMqGUg3UGnb5ZISpLHbU+K2fJOAGf8nGqwMk0
3iuAPXjcSV40pt4kjC8mpnmWxIy1XoXkCLdJKjJIDo98oYexMNI0MjzTabrNAEtx6alif3JOJxm1
RpM6fTtjPVUtWxmEA7RPYdFWXf+Qg8SrwiUofKH/uPCMYgqTSdydQ1LFf3Zp5UT9PUdsNZFJwQ4y
KrKlvZDTO98qe5D2ENeQj8j9s2unDtav+KbuNYRzVcGnjoM7ewYmJZVuakVLLgKrHzQJXhc92OF7
vxB6VYZPJZJB5xzNQZwez8T9V8084kFswErTJUlb26w8+ufgylkoo7n5LmI+hNqKKNhDtxIm4ywI
Jcen/83Ia63SAGG7N7APWnBsRvhZMySORhdtzlrL7jLNOJYEfLkso0YNCNfhMBKO23UHvrFbbVAH
z0doTW1muAO+jOn4kZTx5B6t+TVB7z0szZMHSLwj6nlBZ1dJiulXgs1l+G0NPSckpvCTxMk0J34V
dVBsAZaOZZx2CUDYOn/lGwRPZEx21If8kvvYcmFplWBdZXnaLlE/s6Oz+i60hRqplWRHpCrMqLYU
5ij1H9imvq3xAsLjeopQVSKOA2CbobRi8i9P7xa/uu20cZTeSmnZAcxQ/ReZs3pRv8C/gXVcIMcs
8ylzBLEGDm9KcOTU2nuMoCOxTFK5FUsaJj3QBUWbox6JRItuksoCzRpNynW0ShWhsKvQeZlErJe+
DSjnOCewlbFrx8FJYYgy/4qaC8K6HhOgogomsyKaj9q6C6Wnv2W0yb59zznyanWGKQYWuakcJbtf
UTmHnXVzpmabP2McUTqqfFKAuj+N9bWdkeNP5yobc7yxJFp7jqBcQUCdjrb/hYkkj6kaeirEulZo
bIuzuLBqHWBZQw2RX5jI093HeYcTyEc5W6xxLXgX2ooPuOWIsF14L4kiZxcMGKvneG/J9ZWfKbuv
DGCviRHVAzKpGdhpumApmW7kk+TUEakqu4MLpy9QLitAAyCXQXRYDtCJ9tchu7ccfZFUfZNiIph1
TM/icJ1y2UE3ITdzYNjbxoEXr0zfjXw92N5Y6AwGL3cvWU3fcWyToa6nycQebINkyDcC9PQz8MIR
NcyAtoriYvqiRmQjl+4BcgUPR1aZDn+TWrkwSqCXnwG/9DD8CrbmuXJQE/9XP3xxZ53MSo5+FuWt
rSe/WSZmkIgGHPsoyb8Q/d+A87pqWnCfxASpn2xH2mj+Nkk/2lGSDe6M0hFgNSz+o34VVy403yKp
aBoqRWz4dGn/8DHfOsdpkaddjkwN0D3+JDzU8DvZTgDrvDz5o+vG32H/GjhAswWEX1x0n/1ReM6X
Zr9ak38/q2qWIMpLphPFXaKntttEl6aG3Oayj2Njl3tGQoIUV8rBWTJ3OARs/rUEQse+1MVa1l3B
tiKzb56KP90grDx62f9s5DeNZU8Z2dyLZpEx0fmJn8tvsnRyo1VJ4Ab5uu0U++tdl8apsXuogI6B
k/V87kvfM8J7+Mey/YLYyxl839h8KLo/Ug9pmEIS7vtilLDjzOPMtSd4HUXkG9h76di4lvxhkbSB
kaS4Ujrotm/3pTWLStbLjy9rOJScG2Om81Ge1WZUZ9C2aYeabm3z3Yd75H97FF10O9MsGM7hfB9h
uT2OUT57YWSK2MPBIFpU4OqikM25tu5Kb31B24qQoaOi3obeQFKX2Kd7V9TcgAL7aNvPfIeuJrPl
m8r7M01Q3RmH/AlcKt0DP7xzq9dPBwpV0156tMhtgEsrS/sH+0RpzwSHNUba70Y8FXAYsREXBTHU
+/8nwEeqG3zzwzNJQhIwTf8BmTuWVmKuA2KVZe7wdVMTkEAs6l/uP2D6ALxiAUFimGXfYnEdlQER
aQco7TgHEZYMeqfJLQH1SzEw1rXUbmRI3iBSMQKTClwU6lLcU+YAwwjh3grRr93bglssk5gC6c52
w2PvHmoeFXQO5RminpOMfjyYf9jbMArJbRmbmt2AZmeErrR3WqMlQLXMe0zTtcmNSzXAN+wcpQBY
byerhjfehEPp7ZBAAVmrMrXTuC5olBpb9N6x6iB+i847oVVcjp74nZ/DL5PsiGEfvHCNPAJF9uhQ
yw7EdE4K/DcQMUynF1uv1lhTijQ9eqiO/TM2FxWGSraz9D2B1MVFl4S5IGNHfpvkEB3Z4mhg+arY
7vCNZfkBidQaoy21ZsjXRI8Kur0cnV4x9K6OyXXOgzb9HnpR0mf5U93VWxEM9x5IORr39GBgg4vW
+JSsdJWZbH4Y9W6yMnfWO2pr9rtcH2n3ksxYodLmDWkhfpCIPKZd+3fPUqRpQHoaWzeYdTjOpWWl
80MYmJgUgYuJwe6iQxClnsyN7hqRuQ3bsuti3e0rsS4yM2VvnfUh1hsBvP/QV9CA66aISKJ2N3dX
uZXJnlo8hiGMUfFKpDPoDYwiyiCpR6c6JOIHTohYsFC8+MATorfHDGceWLJJNpchNB/lM0VYzzJA
vtFBoFC+VyNRdHrDoQJg7umD/WYEPkmCM8104zJkaz8parxacgFzXg6mxHumakk90TaG4ANye5r5
bYnVuGlPQCW1nWdNVLnadilwnbLSK0s0y2EfM2wCjQQsQePto7/pgeIZVuMhSdrhVrp9hp5c7WsE
C9IvxqR+9stHPvWDavAFK1J+X+MtSKpH+8dsXxkcSxE70Qd7gEpMz8769iZ3xXgOgQWMf58wI8R9
mCByNq3kX82iDylI41iJ901B8YDZbYyAKOrAm3PqCWv+P5xlSk98cRbPBYjrOyo0Yyhq7R3dkLOK
HUrNIzM5MH0LOIrg+S6D/uzrH8yVc2U4mZYQQ6vAXSkLx6pEBIzaj2ZrDOPBF8v6jFLNUlnIBS3M
lnpwVWW0EF+061i2uNA1LYhmQxR+YWIesDWjOBIePsnQtAxq/VWS4dPVMX4iDAGRBtUbQyqitIcd
QtibomAyn+t+NernROAjCSA2vs3h+tI7BbA44kUUGNAW2PUuSJUnHuN/uE2M8VgETjkPXUIU0a06
2Em3+3iSiRLHxjyXe0OUnOZ/dJ5zYy7JC067sBIsB5Ib+vNVdAntJUOKacisbb0fgwo3EOa/+z8O
ZOSa4q+wqFd8roAONYiFYsNXqXZ/cuDbrnBZ2qLCvLFqqWHFbmozd0l7C5hW1I6S97R9UMnvvWIm
Q8Gxiq1bRFl6DBgnF5AprFLNcKdZs+z2MvrGjw6F7nMXCRJkKkk3KFuL+prxYbpeC5+CVeKV6/7Y
jOpw+CPR/H77xhV4JdwzVLL1VrSbt7VKIcSqBASEHHnHaHtKPhR2tl2VzvRymMZCCVVpEgevwaLz
j9ONy5II2gfRfcbdMhi5UhJdUbwE/JKqfcZXUp+D6MRP+4W3vTSC+K9rLbLYPzosaptpWQBceyou
E1kc9wkhkIJbjac+0qGPxIsaHVX7+oXhj8yNomXX7pho/8NSTct/ITq0sS9CWYi5co5h0eotpkOa
4hlJIJUDsD07zdrgQqoku5z4bKktzqwy7t2w9LopU62Gu5h/2sytVeL0JBC4vO3j6XH3ZAffnsE8
StyzKp/EaQ+gtiZIq2xFNFFRCsE+yofeHyYUaI9pm9ZgGHcC0ZpqDwRbRTlYeSL2BQ4Cf5JQRnKV
tWzuO4VijCGgLerqrIHo9Knz3F/wFfuU0JjUsfRlxbWRh24hVcdJz2v3MFmj5zIQEYilaHukaSeW
Fsgd3PbginRQ5ISekrEQrSAAEZndvAcM0vQAmbzk+qQkkPL+KGyfM4mUtxrhY4DiEbGDmY28gJr/
a5QobpPjDTlz71VtAfNq0oJB6Zt1lklp84UaJooO7RMejKBYXwP655AhLvNa5aauwQdgF7iJhQoO
FF4BC6SCZVevDr6ZrbCOdGvDJNodrG+55GMMqlvwG9i+wUVbWtn3Nj7vAmUNTIMN+50qSq/XVcva
/NbJjoTF1f3UxjO86S7qS+ch9MiKTNq2EhSJJiUqFlPSQuForKdn+Chl4BvGoyNXg42d/rHeNeCN
BiVjPhiuvuBU/Ye3+40ZxKbdgpKzipMpc+qqn4xESe7oKL21PtYgZ0KBYFFw2k1NKLbjbOJ8iVNK
KyqNwv/htDEUkUR6MvoMmlmrvdjyHTVoPX9nYwSQoH6Wvi5r1Q5csYiWdrfWks0AgW+G6LziSW7k
HS6TTREACEpGCaW6kPWdK5fPf/+kL1kAZBcWZQhsUqYuVQRgLKkp8HP/pj38GXMq1edLP33QPpmE
1hHUTAcuRviHKS4peyaRtqKeu+pZ2UpumSl7OSayCkx6saz9fasqAvscrp8iQszuv4nG+tD57awM
dJfWLCb3OOsIPp4rEuiNDWz9cp+95JIIx4IgOC1msQu8LzzeaN/d5kKd7BxwstxSxyozEOOVRPYJ
crOARN0Q5letoU+2DeIWqFKCSBwnFwmsQ8kaiqM8DXt4sqNU15qtWu9YJlbiHKKOmstz+L3ozWNl
YSjn4pTuXvwGJyh+HYqp7i9VFNLH8NBp0x1oFqugVHASyktNICAQ1Oo6A3uP+XDnsDxeUHwHvAW1
SxYNKtHfWZhTk2f9zxYBZd0bEOV1oye7huA12GdYKbvk6PlowfwgHH6g041Oa9mfN4xkWiV/B/wq
0czqiXRJ5+NZ+rNInupam+FwiBRzto5jZeR4ch69mcbJniXEKIWtNJ7d4TXzDEcn2KKB840Z1/tU
WAvBRtMINaPWcVyraybCd6rQq5pLO9ANl4MFMfb3aaW2bxgJCay0jK3m/hFYLEbtcjz96hve+eGJ
RRXPp2gJz9EFVipY25CIYLoOn7G0J0GdzwUBpZ174O67PyyIENncRSH8E3nASqXkQzvMmETUebFe
AVQjaqRXJBtOSkFzSwHudUgZrSDuFtAbkrL/clEe5/Xto8PgRUolFproFrEHOhLCVBx/l1IhvYPX
fCtNK/qSC8rrmNUQw6iVB8lj6MvGQXmXfEerXUigOI38riPVAhFFWJ+aUp7uoV8Bi6PWr0xo3wQt
IUHY1MMlYnKxQxqb7IwnXpK563MhTBf5gyXDfKIbgGA3S5SI5+ha/FQgh78DDWKGEZlYW+4yoYvg
3wZyZyFd/BdhaF88wpzydRxSsiDRan57H2LR213rj964q8VN2WAAosPO8VX7cguQlno1XqGANXMr
DCa1+AUhFdgxTcYNK6K+GcNDC6dqtR8UAsqKA9ivRsxDNXOfuMcOT3/9B6CVbSjU7PUq9fBXOLVB
/vPNi9qFamhQYJX05wBHC4P/dPTYsEtqQl6VtyRDTv3J9Q8W+T/p+an3foi+Sb0BUhTMBHeFJX0y
PuNIc2UDcopUemjYfeG1IrQma4/F1+rldCP0kOqC10h2qqcCnw25JqcUdBzp/y2PcnKF0Ua/TMlV
7s5gkOEE6Zyum/5HBu1t0l4xjhYKN+sx65Q9QIX9b6uHgHD0uTSlCxKOlAzMcb0bD8SCzz4RvhGm
nZNgDiV1Yssf2yXpDpPJ2i4UgCSJKhDOF2py9k1XTdyY6RCpq1X0bd+4b8zvWwAXLY2D4dCQrHTk
h/BlCMKZMlip7ST+krkhAaMDCZrE6hL32FW14MKDljATFAvmo7AbW0W0RR4+x44zAikJcheqJYV6
8XYmGjE4c+LXQlOiSw9+/eCaTWmsz8VLqHhpvvfd/vJP4JWhvGM7WfHupo86ZGNd2JJaCgb+Bgdu
yU+Ey35jqCf+arlH1B91jzigJzpdPi9krXrEf0VtckoNC31TM01YgR/S+c0r/LG/L1oWsl0Z5ehh
/eE5qlfDVCjEWHls7NXaAUu98n0mxIWlPAtrdmu2WdSWxTqvj05hZ7XnjBQ/TK9MMwATshY5vvey
clGCyVWC3jpjMTUDvOTkeqgnPIeYB3F0mWDNHRs+7Rwk1gCHNKWoGFjyjT5LMY27DLr8QBZy3+Fo
p0BC3jWL5tIQ42Kx8Vdmp3Tszy6gZBWU6d6EX11sMOaOUOsnLEqKGHv/XCmo6LzunFAMvg8RcElG
L2Hh8Levx6h+PYg0mXTQS0aDGd1iPb9zclhgxls0TLTOpel/GsHzwM6qcdolmRjC7rDKRwjT/NZz
8Eq8cPikZlqntkaDGVmpW+fBFJVPW0OQk+loznbrFNVzTj720UVlADdSS/VhmSzU9XFk17laLu8w
N3w968/Dgy6HBjYoiyeizytTAny8ke8bxEVr5lGUdbzxEesM7WViYfSmf1RNLPo8y5ngiG3LlQ2T
OXpK7titZnyMsKe4eQm0p/vkWieEcRlidoSbpZlswlazsewQXaLEIz6beJNDrl7siVUEn6vchXgJ
PcBonnr6Jdr+MCNbmOXguDMUMPP8vUx4nGRrg8aKwnOrKbfTRWqjWZgztulWMYcBRs9QJSPAuDSe
+Hk07oPaAGY5QE5i5LwRaIaM1ZePsPDqkHt0wN4ElcHM+CZu1cudpYPzNRUrtRygX8g5DsePwIFe
0WSfvj3zB3LA8Pe64nF9D8aRTDHX/dKXCVBh71xAGNTwbkR9nPIzOjQ1tkkM+FRXZP46ewHfFbEW
OkRgJZAH4nTQ2bE9rhAvx5fOoC2TKKHvZYRClV760z8KCLGcNAm+93y31o1JO/vWg1qZ//25MLB9
KymShYRQsSBUr9Bk6/cSEFXjjKiG2wXgcO8Kgp28FFuOHqTk6o+DnhyN/60t1t122q7AHnxycTY0
RHKjQGMxdhCoq4CqlTkk7yLS+aE7yrspcrHTX30bADEY5wQVXR6+ZzBpIHQ+FKAaXkEMLDjYkJ3H
m/VxctvkXJG5924ZeispDlT4b0JUTpo3kthNc4ZYCAn9USuqjRaw0mEQHG/OGal1v7AM+J72ZZLN
kvXwKs94A4M7oUMwT9OvDUF5RbPl05+q8Z77LIZtAERh/Ox36proeTMolt7Hllf8HLGTNuNrAikV
GZ141goRqWfXp6BbT0IA18n654Hgo4IH4vmtKZqHmMMxLXzI0/Kfvy+N3fOui9mMGlCJ5TKd9Q2K
2VOJa+uXZZXrmAbePI00QbUhOPwieX8IYTCCWTPEiEd+Atn4EAsU/2iu40WwMk7c7VqAcmYsxTid
mea98o44iwpJ2PTBnsDJsLSWNfC6dK3/+XH5i7igYmusqhRp3HsDOmzzVZ9nTaRSup0Ny6N8DgQm
ObiDw5VEAW2ySl5bqNq1KNuJR4jatzMesBzlC9ZWSjiNy6TrqJAq8pHuPAM7NG3MDqYJwjznG3DJ
I4lQTUui37tB/1qkki3ViU5oGAXrMjkAo+pOxXiBC/FhkNEWMQMm2tPtrmydlXrOKtRyMzJvwIQj
syXcjkOc1oa/sL+uOrXucv0i91iinKti1n0/YfHbKnc5l7O7giXRAPPlr3y6HHAmq08pPpWLcYqT
SPwyGWK6yrV3EDUGqC3+wfeT2cu+v2A/jnXvQGqcwnoVNsaRqHcb3Suxo5B7hooTppPruch80UlE
8fWTWi8sqinB0X9sQU3dspFRCsbb2qOQLtspj3s+jsNyGRqUBqVUmvBPhXib9j2qVTL9qUzyPNpe
jfldH+pXxdoQlYTzeTvT+lFkIPpAF+eO3Lf3trvHYNwh1hYQi2nXHwVqLXFISpTE0NOG6rLlyM9R
jXwausnUiddxA8i2sJjgcse6vqQ6Mvq1Q2XVBAfv+/H1p6vlYVMYybsctOXUqe1By2r3LmAby3e1
oJQ0ovoM16ogI3DC7Q9u9YE3V6TAmqS65rZSeK86Nlmvyvk0Sax7bLgFUdwQGtFSElcOCavRjSp3
C3z7IwZgq/I3KBQ4fXq5Wgnwu48RYoq2eLv1zpQr8I8Q6SHdzXD1y//v80yaeDI9y1eOScPfjsue
S2CfSwQkTSREMQfHEMMoRePsVR+UNaDKT/aKsT86B9dSAu6EqQRhgJOIqJx4clx7WJc+CdPhVvDS
2h6G8J1w/u6DgQDfSD26lHbwWmXzMfzFW5aIy8Jf3rvvDv6xmg1moAMSJHbFmvsQmC/k6lMnjK5O
8oq2MrAbdZbLmYa8N/XZmDgfS2pa0vPX+BGEGhVpe7beO+XF+0lymcjVpzY19YCE+GOsAHMFU/Jq
L5sxTyksum76HnYkTy8QHSO7lg+uAAvENtxb7wkcX43+UCc0vEH707MG4RtqmSjEcxmvSd9vjAM7
tsJSp/YKfjWcFQw3e6Kw0cRREL1oKZ7z6ZobQLJ1RFRMCASIed/8X7h0dbFS6HWlJQHBHvx8lNJS
IrA2kyz65z0GjsUFc/V1eGKzLCmW5a1giKqly9PkSRrcVlD7MJLhK5AM1ARhS8+6RwH//YHOyYCd
H9TbgzfgSzGKv2Qm1DTYmBddo7ejagzszdL+SB5dR4tblXws/ROLaCWZfP6ChMdJaaRYJx1mrVUB
DUyNMSWs1lFaDkNq5EOpBM7QCzNou1NU8q/Uwu/gvWCTHYpgayPau+5kCHwN1YGS2JJ2vdqnFFL+
1Z9M0oTHYDQpNJjOcUUKx0nTVvP8x/8MDMp+8aB+7bHiShXhdwqURYPrO+0uCHc7FtENugmjtwVd
7yeyrE5T2QJJKfkdZlJogTvtz1i6RhWZN+OAXRWwvRDuteaZoCK5xkZPdSOX4gnO64XoOkCiTR0y
0lwL3ur+FOcPuDN4qB46E7dLKC9tL1/FAA0+w3+0/cPKezKTDz7nnCfHju5hzxdYqpFUct9UDr1m
I5bmWQM91cipUFM2EDy0+jOMXfJFSvLHbMFomHQ2KMzfODwwqkcA1Rw/o42Jp/KrP0hAZmH8t61Z
hxG6Y+sHidg70bJgfoydLfCTiWlFBMNzyqzv8P1x/WToE3wEH286RmqBDAkIOv1NhPDIB/zqd/uo
nXTXXl0Qm06ei5+gI4gLUZ31LogQetRB4T9fyV/mk6c1qD25vc9h+g14//4/9Av1EGCquM1qMl3Z
wEfoUBDPI9Kk3jnDGvOxO8lnj/3j1s45+CmZrUaYDaVfUZuXQvyxzOleKAimWL++ugQ7qN2gW/ys
qk+rEr26oM1kP5FUqlmTwpRS3vvEcQXs2OrqY/89AQQXn45F5kNfcSuPZswxCLTQMx7HtHLVonT5
182M2rjjw2UP2b17662c9atb945Hp9++fbjO/q7/z61nJ6DX89f5UHIsJJQlCJNvnFNgEjthQjG2
nOKQea0ASKcN55TORaY6BIgZf02Nkt5j5UPQzflcC/NO9xLuNgW0KrwupMj0LOEp30BU+X7K1ipL
wqUrUoaa/Do186p2qCxersBs9+hrVuRhb2POM6/h+GkRfPDYsTlWB8Ad4H4n+qtravQ7ZQTBjzn9
lHTG//kEObmPQ8VB29u1w7BsjfzVruIpl8YE2SZlIU8hlwUvL+cqniWFptWOdjv4sdOTP3fUtXcB
iQqtP4iC3l4HQG5A9KS8oUE2uNVfKxVrKOnhThyKFIL08iHVXbb1LJ632zWiSw1G5EA+n6CEx4uL
9007xMwhUDVSaffIhteZNRIMKt22KnXMduINffpUtIhJ0QqJ0IIQvcXILDoGtk//GbwXee83CsrU
AkR5DYQD+b2KDmUmn1jquE7Z31gr3rNc8L9EgtNtf/8Ec+desYzU5H5Gp1lKvTKJH1Y86GzQncSa
GLTcnxB3GDUel7fWJ2U60PXOlmY5Y1aIUET4uQeZMsmOSzjGSWFAYjaI7QpE4z4lGq1z0bZX264F
u+6etjQnjIsm/nOAlMk1lH2b1H5UhERXYXdgpNk/XTNWpRk6KO/JiUhCLWFityo5hSUeEWzLbq9k
rrSFloHQWMZThGMn0+K1rnO/7dmf8OKt3XdBs1wuY/lihLtURpPoXGcLtxr0OmSYGRj/0uAdTwPt
BTQOR3r8AI7Sr+vQp/LQgbjIQVU+GMBfpJKrJoYEfo0Dz8D9p21fmZNURLpU9eXkb4BLNE/uwxWL
QiTmEEXC9tqiCSgy8ielbiqjuOB7i1U501iNWi/d+Seka4SoK5fu+0uPbwcwwYoU04axIZuXZ8aY
BCBs5CDYGaIf77dhOHC4KY9L93sRECmcUkjYYe0AMcQiMeJppiqo/DcTcaZtiZxoHDAI58TfsOhC
h2FzE8q5N8Zgbj86zZfP4zDYNO5p9gVTg1+/BYv9msfyWmKwqyRNVNW9dkI9WMWYSRjiMNwLBrsJ
bUpd7eZgr0fkiffs4enhJOqYSjeiSRwnhBGYTDeZOvWB6OQK6Gko5qOsc2/DDl0mzDYhtB6FMA5R
CxCaTGNiskKKt4kBLgb5YWL3UAlsLxv321XUh/fA1+dWDDTvnJvrPllw7g3d27dDQurxPazXil4c
Cv4EhQuTAUGwJlevEyocXuNrLcYbvxt9NnDS9hnlXCugIOS9qltvcg1gEKK+X/oBJYud9xcKf3KS
X9bkzTGqftf+Abc3Q0jufoVjvBd40d41ccApS1k4gF7LRRj4sQXUR3m2g9Hx6gzZ82Qm5j5kPwyI
vhjA/cXK1v/MLlDGjYOhwndYOBKFPCc2xwO/Uuc0NgDURo67X0VibZxAoCQfckVoW90BGrZ1ji2d
axQav/dIu6fXLZh6SEIkYnSLMJulENarZV+E3lba67tmiu+BUNHeUu5ykGY9iLjXj78vYrzlj08c
yzuGVZGyyUSlai0n8qWi4F8FOO091FARhKqmWIiiGfV+J3Od8E+MZZm276DYvJPP8/0PZYFR9dRY
WQR5xITdZ1RVpzB2Jd8ZONUfegslEkrxQrMKthr/MJm3jsvxluCnNS/6G0Fyn236fLyyL5x+8ZFI
uk2ts3XYQYMTrFoRn0HvlFBJ8q6uc53l+xGMF61NJv+58qnkyUjex/3LyCOYWqNC41JIqm4TQ1fz
b4vIstykJULmixm3mIyDaiazB4G//F7s9VK58lLx08pReGCBjiDbV2oI60kNc8gYTiOCpWVDtxKn
NPpZeRpaCyOLmToCEsQP9w0Kw2sldDtrICJIoNkRGJ055hCxv7LaVQuGTdacQ6/4aYM5WJeNt2zJ
ivzWXdxjprNB5+mprmT5c0WtMHt0CWv04W2Rh3fImrZbOmMxKWgj1pzUR1RJ2GfoWqKPhAurgug7
nppP89nxhpCVl0VJE+TNQDxvYvVpFeSTqkf+BsLA0oUNLDqUJGE0wZVmNBCu4AQvzRn3obI7doS3
1PJVSQ9dGmz2Rp393rFHdhUfnRcOF4aNBkSlSk3IhdOBdKEpTmRbKEDkN2F/qVUofcDLH0btQdOA
phHp9OPtUPpaYt7ev5j+hZUS4XRoBrBOsqV9jaJTo3hiVlPALkXdsaExXcxr+nyFPixLRmm+taXK
NCOrbvIIQ3IcJ6RvxHB9MxiXHXDjmBuoJgaFnOiMBWaxGG8V8BuaUM19u+F691IDKCqOim97G0Iy
PhcacLqqJQ6anQvqP/PxhLOebqG/6A03Tm7frdkRfjCzOLta7W0DU3EDTfNxscboTo9UNXNme++X
QfcJfBJV5VPiAgO91fFbUFheUiy+g2Ly+DO7ZmguGbuYrFgikveEqANwXRbwjq4ZCRpvLXNBzFXl
P1euqZJJSTx/AqjaQ8D51At5V0gLRCFZsgSEPuLeJYWiSzsxUqnWpsj59muoEUi/XRs4N2zz7nvX
Pt58BbPwCdzKzw0NsnQk6Vc4ve33IG224mraSceXGYwl1KDVKRTcD+KBQJNBnwWo5MCbEOtV/+My
r3nnDtH53VENt7AhB9CtCQH2A9gM4BYEtnn6+4Ok3vChLuZzEmZP1Ts+/uv+okakAGzGdE4fd0k2
cUD3Ql2BH8iVEwn98ZANYiV7JxVX8TMAHSGqnEaftLzljrtISKBg6t64DFGyPrS0AvEY6YwjH/TD
6KY2Q5Y1oaiBTTjYw4An3ZnSSPb4pPLIHb97yB37m8p4mELpQEGFU7xftuBDJEA+rC9Tlv57L9RM
XHNvLY0i53yRCuoVMY93nE+vlfwA7UB4Uk6N6ErwlK/ZO3JwvMDQDqbB5xpdLuoGZSyB8Kr67je+
wdK67v8LlA1lFEzgmyestQQAwqVfoNCMdbWYuf1m14s5Xuxb1imWsOq1397A74aKIKHjWa5O7JFV
u1/did0MvteFYVqz0e4B3PSpp3DUGGC3vvkwLlHuhg+b3t7jFEjt8j0RyFQLVVBkIEXFf4KPuVKE
NuGqDD9VLr2medfbNK/ye0ZS8kbkOQljdj+S0zHHNWu4aD2+PEv4C23e+vZnCI/KR6QEBwdLocpt
+CWtyBSW6zuKFnie1PuJj5CRDbyYHlfaZPGi7EpCvuoycuG/RbmZEHepfa86Z4xNFdteKCL6fiq+
8jftfJH/Ymq9W9RSado1NPnOG1WjzIkQxTbbmA6h00d6VOjYQeRjGbAbOsPh8tkPIFKSp76YKQ8C
M4gzwe/IoPPbxKh9U2c+VMsutWnpJRf+2qERwk7WRdfc/CLMUJUg0GdtGkfFJoir4cyfI8tqbhP5
qtKlBZFxtcvThbuZWO1Ew7v7Ol4OHPGIAI2+iz3mzH3OCxmiV01MIBHC02sOxBZa/V5c7SNkLmzy
AMv7K/U5lnm6k70vhKlbvf0TjIbPGin16Uks/hEEkss0KEO3knU1Yx5/6qx5L9ovoAKNBnoSUnEY
21lTBuIs9sPXr+2cY93VS4j3zvRiU7yhAsidY3uPm9syipr6aYAA3fCO22cpV9h0iEYWFIWJfzz3
sF/svlI9S9kmCs+mNPYya3WV4g90+qcQWAlkc0tB7NKa0R1uPehdAOhY5jmy8Wj1lxLmo/Dv0psn
nZotPHFCl7OLoOfyu36yYbaZ/G8aVObf95CnJ+j1JbJIauGCJ8jyMM72/GHvp7qOxaP8IbkNRlZq
mKKtwTZa1JwQVtetrnSDnQGfuq1hD3n+uESdXssya5k53Wc4Uoq7jGQOSXJZ2WoSMdRCLD8JMsXJ
HTgpSx4Yg/E1TjvvLuoKfGboC5HqibvF6GCkD+9xl70LbpIQHBk4PYP8RzcPnFWa1NckkK/O6esM
5WgcKNwPgXyi3xj4YaCGGVNY9EPZiBF3c5n1XElPHxrw3b2Xw8dZg9qbLcQJV6POLk3Xpu4GFZpf
FK7SogLhQnD8jz29ucgfy8D0pU83wQsIG8lXspYt0TVnuB4rOieLVQAOw05dGceJhnao288e+bIG
bZHJ1GMm1anliW6+2rvFqfwJbl//xbufaNO8yINP1iYOuX0phBTRrmswXrzgzbOKM42C5BHv7SW/
Rtk91HOKvdYa17nZ5Y3AMoA1brKyvQ8zgW69bY+CIscvOIZMrZ9voZf/3/5zroq3atrOGtpJ7cDq
4oK3sU4PEAjcfXd6y562Q4JInR5+T8a0l3bPZChot0f4MXGh9LayapkoY4KKcsEKsb4/Qbqyw5zh
IODG7E3JcfJF1fLhNAM6vi9LUR7YuHOmDOh3OkZ0A8BAM628EU0al/zl7FMZGfCkY4bVsSEw5Gco
uP49EK2H5z5362qcxCllcjC9bLCvd2n7Hm3qjF1YdQc9nCekmKjq6vUOzR9364a9tpLODRNPwp/Z
hRIqApPCexfqIW9fi5OQEZPmUxNC1FuQMPIsUHYFxtlhnWEVu65Pe0JGy5T63cNLDVccgBScmkGM
VO1Z7Xm2IZvh3z1azv9nrmhGmYOWnt4urPP1J+07PPluCD78hwxXJ4ide64M1C1XH/VoFnlbFdPz
MRY28vZoMy1sEQBUb3CB4Z/tflHD86wFWXb813DtLkmbWraJxGGhsqL0eCTBbSeUbUnRMPuYAGDP
IzQUcUk3IHhart4BMi92tg8LAbUg5hemik3LfWrR2PMBhHR9APGLHaOxxMU3MqB6r6qvE/NIRjMd
DxYUEb/YtVM1alrMK9b7KncJEKumE+M+vzeFbw6/zGVZd5z3N0mHQ1WPoipsZje5/H1OFpy4gclI
aI/oQ25Ne4abChJR169WSC3lJuaojkMc94Du1wh5GJ8GttCLOtWvURyui2RFdZQSxFQVpAAHCFfd
6Ft+sG6AnuzSvg7KlJfUJ+DYPnQPMp0U/xJ8AnDbw2uSvHXwPLws0l8czSVL1hyt6R5UscFp+Uij
0gt4+ip/TQNj83QFptl+GEn5INcqn8j35yToQ4w4V47B7YfH4WJOsXQkUsj3Nqd56VaRts1PzFFX
mhmIE6Ea3ffKik3DjJnvmHKF1tk9Lt9TEF9vpgvtFTw0GHWOMf+A0hWuUI8T1nvFBgvQJ9SJop5H
k+BB/ATmnJRj5unpPYYq0SG7EuDxYKTmnWAJSta3KQdqRrOtCu2ezmPMe8/4ahUa+nzbZAjTwjX3
fGzCATZnojEiYsUov3c69dTK1xh83VxfoDCle+giCNNiOFdiTgb8tqoIFN6iNGgHQy+ZTPnYVAy5
DFmGEOvhO5VBNOPpH7ktSDfqJ4JFbSkCifhlXBX7/Q5pik1I0brnlRDMwsmj6q0KJ0XsDvRaEEj2
8tCvPFNauFIGN7/OfVIseqCA3kG5EZrb8vvol5EXANeTlEp5b5/iroe8sOdVokyaATN/5Q8Tr9JC
p/7AhdOTJO3FZd97uP3ZPKt3Fo5hUZGBIOA/vp3eGNFoq/R1rF6b14DIr13wXsr5dSv5sTbvAWto
QmoU2qgGZMZTB9p9Q5JGb/bNxWzue8OAZq1eiXlFIdnNxeA5dqcQ/KXQQzE8mMY66bXG1JbJcYTX
ko/5Ple3gcNOlGmFAlkKM2qy/2jPx1Ki2/KnyIEotCAA9t9zqQZqGj7nJUQ4l+T0dpPd/xw2UAQC
WVaUGG9hB2LQoNERvQ3R9gsYaGfYddbfZWr0pl0SzNgqRVCNnwwyQqiip8U2pCUGWy6ZO0d/trJ/
p82WqQ+sFr+Q55Fgn2+tnrU27xwUqaXcpmqiuU6ZyVCKALq5uJ6Y3JfC3nIq/X1jfb6JE0tppl61
5+mHBd0XMEevA68pLataDI5x7ByD4YCDaNDv33bYDH9ubGokx96dHOj2w4m8QSb+Vg9HHH+jeqr1
fcpamOYNyzfz6zuBBwfBuyPNMlFnGiVnpwI9g7oJ05bNHyVFdKcQT7G7uPV1aLCFKQij9R50J5N8
3QoMuqrphjeX4BLMmAEIYQ6r7NY4HC5zzJ4sIkLAFjhPb5QSev78wSZZwY9YOdR4zuG5Pbn25YMT
diBAIDMIT4RiucIXq79f26qgrnB4oXCg+/rhCr3PEivNSPaqOfBHC5dPeM7tPyUc9h5f9QB1YAbi
PeTbc8ZmmvcvNU2q7vGjulRdjzl80kbwUc8o+q2IxsXmTAhXW9ku5XJmWYy4HGM6NSjAzoJ/XFe7
fa8VnTwk+YQVe58S0vjQ4I3nBPANxrL2HON8r6vF7HqFqMTJqI0f1gqLRv4X1n+nXvqcEzccvZVh
/Rd5dX25T5JpoBbWv9nFlq1OXIHv2861MAHOe1SflwKzYWy5JP8pjZJm3yPWR4zGrFAWr72faA3o
UgTF+oQlp+HvmkbQ3jxjMkg0J+etho+puib4PE8BsAf+INPIoGYqv5M3AVypPcYyL4jvKR5dUMTS
oHxkOSgOPK+pidtbBBXyRQpdGBykRqEO3MSRobgWx4AIGUMDjOqo+6OHfBaSD5sX4daxBl0QMMsi
VyCdgBJ/MDzuA0xWL4ujA4eyGB8UN8HzIaN7c3YKYpteV47PtgfpV23sZdLKwRpGevfEd05qg+yk
Ex41YSlQv/OKS6oT+kdGACTmy7JMfP/0qHk1HwYhmzXrtFT95zpE3c53t5KDqJrATcOvgzCQOhNZ
4SX0v7GRfsI0O59K1CxBGufTAAFgNurTHxgqfEvac8ku1H4cJrHsGNfMoKo+0zlS++qv87PYza5g
oygGu8uWWu63nlZkvMz12lAA5x7Pb9xeVZ9nfUBEw5/nKr4p4ab5BU7thNcli7Tz5kWOVB/lNcuH
FHRpYWD1UDKKKFeRdFR6iR17ZAwMoa8QyGOuOEMl3QAoedJVjb88sZXs+/Y0hL8CDYol2fBkh+Er
NNaKLuMfREAE+vUOiCEGBjp4oqNmPtRDpaT4099wjYEQRiY72vCBLqZw/8cWprG9JA/HY0h0mXw2
iRyBf3LfOGU3/qeiW411msGrOeCuqk3kdnsmAMDw7VahkU7/yFP2WJ93yiAAQaYNunZCqT7TdXdG
tv9pM3Oagpm1+UCdatd7qFpffuMowQLzpKvoYIuDpih1qJdcdct2hMR/NJoYSMkG8Vw2RZPD9Pbp
ujSgpepguHFcx+cAJstk5gKD4AScor0C16UqbdWjMcrzHUUg8ATn4FzGGZrXe/BZaG4OE0ujS+oY
YpRcOI95pzqnn1pZNRFaBx5mOw+ik9GrMTPeBLyptzyVpvhVa1hML3WlqNRKDTteQlE3tpAHs0sY
XHzBD3RH54U6opLzW6spDKdPmP0c5eWKTtBw109OWVst/FnXb/zce1rkgLZiuq/AmWHa6IV9SVTy
iD9DyAnKC0+kzRyx8b6J0UJZ1T4ccaud+OdDlnew/ISIEagjevjHQwRU00zMCKViP7j0uupy5kzq
euAhtKFbpzrAMJqJfr/nHL3cWgPJRKrox4pHEZE8A7I3vOLMuwtWKUOLYEwVB0CU8NftPYWX6loO
esn74x0pWg3hGzHU5JKN4x8hgxRBZ04YhYCpZz+C8LAgKFF/p+zBpDqI1tU+wgK4X06nQsxaSuxa
qNyLBmEwOgpMgDSnJ7rtbTJYOr1lYnC/gU1Qpvh+5iVng3BuhY1G65TlN4pMpVCpx6tI1U+X5Mw2
zqAgxZ79uEM5D/ESjE5npKtnoNMYN8vY/iM0zPmQPg9Kd01b56v3srKiahAu4fb+VCBKowIWCoyL
j28QhjjmWSmcN3Z82okgg5NrlIaIun4C9R0mg3UXmtnVsEQHosQ4VKyPiry5vpPLrchIxo4HExam
4uV2+CgAeukdLZG+dh/2L0IatXooYBoHImHbznfWo7+PlujtaH0KK7B8JLFSazcw8cDNTS3B65bZ
jb0+lu16duxMlRFKExtfHxK2Tl+F3kH/phEBI/prT/UJUA9QWGd3wJ/63npfzb3XoSM5+pe7CvEp
08xoC4Xur9gBLkqYbXkGgtkXhOSFBh7WpnwlmOxvNWVgNacVfUMtTp8GKw2TDr5C5Js/xm7FTidt
mZpAQkXs33a+AwFSL/7aod/adbLofml/NfFkVfkTgzLuMHiP+c4C1It3LJpv4XQfxKXd9vWR9e2Y
CmGZEXw9Qpl6Soeg4quAVLXxDTf83MdE4jhxc7JH5UrWdbk9+vYkdjjJygdOZPuezrdThu/FVuux
dgspFaA21pUEgOPthb32KiqaAVuh3a2pANASecgr5mLk9L7HgjeaStwpig9BPyOh+clbD3pLE45m
6DseHpjIXukqa9U559vKNujyl4JGvHiAThfLuv2StJ+MieZXsnWaaHz3FficQoHpBXHDJIZBNu9k
eN5wdp8UYsHR7AwuKmf/kiumtsepTEtyWBP5/m5QmT7dMbvSdM53iL4vWBbSxrDyeEb6sZ5X8h90
o0q/2Kcz/F/rDJPeb7mQrG0XhAWVZ10zbV80zcevWSFltdJw/62eTpIZlWe74cmDfUU5SxgzKiSf
ioSDalO3W33I45ygM0jfoggicFNf1MKrwusZ593REhLnkdnky0gXWc+EkeOA3PkOzZMv5etc9FMx
RCl+TXxhRQw0qJbQNPJg+Hm20DJz0xu9+8bfDm2+EAGvGAqyBBuUpf14ZOG2kyL+M/X3MVFxiS2O
LYTzzmRkjX1LjZkILjInGg6d+dNnjouSlVgSd9QCQnvezalDeHgxiS6mK6ijtXK89sMKUuL84Mm+
3Xh87lUhAaIqsIVeXEvy0iVBnvGiDqwuYuBm2VZzFm754uwOEwVuWhfWXkfbE4FrpM5+r2KIxXWy
miCe7uIubmvJqj6hogWn025/Iypd9jI/st+lvMOm5/gT0T3KU0yTgZb0MRJHA9zTK6hcTurCN6fK
+PjM7Nxka7kQQA/R/qdv5QDjdUXTJnJwj8imST51U5tPSTO9wDlzQH+C2kp6U/1IhuV96Z5tjxCl
LZbkQ+pi+zpp+AtHK0ZvNoX+tr3wf0byV/vhhG2czawmvqlHDN2IQxrp0olV4HBmlZQNlEjSyer6
DgdopsV/30CXEq8GDAD3SviBxbEn73nUNjzFxL0AMfMZxeAi/+Orp7OAw/YoJcCI7Ahy6Vx6CBnJ
8GQQEfLlZYuJchzmmQ3XNxIs9LX5yjfcGo4C3WcyMqLZ3xUB59FVvkdpb76EP9d2jjSCMRYrVB4+
rYoIsDdYs/KhOZpfPSWfvAL993KeUX4f+qIfcxs5dFGGsa6Bs5rczpjX036i5uhFe9RAyaBMA6wM
rMhZh8XSBwxzy914zDmq0M6g/MHlriUOpglPK83YI3YMqxNoJXilusXhvl1DaZUPEeIi0HFLhGJd
tigYKdPW/p2beyBtC5QdzI1I/WCGCzbnFgPdEya84mCL+Rj2Eaby5mrhz6Sj/cpDEMclFXDHl8IF
HjRzh6pL9/F2aXtOHehXBRrmAxLXibtk2BNPKA86TDMzqIiiew497t7ONlFFHHkilFvNDllh/w04
iLH+HMQJN9l0KR1CffUimbh5KlTNF0Yu1ZqsFaA2rGgZqmzpojXHYWOCYCuboehCw04SqtbcZ+O9
9YplB85wYvR/9pdnpUBggDCgbMfsih9JzD4DVH6YdMdeOoey5/8ez4Iv3g2BYhAhIIfECN6EC94P
jPJQgROxPLhWwODyO877RZgvtZc017av+BbVNaq8YpNXAnPdJv8Z1CErAUascoAluwftAATzDOby
f9FE5dTlEMKIrIgd67ZIdJOJxI/p5aDCQ5YGpNjKRHRqi/nTOo1vEUBfyFKJZWOOAAgoYqevu7sO
+5cGGQMCocIsnLze9a4IMgbxWY37SBYCrj1LORFHxk/RStI06AwQiu9Y4XMCx3Yql+4IvYJRwnTq
Dq23DwFuoescg418cYIQw8CTwRhn6SC+6CU/U8KRIMrfEJtqDCHgpVpMd/E2wA+ohHsuNq+ttcC5
/MCeQaF7OMs9czMb/InmnoenLtX7AvMvgZWwpyBNWJbmABrJp05ip+UE9/tiEd9zj3gbbK4ijtL1
pn0DpiAVA3YRfbWuvV786MU2ndj0UE9Ja9EJWkvsmR8CsTNRNayfZR4vtrvxaa2o9IkqxVUX6XrS
7O+U981GVcxMi1x5bn2deOdK+e4bZJXM8Iy9jJNvTRpzgObTuzo+h+iFujZfHoXXxwDfiaccy/Ns
OSoHJIrYVLfqWDTqGSlk/jc9R+9sCyXaXG9XMqTQX26cjENn5dU/oZsNvL9silIMdEgGexEnlYOZ
IMIcSF5TeE3cYoMqtF03imt0tQc5ppaLtj2WAJsOpNehh2P+vWCQo+Wiw2vv5+yaIss8LnsZGsf6
cyT7PoIth/iGGaaJIjUV5BuTONS9azHkXIfufPeRowCeJhZj5aFBLmTJmVBpFvYir2SVsiVCoBTs
IZWsdkZLPVLD3QJHc6qZFEsDWq5B7C0F9cdAb6hb96q0qv2W9Z99ZvpUkfmiILlmH9oEnrjgITYL
AMItHf+1PzvgXYwbIaxda6XkSB7naDXvcRGCaNf7qVY0kXdoE2MsPM+BxlqzvOJXKfAM3EIyR59m
49U3lPEK+D2DeNKojwPO6rq2nACHtpuAcOA9SZsF99U7eb4aCC6Lq0QM3pF9YtmeGPt1Gca7Ft10
PFxJUV8aQE1N6XyMWHrjswVzD4NkqyeQSUcO0by/khy0vE55cZjuaXuh4iuqI+Ks3HdF28ckNrcb
TRH8e6n1pwdb+srjb88SsPpqTyFwVSgwZTpkqTSyjZkHJt4EKz3pSAmsywlJyk5iBtKxG28tA8S6
R4wdcnK/ermr0f44QHuqkwkfutwU1SZSFYyUD2G8w7zO9gyHHkFCAwZ/+e//oO2Dssg+PTmjH0K8
4zRcM/3qxOUo8Xm34iClTLxUrVEAJMwm/OCRETwsHKDEjjxnHNVYnPTbE9iTkGPRE+Pwe+rybzN0
3hAA+krUWSoCTUVXFO/9k55PeTMVsfUia601wjRNfmhVMf8+gzez/dV0KDz0OX2AYnfII4f6QKvM
LKeTJxxsPojHd/zmTj5ESM6hLTpnrXKNDSMO/mnJX4b1Tz+jutV7+wSkBRttc1EQqEc19XO10+EE
6lI5V7Qrjzs87vp7PLgNIwatdZrprTV1i5aLPpseD/bIKMuZ7vSjlwTZrCDHzXKwTCfv6snfA4Fs
uuIwT5Xc8DnOWjZrBdZSAbo1v1AcdYcJmfj2ROjZ5JICbPRl/tC7L9pCT3F7hjJg4TR3SOsfgG9K
XrhVMqvBtyCk/UOs9elQlXPoKPh+SnYA8PfJq84vfEsdjo6Z22EBbg38pGHgNtoneCP8cIVfGz+I
zohD5vY5xrkXT0eRqkH4JeHG4VZjpEsTIAxirCLDHULYYewEY3dWd6YrPSWmJ4mokySXshhiel67
Kv+0VUfAMM+zj0hMGUtugs3St0nHvIxZh3iMUwEnnJvlvAgQpAorFeM1aEbCGMEqllKay4hXo8ro
4OxhY2epOWIwtGBguLsBAHdulz2/aj4NcQoYzAhcW34SaO+8kWzceHE7s+dH4B5M2Irp/yOEm1qT
gKEFyUn1MIDGnl5in5ZHYdqnLaZ2bHGmbYyTAmbw+Xs7trYqeV/gzt8RvfnHGWfnhxYQJN6Cyn7V
1AOLWdMzVAOV4VTUUeX6QBdUDDcyciH71rJyMTinpgNbLTMegB/cg2eeheTWMUE4W7jpqi2qdFTu
bKO3SD8ukKtI9gR+oaeFC4HjkxP/LhBxZUhY8Spl+h/C8ry8fQHx1Nk186rYtry7SaF6mC22RqC8
Nu6FGexPSAQFMvhiFvaMHgRKj+Y75Y3I/3vITJKVF7SMo6Eo70ve41aOZKrEeJT7bGE4ZBLdziOW
eUDAzxkO1Gq7fzvg5DqwjupVfoYJcqUj8rCFuTE1AqRG5nut6rCO+OMqogaZ8gZ/ziPvbWHWH13e
X/ajzkamuSYquOpjKAa7Kb7SWB5tr8mQeXH6d7byleApfCrrk2dQHSSHH50bpZ14WDtBa08vYyUm
8YYzQ+ew1SLDCmaIYL2kKqn5aw1hh/e7MymBYXxxze+XTlqLcw1BGhXa3Av4IXA6C+7jMczNV902
Uzf5ahcK7+GYpPjGkRbCY0a5+xaqfxFkwsfmMzxyxUaoJBMHUJg/tgLpxoFpE+hzedBGkbdm/J4v
8Y3Rz/JQ5zlqMzAXjcA5P9YLT6tH2sanun14ivLXwX0hAv68QW9/hXZHT0YJd8CYoCer2mZcdtWu
1S2CprmDFHv8LcUhiwZJJC0D7wtGdXTUz+c0q57mG/YoXvTHgeR/tExWKR0eR9ZUv1KlYVIvwD2P
gKIK9rWFuU7JNA3v/PeaSFgAVobj1oaq/aT+Tf6SeF139BAEysNkEDIWEBIQEJ9MMalDg7BDNvho
mHTYAsWhD+ARXKMgNOX5npyYcOzRz+JA8+XUFdi/nTzZ/zp6ALdcAeUeAsChXr4WW4Ianc8FgSQb
rEdXUWfhf3a91M0TP08eu1CyGjvZEQXXOantT1pMg+5C9X4ZuZwetrEOe8XxTLbpTKWod0RkDhh3
K0Lfv+gsXQ9GqYRAV2TgT2mokOOJtPLVzufsW2CIdJyG0plyXDDaOLw4iz7Nw/bxITVH0N8KOkZc
fgk/ARB4e2qed1ouzgMXyt16Q0ms+ABDZNRKc7Z7lsC+6FBdXdNNQrt7e1du1oTVRuJMzGXC6MLu
3QbeqBYd0WKVDwFpepvjyd3RJezBAvuZywJmuHJGAQFxNSrGJJsuXQQ5mfH8smeeJwz+xqeD1VyO
//8Ds3C7I2VzbuFSuCfWCStc7xjbCBagedR7+xnpt8SNC36ZCP4VTaXK/X8VshIgKwfyJ4GFwu0B
UKuBieB6UXeuc+uTXltXlw1tqZO0cSmzi22I8VbZ5g4shN/NyS4vsuybD1g2+MRrDnHB8nmHIftU
p0bJY5Ri/vfmqrVKHpfL80BnISZMB34EFc7OPK4x/OfK85EDSxmDNVTx+VdwvfUI54q9WsLswkad
58yc/U/qi94IyG7HoJUw22iTvpNqc06fiwn0W8UDmoAlZHQ++tCfzJmcuXX0s7R2xxsyzxv/BIws
Nsodo+YnFFJC71H66kdDNX/4abu0gG4tFiq9DYgehyhKOGKi08U0gXVtkmi2KQhTyng2Shuj7WT+
4lG3Fd8LcPVgI3qSKywd/0IR/rgEb8U0RRD3re5mmQE6QgzdNXJpAMQrPh8NYVhhE01ZL+JzJomq
5g5thUWbYmHaQWszJL1wlXOQT8gez9/EPAdozuM4yydFrxJ+wpQHM+YeGKIyeevv+rGqBjN2C0ec
J1wJC+wq0L2vaHEU1LMrnWN2JW2JY8iu+uLpjG4BUmm75Q/BC71yHIH56BgPMGrYBdUcJt2dD2Z7
lL3eTJvBp9oaQQkFKNSmBIOuPQyv3wpLrYuCGqjJxHM55gf1BLujk7Yx90HRtWjR7tNuCNncnwYV
lqJonZngoeFDPt3UNwGbn8V9m//o51gIpxwfpKHrNFd4LiW3gv6AfZYJATr4atqnbgGKEnqsklPM
AWWRAliPeWukyVoZFC2+BAhM0t8pY3E5tE9k5V/8DBOSvf+iHodQxeFzz5TD231kv2ycyzFA32ih
QTIaN5ewOJwCnpz3W+0xAKT3t/rV3/aIqaMSzs/E70xZjtj8oeEo8/aHGCAF5NQLPqaSCNbMhQoM
l1tdf0ag3QzNzKl3xCdi+RObUaajEzlVrxngFNAmq1I0/yivYIuUd6+DAIdzPboS6nfyomzA28LD
disWBZy0JNABoIiinL511T3KRnyZtHCv3EnCKryrYnaJkuOD1+6aYU3PjbtMTfrKN/EanWEvpTQ0
XGNPer3OtTbzbmO8srY1Jwm7WTJETvfeJ8PjeJ67UQyy2GHrFn/Mktsa3Rp3spk1LEkFi+z4zLAR
rrsMmbMEO6Wi8wN+3PZxIlv8U2nf8YBw/tDNDU6acYE+zfZpyK9IeucTdo6AtZVNr9/pNQYGmQnN
BEUD4UBL2Syda9z8FOEOUl6eZcBMRPpcfL4ArIcIdn2fVj5mKns3zHm2GPEHXzuYNZ6xLVStrbDc
fWepuX0VB/zweGRxTj8290uIohpSfNeliByvzIMwxnu5QdbtFk+kFpNTlZPJ+zBVhQE+gXWXIE3V
4pv4j1E2x4WIhuu2n8oHgo8Csa6a5rbiHoRy7DzaL5f4PsbH8xqDhuOhFO2Qe2zWQ9kN8oci5pfR
N7HoOw2A9Suf6LuA0C5rsOTpxtC64kGFgBiF+Dc/R3S0dyafkqnb38LRoTOlzQ4U0JtsV5RTE8QK
jQkeD6yDSvH4l4Cx/B9aJxrRQuJVAP96ym4uK4v4qZiRd4Li2kAVNsVLPH3w6p2+E0uihL/4Kxnq
3BuAGnQ0lOZrxsPOjW4+Fa+iG/coTpVdbMW/4FcXKn/GIX/tIhk7dXl62fCfMj+5PEC3Lsdnt+ZH
VkCZhPmIr+dVlhJpePZCxIrHe9VfDunmIxA/MUSF3sXOb94WJKVQmp/HKzto5WYxcCHS2eSqCFfX
e+oIyhxIBjWy30UPNc2wtUawSlE+f+qDAoSbHrZByYkmfFLU4HfhPG5wNj9rVV3fqAIiYagd/cYS
L6SgSBrt9p165raSNSIv5mNW9hCIql4ophoJuuSlMcC0cV6Ob1LPaHGFcJYdVnEEzvxqGxx5m3Uv
rtCdl3ELPkO46ZIROho7YK6nXJpwmrtdk1guWJ0wyTxXvTCPyKiDMk7bRgC/IF3cq7vW6D8zUTPh
raDAzIK7XHL9UGLaxERrkydf6N2ImwqabI356b+L5hG6qOJc+aDKh4Ie6Of24R/qUBIRv5hjOKJS
3PdZj+8/FqPAhdSx16P+s0aEFVvCP4V89TEhQUdeVFFADqfNo6pjoNb3uHbnUX/ZPgmLBMz4LfZr
jBPlLvucw/tuZYd9vJjs2jk2VIL8HnqvI46kYsygNldzqxUhSir0F6nWrF1w6hAoxNTkuO/AUtUj
LMHN8iR/UwUv0D1G+0vKAYFn0pVolADsPE+8kHClT7DeplvkLcsrjeIC3F3GYm1QmXImgenFUOx4
wTCKMFMSoWnAy5JaS5THArAl8KHva/odQLj0OJuDlI+N5MeRoBo4k+j4f7KzjvVl2dyePiHty9J3
szHCB1fV2herikjotEJ1NQbmguLhKmh6U3rvwAE+3cCy9u03yor65wGznOtcgCyyhu/G7WrCbwst
Eh/TbOruuWAk7vkviQGjXRJF3xfnwNttvKKZ6t1hUL3Lb5Fifvyy7YOg7vBUOGKpEdCvnEUQlm7f
+QKbaDbIXOLU+Xw6liJ7F45oMr5BWjbg1lS4yz7HghccQ1RR/YaUGvBP7+m+KysD70+BwjljZxBv
IYijMFOvAGcvTsqSb/Vl5rRUTjigwDniSvSLzUMgBghJh8MLyG1dHHoKDAXE7ZppquqLna2m0UyO
dEyukbqk1X0J4oMhRtiQC1cOPk3zFAgY0UxhdwfPQgkP6jR0qKConRswDeKGW8oaTcu96Smvxve5
YkFYrcQx8MHbVKyGv4k00Voiuynw2X772gKMnjzpKv1g/3S3B8Bj8On7vKoiO7cMxupUVbwwNaar
xIsZgGksqDYcfpIfFsK8WU7kjPjVJewJxuXJcjAfBVsB4J8ZuQQsl75gzDNqoDb7Cpp50+nQGK5q
q6WA3Fvd5IwaSbsRTcasPxajWpQqgTgRh5ip72PX/wr30DEVxmsXSr1uQTi27AaEwkrdwOojr9wM
j5toYrQvpEMZSTmk5nJqrTyJ4TKglGAA2e3mKatjeOW6vRUT79fIC4G1C3ZPJIr8+o6Hdnlfr7tY
4G7TmSoS+NGVI/YpWx8w5mlLDc6o8AFHWO6KwIrzabTtfgSb+TA8ceVpYHG71UxFLAqi6ex/Z0ld
YIKcSRIwt44Rjx8ZrYYJ+91Xyk787XBixeQjKdMvivu/0sWfE61yUv1/ZbyRYg+h1PEqXo/EsBFp
t0YmbW1lORM4KmGq/c2vF4k1kFvRQ8yEEtGGbxMw9t/+99gq+LgwPJgSS98w1kbxW7uo8F7c95XJ
ZleFxxxuzGVSCLYHJGtuF9CeDI1Mvk7IgfkcmL4N8PztyWqarrmkhDTb/YKfGwOLvMN/uazXwA9W
MetlCQRawZINpzFaenowLK+fOb8uiZPy30VIr6aYQ8tAnkKcOYtV8yxJV3S+EI2dZRyiymCXXac+
goIgqCDLKv16XK2WY0SbFIte1/5KzTWQsb+5QXRuE5TmL/Dao6ThPcNX/sRdwogaTZQSg9gqrWLi
nvfG4wIdhW56QQMxmgzMOuAwud0tUvVfxJ41qHKQpxk5BGowvzvk+WZTQ2H/9Xmo5MIaa1wUqWM/
k8dR4TF7QG9VoSDGe6uUqLo1gDNs3zA/jcfXmYg39mdJKQ5mfqhi9lIj/jfb7mZ4xOHOGDhrHb32
CU4cjZ0sZVIKv0v1L50XhYGutly/VwXPElAOONrEsjAq9MWoom0SZLFbIE49RpHwKPRFACmCaL+s
HoIfi44YQ7qWMqTedzAfYNPru9j12f5kWTbocKjjt6R4A4kJWlaLDSHcqH2eL7vlrmwS1sp7+syP
AwV7b/b2LSNtSWGRkdmhdwVcwnvdv2tbL51HNu0cU/nvpR01qXKUsEf9DpzIHk5gpcIsMzA11krm
lL8AUKW3LWzzeIh0NNIOYh962XGcvMdATaQU489519TiWhwMoN62dhaboob6BVSxKqpJjam9l7f8
UiyXRvf6NPiHGPncPI9nU9xZnMWcOqfUiyR/zsRiSX7uLIc/s7B7bco3zRtMcHcVaisfqRbP8I6F
PkFT7c1EAAhXwkeyoJVo63/ScTmwrmb73ZiHFgTDb+AT6vZKV3i8z4gLfhMhc+dGNadc5sQZu4+H
+7sDqLkI+itHvUZjAKadbVE/MOSViSEOKf1Wwku4+SiWXChIHFKLaXemT94TuW+0Bj2KxSUMufxW
SwwHIaxvwC4S/5bgmx/qIWOsbCW6zR+yxiir3+HUVkeEf7TJrbumrCSGA5i0UutZURjM9q25khjO
/T4u8zXwFTk6P93AA85Mq4PJlgw+CKECc03FLXkBqSDNriBzg4yFmeADdv3jl9zCmdCWjn761tcl
4vSQOW37uj+W1TzoEGxHrUoQvv0E2UMF8wpqCImFO8Cvsc9u2NcfmoHOcvwZAYBVwGWcwlioRXkm
mD/KiPW+BcDYdy9Gs/Mv268DZIsGG9zl45RfctxeOqrcDYyoM8mBuQQdotrzK+KIWd+oJ185jTjX
RGPpawm93Y+n9GdvXUKEGBbLv/4FfC8JPuPu5LH3Cw4PLKXTBY80gmx6ZPaGUBQavOwJCQr/Ayc3
ENKshrPwdPSKx3lunmaijHJPiENPsB+UBoay3JCEIYKNzReQ7NgdM95frLUhr0Y5foIUDakeJn8Z
czekhr5/Qnl476rVuUVGX+U5SA+2+F7cMblezUFRi3sljRjMzg3URoVp+EvDOQBsYZvnclV1Bb2J
un5k7sEdeUjh7hDZ7zz3+caOC17vsw1bzut45vZsZHz/BpzC2V+SyOeFeryFUuAvIkIqbJ5yXtHI
mtH56tr1v5cEXdXcE9Mnd1bhSPNtEmOz71aU36WpZ31+i0UQHJkIActN+LpU26hKTG+VwmziPqrJ
7alfooGBnPL1NDpAW1EXBYejDsqe4RHPFNwromM6MsztopsmN6K8ONAlfFbBi3RJHrBNSv0M4mmD
brOm+NLaHIa98Ki7ae+uMkR/Rc/gf4nOer3eOU0SEgSk1hvr2UP9U+8mqjYvVpuWVCKCVzILHPS9
lHmR/UQMsLGp9s4Tyms2RYBNLCVd0khlJyElLmYmJc5RO6TymwPhp6UlKIRCL/v/lU9O+IJxAy/2
NSQ4a28WBCAMxNTWTAJjP03GM1vnX1vdxN/Nz50Y/OtT8BEV1zTquRE8TJQF6/6il1H6Bn4LwSAW
EPOivC/+FOgugYliBCvacMWXAVtdcD455FL2S+qokeFGXJ4eUhpCzi87F4RIeniFTdlpVQC7VSDW
7kZdz/AEemi6SuPtxQVg4TMAaq6b7koiK/tmRO4fw7CsmcNqI+3SLDTYHvfe+5CUeSbmHYi5RiQv
PUHG/IM0BV+I3RPGGPYXlRCzOkuw2G516C2qe8M9xGyBm26t1la1BfGMbvnKf/AS9XXZ0ayT2RmX
EwgsfO+gkS6rY+i0xeLsc1l4G+PsLlm08XjplyluX+7MmTQZMTv1AteYkKM51ISWz+8sz10Y9SUO
0sGb2BI/NsZvFRelbafEPssrBVnr1UgCDHP6R1plpCZHK+1N36ZGdPNiAcxJ/bM09m91vLs6wioZ
nDuMEOS3r6ZhANgzOq2fOqXQKkDG4jVBAWdDoGZD5LoPOBty4pO7VxMnIkwcJpoaKTnXaCbeCCfu
Qd/YGuas1NJF87HyCQM6evrsXcypWNw+yFI0J8etJpxMfXSP9z3YSM5d+nElw1sVjdVdh250M61V
axKLHs/PYqd8Q2yge8Iaj4vfsV+kGjLq+8HZBLlHuyx3kb6f+3RHrglxREtgwIvZlnEEVzuRl9rG
+QDq7WKgupEZwg6G0kIK6lv61SJnSVABcHuDoi6qLmLKH5dFAiagQ0lGwfGrGMdemCaElxOSg51o
jbcV+6OJVCmbcgSk5CjJLSmY+YNEOEb//E1DsM/YyjR9vFxA7WQpo95dXr3WPvLoLLLch9oU7W/m
y1AWdyYMQYSm0J2I9huG3lqqXr6ck+m7MiYEIqsWPMXYeoxz9BrpSnRhoo6OXKCGd8i6dHA98KDb
cAzz5KrJOARTy4DBeg75DohbI6Zv/dr8NEVKZqQe75eocBpjA8F8l/oYv6yRw23GRiif7pKILSun
f41TYnoVYRhc1JMLBqcjax7nwBxFSQZRVpvflAL8zSIpuA+ifdrF0R/bL++XxrI4GklyVeqtocVq
cD/G//XJYkJimNnu9xevfCdnxoCnOCmSlPfAUEQXGiZDHTn0dhM79jk96i2RBALQZL6Y6J692HD0
KT5iCK/2khds7GAXbzx+RZmuP7Bw78DO/49MlL6JIX7BNAdKr6t7M4kZFvaWrNmjBtf8eBWyB/wS
LFOtdnApyicqsJ6zzu9H+F5Nzv+GiRMqzKwqKnLohOOJ6WsrprF7v1Fq4QWK5Z8dZne8ZddMnIek
HTQPtGXN3HlPiHgjeLvY7f4xKmQ3gx9sF2U+RKe5SkJcLSAcftnf+HdBZKW87bjBmMac8lzH8jMA
TyN9Wd74jBqAgSUOmPn5CabE0hmrtPgGh5oi6B1iIidzlzmkPraGd4e2nXsE5MlM9//M1yFfMfTD
Ce9MQq5U7PGeTZEok46WhmnuiufcWXoweoneLxrdZkBnlEaR/kWmrLHSJzVZT+Q43/qO33LGGPX/
3DIUQJQd3y/XGFpUuNZQMiXpIIhBdw6JUSz7hlbvkMgQp11fKkoOHGKCehNw3AjLI5j0IAGgpuNE
/TnqC15tvrOetehWVRm6xT2TOyBILFCCgKgTc0/xgbW5Pt8yzKxpeKwPSeVk054IH2Ne5WSIqEMq
lxgMQ6HSCd27zOcUno2dqJ3AjEW4+KDrZqHeSo9LNzB7HCGuq0hUn4wHlbSbJb3KV2WmN9APreT0
UXIZYXoUegW8hN8B/NP7FOmv+mZ4EXlXoEGO+CsNrBjNEVUAAROKCFHVaTMrPQqEgnZGv+DhgrLu
IHv1smqc6LXtyRIiHqSjoKFdBCCrmbfbG4IxBQuJ5uah9z73qVh/harTfQerlcWV9VKvefiGeZFY
+wHDRPyYvOY+ML4sSbQQez0bnlfJgpT0NGN/1epshlgm+7pMW8A5MTBThZFY0Qa41SHeAOZ3YK0+
pjsKbUfL7dq1Ee2oxeVa0knKz4nRxu/HVriAAHPRNEw2QHohNKeGw08q4j3VZE/h8644Axe7JQud
+GTh5UUrmAuDXyp79m8fUwQamChBmYXi6f3KiF0iw/6/TnUQhHJHbc8jMivlpOgF9I1x3qQKAbTE
lR+VVHizJfxSuhGJ9GT3sbF2fJD0ex6TPZMjzuIv6vShIWwKv6WaINvERrJTgszcFJ6jCwXniOl+
EP6bY6NkxhbrznCjVXprkN5HLLhpRr9dOD0sS5wJNr0vSzP6X/lf9tNMJ3JyAhfnXk+NTspOBaYn
u+yP6kywFBnPEHLCxn5B6tbJy9lOHFI1H0SdQn9ijSyEL3KnLdyEuP66Vfh2v2kwnlke5W4rjYHf
IU00fGlDFQYG2TMlsG0hPFeE/NzLjH9IZT11f6sie1+Dp4ucvAKxb+gwUIFC/gz02DqwFdt6nXSb
zhmx816jYWZruQYUluJq8mwM+oM8F6Xg/v/IPNa2yWiBiF4A5SF0ZiZNOynCPGwQC1u76AgIG2B6
phRkTqnZ2TjtDsZj0A/kjwnM8IQgJCyotl/adnk4kRQxbmzpULGCLXqTWVqT0tDZDxNvJTsiJx4q
iFfY3J0donawUhplwHPx/1oeJv75oQysb3j1tih4NSbRTpXINTN2Kvm1jv8Xtzt1tdYdlXuJ/A1V
NNRLO8LZj5fFW9LEpHNfL/pSL0EVpMXOW277MCW9slPPNeo48N4Si+Yl5A1dOJQDPeL4XYIPvo9d
52UEYOj5nzeqEhJRCA9871Jbfp8yvarkXtnAsj+u9GE4u7wToZ5pBlL7N7EXA//NhGcPOOsNlfhb
hEp4uyWAtZribBWfWZWLTcUeKmSriEy1ESQfF7B0Tj0UrtOQetiC8sQcv1qzTCEoDkB8RSTMow08
lXzFe2ItYOgsfMs5RprVb6irtyDwsvTCAJwYizJAcZ6tCWx4WNf1cXPQn/ejMifGwwDp0un6ZklC
ZD95b4D1FQyqDQNmodr3QXDs8KJ4/ihBOfvsoQAopQMYRpkz0i9QIrz+Gnqgd2Vy+MSgq9E1Ehh8
LYZCXEm4niY8fpKICMT5XdEE7DPgzGMQxi7aBGEei+QIhss2v6NFIF6T1LA4eDESkIQqgrdAxAvi
Q1g4RrubJmS9e3IzvIzWRsQK9uRRz4gQY1Rk3KshtiL7ej/4dkRjhqcduv/HpW2GuFIV2QkWJs2J
vlkZxyblwCHlBroulxI3XMfMaHWhuTQqC5b8rrFMm4lWZvAtrZLnkfczx9J1GwMXMHPmYOFr/Htm
FBT4etbyHHXUUNOr94LUcxAV2jZBHKBmTWeVwqMHab2Ni35pFdNKGjhU6q4lluDjy5gcd4ZXxIWu
V6CC/0Fa8uu5vC3tGHpp5cJxR4nuoJZx4St5/IfeOL91V1CcZgNobGXUtAQ3R4z1XMTfomQ7WOyj
+QqRYgUOpfz0XFjJ81ED8Xa9zG+P5EeF5yjps24YeyWxtkkyx3g4NLYNHUDu5nuFK5R1C1BCvEuM
bC+maaHKfpYMm4xCJhv8M6K6gSY6N23LQz5BwEjJimD/dSZwypyAjsMvCVC034GqDn/o77gzoKYl
i8IlBYy7HuZXqn4vb3GfUUE9+NptRZX0fq91X+CBL7pvKup1yPwy++e3+nFrKDV2NGJk4tc2EkWe
qReYHQHQ9GpjF4nJoeyOFaTZWz5Q6NnX3XrJM3bnGANoihLZySGu7151ShubAQyKYIEi6lOWK56a
12/sk1Oiev/lDPPygtSsFRtHOUIcVqZefIxg+9+dwzZ3++XbGJ7VCDtxiPeGxQ4upeYSr70x7/Va
9C61hILYtOsnoMhU5mN05NfWNjpdOIr2OwY9UJigdMtjVXLlRLPrRCHv6FEZzKAVGGQDXqDwqwLC
8a2LHUJreTdVk6JGIuEZfzX7FX/KnY79h2a9I4lvlx5KeyU9bxKiC2hYW8j0a8LvWN8kukiljpw9
P3sFXPkPgPM0Y/+1+bcChWdOt/gEIMQNerWR+yqPuylr7YEEKVDMUfi0XduaP9H5NTyHE00MJ/wc
m8/aWSWoUdLX4p9AfUL2RfLF7wzyUUJjgYOQdT7NYXoIc+rMMYklg8K3IQnEIFGWpinsvD+NUAXH
5fnKcQK48PptM8wd44uI9Z9DuhUOGIzmGU/S2846g6hhomjpwDuladMbZVmhuaN3tGkApoeAD+am
0klc6/SroNTqR979S/kC/EvLbsxAPKmJGbMPUIs0WJtQmFlCeqQ/VYHANGbEnjF15sFlU/0wt8t0
wm2A2Jx/xsMDzYJi3sHncqGMQADUvVlLwZxhTYn5wqQNJid68sj1VQm1SJNPf05jTteInd5nxX2D
qOzDdIfAA8mmD10lt/eC5yv0OTmvpx1B13avsPd8qp1BC9G/N21sv37TYeA+AjU2xEPUmo1Q2QDT
gTBRcMTxGs4/yKLVT1wcOOM0hP8uzOIQqc3DoqTk2j0Hs9xHP4Q/Ev8Q0vbZAEfeJ/BHkoaHcSG3
6UoRqshojyZP6Z/RgTBk4bcmNYkZczRJDuxJ+8b8/oFZ2rwy6+ImhMJVC0Q+VaN5nx611pcKVNSX
dPYc6E1scaFIIbHF9BlQiXLIvcu24crYm1NmcEZtVPve8897oq5VtxefwKqOD2Vo9vpbGA4la9+u
yiDryDNihbcchsErzb1F5G5q7G6qSUXC0+wrx+anGvnVL9XzvlR4eMDGKS6nRH5ucTK+dSBuJmbr
7e1JfQqmv/lGJwmNAgjEHEuGloNW/zo9N0Uu/QYOhwN/IymqmdnzDlShvW0PAq2mDzzIrGhJkqEf
7rL5rCb1nny5PyDhwhBR7rdW0pg/+LnLJXBZaHbPrhLPQDZ2liP5+XTl7n8nh58xnS9T7yZyshwa
y5mrLyb73v3rjdlrBI27kR4yFDffd5pP2wWvD3wAEFlGzw52cJKQCYaglq6a80z4gjKsmkWQL32y
yseJiwRMf3tNgGQAx+Klxb29XfJnAaDAX1WPkck/Qt8jKsWZApkLEdZT9y42+yogjOoYsdi+aXsk
s3CiSjchbDG0ChrYtW9a1WHhkXwbhHdm6oRSO1tbSXnVR+JNDkbWsp8YHBj1jIi1L5R52syXQ8qn
5zMX3jMbzuPrOieQCP6e4R+tLK4Jag9XU0VzpdD9Bx9jnS7WD5uutJ93T8gM8O0WJfsAtP1xv4gt
dGn7f34anIRKWEjfI3pF7C4FYoD9+PlmI31eSFZvfMN8e2oU6Ccv7Uob0uhso0udcdoWf8KwKHtW
Y+dCZelvflQcPc29rttA49wzKF+GStMXaMjuLvlD5ox7N9zEDojLAp5MN61shgzhRBA7GU7Fo1Ac
TE/MVKu5t40K/TjD1cZXMeWA6qQnbpAyFs9/6wFwIhAagvyeM6guV/e8vFs7PqR6M9yoxBYklcBT
zZUxxiQIIe53y1iWPtSYwsddzzCYGkYta/ppAfWaPKysgJCpq3RwjH3MtDB+bi4OPMAQoFhDO9sO
6LQC2ViHVOgMPaMvbKmq1nEfUnWT7921+iT6wJ4MAeJfgMgo/xGxOaMqNfmBsD9cG2ZimDHq+WDB
zV1ANnLjFt5otV8jDi8kHxI/X3mt4zfYm92ZMddjmUBCVyjAbejnRVFJly0OsvpMjQvvW5vrmMtV
xwPOcR2rFBN4dMw7A6OECEFZBWO0uG8cSQiAsPht9UwaUou2ytrAe5JOMIFWXLzxxjNVsNito4eK
szOUvBaQZZUjHBwWY7siCoZYtMWnQc4vd8fBTr+ZPjDDf048EsMLyKC4rckDBG7B9LUhYEa75F6J
j6QC/aXrtXTjJdJuvgW1sVt52oxGYSxAEXzLrh01fsjHinqmXNcIxoR6RVHn0RZO6NytqQW8tqMO
ntqGpag07EZKdSzlmxI7W44Z6AKFbvUO2xMpNxxtgAvW84DgLmQmtXcr3ugzqz5l43QE5jBU8QZZ
iuxZi4yVT1PNGXkdEhavmvwLvGJb7W4yl5V09ap3addZcJo7JA0M5CIWEpfbNSXQlUHt+yRqDyDC
D9xI086YPYzMIDaJCMGYdgxj+CwrrSpbGgr1sG2xiTBr8HRvCa9HcCFZjMnP2qOHiz6gsJTRWCNn
ex3BDUIJAgIyX00R/Gy3PvQ3tmtaBjqNKUosXVt0LZ1Yqt2Q2VYppXOonV7Ur3VgQLnzg0Qcn5/f
CLztgvf8K5b6L+QBmcjjJn+AkXfx/ZJ9TLHDEfesEHkf3+qhO4sxx7CwBhMJNm6FRCkX7EtlRav9
KNHCA7qr+0QjLjeyM9R7xGcu2ZyG8LgJhC0vK0hyAifjYx3hgwytSGwfdjZ1zFRCiIw1Lf+/BBzE
qqWy5RrZlOYEwxgHyQfGbtxqmy6q4avwAGUjS6kdfVJu//u8y7M9lNquS2GmgPBgBAPHQAsfgUaI
JMXYkesjBlo8Ka2JB3nFW+L/ZOQdliwzYs+UgHK7Fn/4DuWl/eQ9M3Unb7cCyglmx6xzoMNGoMvs
df8DQK3PCuteSjZf4Ibm7frBxeD0E3mqXfSgQq2OUPJAqtcp/+uKJw8XMIiLNoL3caFo2AJPqjqX
1BP12uE6DNCwQKcf9+7/70ogCcy/ZnNeu7RF1IY5EiWYLmbybMJGY5vCBeoD0HGNeo3b/mOAwuNX
gw9XJdlutUPzszqcQTalIzI/oZJWBQ4uWrbZoW2mm0SckwqyqxYito96iwBWnopF56elKrVnPS+6
4kqYVl4/JMl0GIOeOB07UTAycNS8EC08IAizLLKOW/W5r1xus5XwfCyn9SCJu/M1B1HIWm06WoUe
qdJt4gxbrHLchbExN24DQfA3dhid1Pi78/mR6eQxO3MJsFSL4EEFLtR9AhBECff18RoYMJRzMyOT
IAEnBP5czG1HVc2tp8k6HvXh8+3iUirj2d/Ak/E6caBnWwR2T1MG3UdBmjWu32eDzADPgZMsVIBs
97uJZBcWMDK3lZTdVJU47HWNGR/6D1nmNEkMb7eawhPgNiwOq+hTa4P93AADSno8nnI7agdWt74c
GjsLH8rdbTmsZvNWoeZsQXMINZdw66eryu8NDu/Y8mbIt7ZCOzZSgA2B53K2YOWiSaOuuefyFAPf
Lfc7Ru2Hff8fkOidK/dE3uUskLsEtpP9aORsraW1dp6ovawMoF07+pH8YELX+ML9uj8OyBVeY1HJ
+fPb8uNHFhHY/+mu9FUrul1YLq8DpUdahYz3tYls3piFNbOn7hf9v7TEv53PNosgqWmBNV0u2Vkw
utZgTH2hn5KJB3CC9t+5ZdXPuj9FOO34RbVYZ7pLhiO5ZKu9HGyGQJynK6mvtsfq+0EnS8oBZnJ+
dgpOD5WrOKNJD7WvoW6dLNFBeQYBo4xLcJJcHFCHpkveQT2n7FzhxMqDjFy5jxhqKezn4jBGqgXn
lTN8wAbzK5kPQwzMMsqI2ItnMr7++4UCyIf1Y9JwacTFboXI3CYg3PkuJaULyFY82vokIpkPfnY4
MZIGLJ32HpuSQuv1fJM0WZv8ylVwxHMvPGu0NnNQ014IK4WnzNmywq/Yv0ovZXumMGSGjePIRHrF
cVs19zkqh3QhRbXr4jFsDKJnpjs4WUsA4Br3whUUYBR39aKrtBCocWuuXIRmcE7bTrVUSbA5N/B3
r+1qyfHOOJrG0GK4VZOI5aj95UpfNKIJjSPWCF6p+SUYqRlirytUgRcQUIwyR2GQGhtQiij9b07W
e3AorDEUhjRx9SVDiQOWMq/1b2qcZYQqQHbEzzNVTqlZCHetuiFPSl9vzQKrWCCoEDWWrFOhUt6C
ftL+6qiZ+ZMjMXmMov3rxBEqIWLs++QUgL+rFoTVYdLMuq1jRIbzB03+Xz4jAEcSts5zle2oI4v6
05aZMOrMyCoySd69Zc9AQax5QGOqbP8IcS5fb9XLezkW5kYFfHIrx5UUU+O3OeXgj17zA6ZF8cWf
etI2hTJVXg5OCURVL10DNx+eCU/BN+rQrNHwdhJvDxTjkocoPI77EWdgilL7CmDcxfgzVcuhmlnv
+VBqQQAV+YFUGnUMOJvFmE+ARz/AtWvslBw6kuJkjF1n5dA0tWj8ssjl459msNG+5WQ5ZWKst73m
YAmqA1KvJbHJ759rvFgKa2/RUY+fNDmEO5ofuIcAPiWeqba3u4Ok0kcLmTqqANkF46ognQIvdEkK
vwZNAdBjLKGdnMJgjUFlPXONnwiN5tZynw5ToLapFtgtdykS2820kMfg9XQMTuE0QwK6Lo5IfoSB
qEvKib2vAMmMswIJ0+tU6J2dFvByGdQQncRY4SV7tuNb7Y6dYTVjEhqbjaL9faJquWRttdaRwl2q
LlxjF9X8W56l5mW9EhvX9RVF0ltAkGI7z4vyayDaRoB+3Vdmp9pwPg4adYMGCAvICD8x8ynADWwg
Xsr2CapEWsDZvRifv6GthuqusQu1QsJRZ2/c8TkYRYW+r9obWB8ruR3uZ100YF2wIPG5K0o2BsYp
Ryi6Vm4p7j8r6O3zwKcl9IQRbfkarv1dFKAFFCjqFqz5qqLusEEEkU4T92eb67wl0xNY0O6vW5d1
SgUde+1oFtPUkCEcoKxp1QdQsincTsFX9W2TiTKJUYT1DcGji6qyN9CSWWlVKsm4JXvVWZ0XzwgU
0kn95uXq5JY8haB2eV0Ovk+IHL1vnFsnJhg4otv8YojHo2a2Gvm0ZiQFMY32Vl4H+q7LmK/hYliK
uC0CAgFAcge49/F19UQ+CccOMFrl3pFV5vaq/tuz3c3jey+pJS+hlRpbl67URPVpoaDvl+vKiHPc
xi90IdMWYUFwDDvjZ4WfUCjr0FDOjQduuajq0iToa9s0srdHCShKPC7KmnKAcaaDB7npz0vgXR93
/aAs9to/pgBPHus25KrPRtZ0bKS6lKewg6rTeMetaQ/nb4bCmSuJ165pWebLmfIog29Pqbtm0RIi
pPLkqqLsFSwCBDEzc+o6USS7D7QsaMEeQPbflv2DRbNWyFV1j24vH1ZJNUt16IJbKkeWj1vX9TA3
352hAX3mq9mG3r89zJMHSkGMiLcOurWSPKX+3xJB0p7AESWt6LB1PVmzCYQYHPE+pOXDh41kYAc6
gRGkHGb6Ik9QbZiAiUzlvicOFvqAgSz9reW5/+bxt1mwykmR3B2pdexLcaL4R2BmTdXyvoVXL8x1
ZJY5MljHzrmFLlzmGzfimAgJMKkyc4nKed1vEIEvBEvksUpppvDyNZ22f8QMHs+JUVbs5xhX0td1
JuYbyh4C2U0oSnU00Bwawh2NDFWiCPqeJJhPSb05IgoKhQwQHebfpzuQU9O3OwccME0sG+bLiyuu
WLVHHkQpc22aMad75ZI+d5vPB///E6d7iNbVf5Vw7p6sytO+hinWUDJTdLXgK9pmiusm0PAZ/Ezg
tzJVbPDYISLduOTunq/a2+AjqwtagJ5fUOlAMpmpRt23iKn61v53TLXZQLmVQzxhvHJYq00CSLpu
1yCVoR9l2YVqWHeNFSFrHHoBdXJhGuSeFjdkRQwDFfYGzMEOC8F5/JGtsB8E7rRHp+uAbKrMZWpH
mkQPkowuQ8e7XN6eiBNO5F7pVidj462/FxEfno7ZIZX2I3get/dTMUUuI9yx/W854NA27Ijcy/Ff
Buw9ZGDzpHXEE3xb5MfHVkgybBDvcPjmNDTcap08sqN8hQoksYNELdmqEOs5jzbX/5CHkNVGuCIT
PxnJaiHQpD0dFOMyhQCBrWs++va9N30jXRtiyD8L9c7GwdvHkQt+SD5FBgTjmnAiTyvZI6xdh5Ak
og+G9aiNS8es9zYzc5xZJ/ruEJnS8TmHwVrqtGgCzgncmPbTNO9hh32VXvH7ztKsf/gy5z+k0Yg6
UhigQ3XCuwhmGkixsfUgnt1kjVhLg0vQ6rq/hmn5kiOgVwbzg6LFRiBtlnzkHYbK5MNzap3Gj9ah
W2B+mD5zdYuQ5lpoGNiW+JwRiMsCNmxl+IndTs1O29Ig+ZpNj4+6KwQV7meN5OjTA4RvM1GH/f+y
BPMUIaj3AmTMPI9RRwD3Sz5gW0Tq0GButl6iVIL/hB7MQHVz+EbnTVyXeAgdwWkR2VSTXwAUmuZt
/OzSOWj/7IOP0KPMHz3TZ+UEeoJS9Q5dQ1vc875m8RVTXBijpfI1Q1yvgx0V88KKzK2I/YmVTT++
hswlPldgiPs0JaOkxt6phuWEB4tf4+L6HPSwMVsRiw8lGY3KiEa8TyCGovaxM3MK5r6r1YRk0bY6
KLjn/hFbEJBk1qrRy7uzj1plGFMUu3SCC6/R5oACm51xn0MMdxgPRVZ3FfAZ/zHhomQcXS/xP6z7
/xAZGqFxV+pq6NlFKFeNzcOlz2pInrYGLF2nb7ahu0qrseyGlNpGhHj6wbvEEaJRxKqmq+xexcSA
15N+0SCUU7+1UHL24zXppOJJpm3FkVFc9fiIMxG/pL/e1MSt0bLZSJ4ZciAbBt1kfmSEpT00mzYo
qE8J4eImOsSIGSDwh5SyHYo/b5enD71I091LWnYMEEboQPfsnqb1dE3iG3vcDCZdOithEZ2cSKR4
ynoLE7Q62WLev4RHHZQqXK2rGDK54p+AKi82qqd+18tcNva4oZFZRVNBkxxHm8ttNSWaHvdFSwVg
JBeZDClqh+xw43BznasjP5F0ZOY+jQ1ik3BDB15VUwMZq8rnVRLlgdxn2ltTxRAcCdosN57BLoN8
ys2M+iq60sjubbnovV15qAoRsCjBSJCg+X25W2gJxUIVKs9B6eO0aGxdqOXX7y9QvlovoV8DhsI6
FbInc7AnYPA76v3QWBPJypfapBUjXvCnCQTI9onxHGPmkSv4RBXZEzeUmmIBnBdUn4bRDhXyzulN
K3+zP/Mgdax1YNq1Jvbw2iWIhb55LPu6L3gvMiJ/VXHCboLTEziiC0NLzuNl+2KkHmHhFvpfVowd
L3pFp16LwLPAIXx3yn+gLAilNv3Z8e+iimJz5GabodHekHFIUXip4bds3d5Krennx5a4UsP91BmK
UKkR5KK6ZNqbhPRu4PNEcpHA23xciVGnJIo9MwB1DrJ+Fn7OWU6ChhlPrgtns5kI3QZhFk50Zxl+
9NoJlyDq5a2gFIWrWbMs0pL+DUOZC6lrmeGgLmV5Wtv+diD5XCx80vV+paUeb3Ulf0tu4a8VHxP4
w0oZvjYx6hhAzBLHl0lbitKLHF4ener4Yh604VUx+NKW0YzM3sQ4qcznUenkyN6e+HjlzIi8Urcd
wFvZUQuTg9TZk4Q6xy6xsonVwYUZm5pm+doZtLq3vPmEnATWC8POlBZro6Uvle+LfVZDWqP/2Qe9
O9Q9SL8NYASrz8CXv1Jp3zNIao3648sCx0Oq/cJa6csCz6lF95Vy0oD1C60JFQL4NW8aXrzLaRCR
NCnXm/RgxRC/XFFlB/MBvpZSQGF5EDtDLhNlYed9FCEKwZEaWW/muxsgZ0JQjGap7Ds89844pfnw
IPUawd9/2w1Kmau8uizcVkt4noijWtcrFLAvB+S3OntUq20pm+6Nb4IjuF/j3UmUz/0zdh4WQySk
kLKj6u8BjeSEL0j1+EscMQwrUvu3dIHdqcriBwNvSYqo5XiajI2uVYShg0myldHrQ/zPAI3pXYfs
MgOLdd9V9UTGYErJEv/hCb29gPyqwG9DI3u1fzirelv9Jo4ZFJoRF1cbMcGJ/snW27j5gbH0kFpy
1QtXJPfhAoAI30Dy22XFTK2YZfbtU+LHIiGSrC5OdkEhgfQ8vj/2togBTOPwMZ40qNMusBze8RpV
+NrIB5aMub5hd2Yr6LVIe3hwIPm/BUbiJ2V7Hg+p5sPcTuCK7lEpKFu0Z9GzblhqSjbfX6+YsKOJ
WMRdVGWeYhTREfHMn2LDT59TRX4AUZgJ/uTTrdanInHJx57QApjmx0rpzFPiYtRbSbQLpJI7PNkO
Om5GllwvzliOl6/yQa56TBZJTx/K+QM9Iv9Ec+AMFaxk1eGH29abby8Ut7RMOgawbAzDuWICXG1W
I7S4ZwYoqHts9umqW9ZRVkS6DjexNeyxpkWSRvW/ifWhhCPeCfKHEIBV+YSwUsGq9T1lAVnMPZ+r
hkS2FIJqztctZnA1+XBL/pGvaYINe2D34UIgYTo/U/U/3wfWKku1OeVhcfMtpfrHByV2wObjue48
JoirWYCqVpSlydtsPflQezjl9fkvHJZe2XOBtC9V55qdRvDBWwj5PtCt44feMSGYnS6WXbUQjd3E
zTA3IwelOqdGG+ITbVfD9GmcJnmk+04me3X7xaB6aWRyX6ePXQMRRK9WvbdQj9yULSPiwQIH0DAS
rh/MMVpUQFW6zsjTqw/lKT1xcmY3UP94LToaOw706g9L4GpwCoa3hQjeAaoH4zfg2uvsLNFnX3Qb
VDTPINKwpXM7hKVlBp7QeBjIi69yie7WqnPRJm0akgKkVksEnueV6LSjeT1G7XcFF4N6/ABVTQyi
6936Er8lPpmd3bZ++yy2UfNAKh1HuBsH6K3xPrWVC9E2ChmQKI72H+2Cd/lURLKg2FbXoB8hUJ2r
Ybn6RswWkFn17NPaiIgW1K4VZ96f8E1Q7OVi7pcl0Zd/FQJBXuleyKd3g+ZwIBdQVE0ZOy4thh7b
mz249/IXiDCB/tgpGiznJbaPkyWK6RZEZnU3ZiljPgxnnkTWFgd9RgYHP9VfiIrEC0j1Mkc07HCT
FDt1CsZTCwwnzha4ysH6bfY0QJQDOMMSQIwrAZ00Hn3jL0FeO1hCDHMCbxvQ1QdSximh8oEyBIbP
ZH4cOlqt92KfOGwoG/hZ+wBm4RbzHUgn9//UCFo04UFqcCQOKQPJPrEVJUGrEANkt1j93BCEGc7K
5tsa7ZS/l1M/F4930cekPSiv//C7S4TbD8YyYzgYUawpe8Qevru0N4zD+wr30plpIO/76ccAQlG4
2SIc2qR1fn1gt7wFuLzSjok9ka1QPnMZCpdCw6TnWC3AdKGhoRVMnSR4nYgg+oSQbJ26l4pb44jy
mC5vObe2XcrcBtlpCPCNgKSuBmuCUcsRvxzVP+AV/OyI25tWzWo930rwvgH2IlCLKrOLcs1zohY8
Nuo8CpZAUZu+5da+7PwAYmJzXmulYMzTDSHi+xAQn3xsAdwVhLDlHqBhxqV2jL2o9vzVbpGTIR9E
k321EOf1lJadvq0UIrFV4a0wNQDbj3b0uZMzfpS7e0HrAp1iNxAB1B2a8GCtmm5tTqKojLTSBkhh
L5nwOymj0BQAmDs9kyD+M0LR90l7K7xvfPWTEuYqypF7zIuqd+dM42X26jUL44HrLVgejX+hNamQ
zACkoVtcz8aD9hsWd8iPLM2dbhRE6dFgI5RqP1WXr7MYxcM8DB2OlqjB0EcbBCzCR25seUxiIdK4
+/NVwjbYUMIWyr+q/Uxqp+H/r9PflKIYSO2Lnx9fEqldJksi6trqOY990f8aOXIoEmnh6Y/BIDKS
V67m9LIW7SWtn/RSiBBE/CgPOuNDm9vkeBAIhu37T/YAkvpwbR3A8RgfNnZPuyqMq3kuVYejfvF+
4254D5kJQ6uBcIeOnx91r79WqN0bWV7DO+RpRzksqqErBRS/urjmbrJv8Y/nuMUMfTUhcohIBDM2
FLOrWi0bnv099zk8AF28MOZEqls0ffVTYa16FfD4Q+v3udTdd5UBtxQUNeBSEnVbP1a7o+STfiTP
CQ23YJVNVIVh0+LVcZygiNpMQ+3gKBhmthNMqzEcvRixOvdZNIEyyqrQwSMVSePYfl87ySJe//AS
HfNkpxKNDv7Hp+TYyA4L32hGkngjZg/dwIyxjCOGMvZrrIyApu1PyHoG11U8PFMyA4v3ktahyUlZ
6f68KsPs8e3ogX3PZmCjFcgmbxZZLo0beQQSdAbGa2vR/iIJfX3zuBxy0qprU/SMrHbZo8MBgmsW
L+1CVoFv8fyiRt0eR1R1mkq9/je+togojZ6GN37l5UwJaLtKlQ0E/0OciIAtV0a7Uq9/HwQUEY/m
s+a5JXMQxmgwKbSmA1dN7Cgs4YFtenixhwziDBVPontsjyBBDgLM7PuI+xCH/CrbDop6syQdzll+
tVjQII2YP1+j7FN8yj+SGH4W+SPGfWcY/hl4lhY5PKklzkGGaqP76kTmBFiY+EzU+ZBiliYo6h1A
+JvhH5Yu2fK0mhYSqS2IrkwnFPoQcCNlC+bErvlJqhkEW7N+BsB1/4TvPVgQHeQ5zah52fMu9ioL
vnUYSRIqQirSJ2cM7WPHty5mY7WZUaToRacWNEhhWvxVdVkRZfzDnvv+56A6dygegwmc1JCRbRbq
tSCWwYJUJbuCMzH4B/gFVWgEP0682kIo3A62Wfg49c6kuYqzAZSjwYfQKaTc88CJ/wXFMX2XyMmn
/A6L7sKgVLrJAWbzsL1yazeBp4dAyhnudW3gmSbkTGcXyb2cM131pGuJAcGbepik9bdIpn3wyHI6
zjAd15lYf9X4QpwvWYnWSLb0K5YT8Hkvw5Fg0xjVX7FevW5SHudBfv8DInkZNCoOG6PGEW+ijB2+
Ro7D8ZRICd9f/GTSNxCSPTk999Y0M3cy5+HwWeYPyP6ZhuQH9xR/lenAxfBOxt56DX0pl3sVmvwC
Ixjvt4RTPZcLaRQ0cz37+5Kp19kZtL/2Jql7utFsprf49VqNVzVLX+f5tZapFh6y2oXY/xIJOWxK
UzwAH/uXDXK8KkHdIMEYI5YSPhfLOfrvd4o6FKMk8nxrzsSEYxgrj67ixEzK37KjYERazyCEpHLs
lfXGz6/SJbvfsX3S2FE2Mb12nUlreUbp0tE57T/++cdEcvsJgObY+WwTUz1BjrjXSTJLEL5fOyUV
SW5BJFAGdMHhli1qEJ3wjDYVieM98Qc5VuLulgrLH9Ba5uCb/ecu9Lu9Zo5WMF7Klqox4n652JP8
zggclglp+7Qj68Z1EMprAy/nANh/O7idNOe8JYjAx79oeA/v67midIMgEHAKaBbAP9F5C0Dfrz3F
JinGIde6t9W3qAMQNT0vhWjgp+pB0vr/I0iFOErpp07LCQYwrMWIQZwFE7YzkGrigmt0U2gJ8UqO
jSCSu+oFplZ9lrhz+eSF71zRIdIHmjGVYxwut4k5roGjOSf5QjDeaoy99B7uZ0Io5CQGTuE3ytiv
mok0Y7SvEY78T/JT43dq1Qdx3Z+aMGtFp1JKzGuWY6SLmFa2SJ3pqE2po7L3ZWxtW5jnHdvcK1sj
i1hbNQN8HaXogTucLg3L9QMS6RfyPGHb+oxO/M6MQr4aB1GhrX0XnIFNoXf20LjB/+t76hIRWEwR
j3cqPp9V0vSTvVPEtsllsOJS0+GwPA0UP9qYHwp4HrO8FHxHuW2f5KShxOzYhpXlmPbrHAqNczMw
6XIIUoLglXVrELLhkB7Mp8FW5iKhQD/2gg0mpjAkQZ5raVfw/8ikk4VVXgehiYLKgKDQtgd1yuvn
kXCsolF/KTtYB+CmezixqPkJwnOvJM2HbpTQb5OKAlQ27GvxKBMWZrDIsAIduxM3AwfgHf4uUkH3
tZndnTya9Osu1L+qAAhXCKqdVQQfC9mXY+TeCfmAZW9OLtCF/Vlu7iRk3F8DpJUnMYkWfVToYcWA
Pg7dXuUJdG3lkkeVeyuI3RxFus+2Dcbtp0AhMSAi1SsC7whT0s84JJzP8YCMKIv9IaOWabMksfuh
aoI1quniIsvq2+fjCRyY9DiipB/kg8FRvCdhxrBcol99EZwn3MU8loQMx1n3cpEsiqxwcwQcnOYt
i59mQrndhEvRu3WGle3P7ORZkRk5/boFoMJG7zTLXH5xUP3ykPyIxdwGJdk5HIJQbZNLPua32Sud
BZ3GT1bE5TQYmMSSpuI7GGjGeK94wpUps8N9OBTKE2xPJYT4od19GXo4ZwUiCn1kACZ8w61854C/
V4dHzkWMeAFNFo82tuqFULqmGwWE2g3s1OtEuuvYDhwXi+PC4ryLlNpBuSLx8PfYCkIi8T4nw+/t
dpqFksaib/MpvTZLGrYeAJbHtlWkKcgSOfmgN5PheBJPojH/ojXHm6vDQeS4o0vbojK8F3gXaEcm
mmtuFq6fqblkCUrNxjY8BJRBOGhZ39CILWpIAupEkyf6+tzXznpG3KOBlAEoJXyFbBfX07ZSGfz3
jGpcv3d/OyIHfBC+t6e2t61F+JU200MhjLVYUeG8v18sY5y4cXKQKgYrnVUE9n4Go5v85xBPf34D
OHPaFxf0buP/KE5dVg9l8bu0tC26q5hu4x2aUbw1bqD/Rmlqt2Ncn5Lh03uOBMT/64OoBgZMB7eE
48X0w4/i+s1exQ8Xf8KBkxi+4R/1zzJ4Fqy2Jfw3XbGK+ACvRANGH/88H8msLWoCCn1YOnybPSpW
YickzBDK6IwFfZFdv4ego4lepHN/z2jVDNDexPo03/5A4ceExBdxaJiamCKEZo11bVbnBQCCrD/y
7vOtUOghdceiL2cFzYEZMksfNP+E7HruJXoNs/EqJdoWYgNiZw4DFx85ZF9QeHMMznIPzBnx1I1U
5B7N2YwzxY7fMfzVPYwuHGENo7z6jWzCj7zm+4urbZ2YhzlFiBaMffiVfJq1wfAwbgzNJxwegDCt
bKqUuzTGbDURbdkc0Bz0HErZWEcjjucYUY4ojyoh/YZXPFmHYUiXaKAF6hnhZyRoRXGnfrVDWsW4
RlbK2odAG0DDf75pfGzFec5I6N4kCceNns3fZbWjjulh6jRrCCnuzxv04WoIuZ2FmyWsyDMtm6q/
b1m1fXu+iXShdPFK13N+JrtW+GN+73TkNP4wZQWUL6rvp+TyE7cQ4tGpt0YTiJZg1mlpSldwiyHN
NxCwPQXT2xyNuixomHunuJkPwr3ruZ4HW0aqC+fJvd0vj4HzZf561KGXRz4WpojbbbaonlHWeZs5
Iw/nwZC0otp3SBMTRKBFyikBBGgMBDF4WzJwGz5AnExTiicYop1X6FQpUBCXGH841wmajI1BO4eV
bFbC+Rdvahs50GBe4nLm57/O2CpROzZoZhf4V9x90pVeM+p1Iv4aG+47Cym245+Mu5d2avE77vBE
LoxGSYoKRitDohftjCH1BfiZhjLlHzGJKMIqZX8W9JiqlOgkOdTk5v6zNVAysqI5jZPPvaYfK0aR
LdEz/7xHUtlogGsPO0olhmRiy872bCxJpVknMyIkSIozq1uaseJw28N+SJXK0S3cJkPxkiSlY2TO
7W1ULXCgAezShaxjwr+REp92Ij1ubFecJi3vg3tniAkdLNBd/XaB9xxTSkXfAFvO7Fn1lqH6R4ff
FvAghhY6DwkzxALk06OyL/W9EIN8/LXsbh/jV75pj/qc2nb1b9jKfgqAUxEWYcWop2jxe/vS4qPR
DpZC+u+B35iMZVw4/bFcAUPCBwV1Xgdf4yb+jKnNCxyOBAho59fypIXfngpYWSOa7UsSadI/woSC
eB8nFCRsraDQV2MxD7m+vczBMcnv1Rg7wqU2ne2JBAOKeLMJjlyMt/n+Xj7SDBQKT5afQQW9Tyog
LMq3Gre8Fah/AD1FZfVLi68aCJZaRyBaGCbo4THkvufJkqdoCP+AglPHVMp5Iek/wBR4duoPQd5d
WQXekkCtj3OtF82pYCEdxVWZbrZFLM02tPNbXRbwEx5PR2a2oSXEmJ7Nx9mEBnYCZb6L309MlRQO
cEk/adlxwzib1zh+n+hcBJfiMpKE7joUSBV5Wvzi14D8QmEWjeMyoobu/Lfk8zZKGYIdqtFUW9CI
elhNWiwDvf/BvkZHPmTmRyCilvD3WKLL0kLg7YFaD6c75lFmrcYAg9dW5al+l+uysApPo+KOV0Oe
HAp+SZTB+nTdMn6M7pElG+pmhOgVbXrtSDQgkE4Y0+ooWsDPUmU7XrtyPULbcYl/pa1II2edVfNS
FF07mYi6oq0eZY6M6846SLs1IC7iWmQ+RxfwjhWkbMzryMRC4SUcOLaK3VifjvcLeMAEowUdv9M0
QvQCz+oqwa+t/qXWuULrbKQM8w1hRJPCqgMcbE9OClolPKhbwpRuf8CBOUM1quoNwDNCongEoK29
/RXz6xj63Xmg51MQ2H4Qg+tIItMQihEeKt8R+5ylZIKN9YAf97/sxJebt8Q4L/hI069Lx36iomam
PtosNFHKnQZFNoZpvRuKOOjMm7BGGOiRbSQaRVbb8K+joeNuq4qKbUbHiKG+3K+QhUO32EPVU3Gu
tKEXjFHN1sBjDfXXjGsUCIMTjoicJAltIUJgNu106pp9MJrOef8MQ40HfLnDevFAbSSutl9Eqoda
+36zhQhpAp5FmePmrEIdXSaJpZZ5Q1iWgV8T3cC0rC9+2xu90KeCOSf6kHmmdImKCdI2y9HtN9qg
Zlj8DCo06Sk6rnZnPLlPxz/p6htk5OQoa7qKoKxo4Ovor6fMRntzc1TUD/KNI03r7leYZ3i3vA8c
CuKWJvs3qKzygpVao8U4lxbBw7rRt6fJDL+s2agPocXZ1d6cKnX10fO7FhimO/fylbL6L4ulj/5u
hLRcx8BDmPGc/wlib6CH/UTmr4RwQBcGvlO0yHQwE4V3nr+YEZGa/dcFLlCm//glSyvvwOisLzY7
PgYo3kW3uLuWzTydANZGblBsjKqomeeYMJyaD/ZCTPeGNk9WJe91tZHLvIAujla4pDopl/db9eyv
qK91ya4mlz9AKk95+bhePRUDv0iQXEcYewxkE4Stozbf1fLQT1Az/WtBzKphpaSu437+DWprgXrW
uaVBtsQ8yMAoNXvnm+8AJZZdVfgN8YAMAkQqScakXLqbajM36+LzWaG1Sf8q9TTlKU+eHdq9Rc8B
HIyHUcUA1s7p6CoFq53eAbZRhQtbg9sZDmpgI9aJjUz8kMJo6ORNGGZzgtTRsPH9b45gKg3zNYLf
JOAM1QeDdez34k5uO6MJDDszyN/oOarfNf7sJFvBWNWsGYCTn9oPIwoQFz9LqbKmhWxoferhvEjG
cZBAETXgwPcY9UOHtri+pwYzKS/FcLUdTtOjvEp0TjvxJV7P2PavDBAXXrKgGto6sDNTBFXcCuun
sd1YYcln3D5txU1Jgty5hqauL3O0HeZChBzqZLLrvaIBGykn+aOaBcyfZ8W1qeOkcvSlhd7qHKKY
VaFH08SXWLlBZlpBNKeF9DHEjjdysWuxZul9Co4JnKjo5ioPM061TzV2xC1tgVqWQ7bFcEkkpJML
vsvA/0/vfLNDMwnHVr1swmwaKxnQziKYL5gU1Ojo6PoouQk0nkKNppz4pmc2RA6Jn77g4XXBfIAI
KkLxnGgKHV1f/nXUF3LV5pZlx3IVkniqATaWSQM46fn02Yjk9+bCYBb9H1pzdDmzkoe2HraEpm7q
jgYb9xjEBN2nTvpjVQTNUKG8mMdQpkX3ARDM6t0lDViIVeTWzjbfB79sgtEXXFnZXh+VBy42zeg1
9JOSNSvMhp02TnIrTbW2P8pSX2ffd+Wbn2/pvtCS1lUIv7r4WRIPcNYJwdm7RC41UkKeOZ7LvTn1
IQBAXkdhjDRPs8TP2X6PZTJOyCnjDw3tXAPDwkqN0Si/hmBvH0h6lbUmAzW3MUZQ6zGGtQSHpwH8
/jKv5BGDN9VbgdidH1mPZfYPsAphFJEI+WJWvfi2JAKlPr5XpwJBzIIOaBbina+OUo2WZFniVnGW
H3JuxTRIk3Xz6KDCpt4VN2NT78QOWm0UhslwH90W6yl/S1OuofXVzLnwuNNKNTzHNd2UTqvlm2Yn
rjma1PP/8CV0/Mbg0vhmk0iGyanm8e44JoKPGFDTkZdnLsfXccfVFFDs6wFl8kqlo2fhdYDu7/Mv
T7CDt7J23wEBDHVifsx0NH5gZeB6uKDuMB2V5/uEM+5BxNgUx1yP1tx0AbkpygYoYJhPVt64aBpO
pY0UxqTw9hOsTJchQW0N91ea3FbV+XuKcvPJInEqe3Kjm19DaBfHIpveG7nMumTa5jzXwr29Eyqk
RBt5ZlgUI41l3EdERtNzGfm3pEUTgdsw2xrYcjO2M1yPgJuZ+PC9aGhLpGr5pzQAS2OeVUq/l6yW
zQkM1LX/sEVIzLPoI5EXsxCYZ+X0w8eF3SxVhfiLo8xO9oK8vgdW6SysiqejKrSGqXPnaQcviJn+
yjjmiNdCYJL3Zjs+IBW067yh0D8nUuf5TuY4wTDCPl10ifzuqU77pIAxOSsptJkxb/GEw1DJCfiV
+BtQjvk+rkLHqv+sonlkXD4Q9IkQYOjWHGyqD15w+D4h5wnxaYai5Cdc+Dq8DHnHVzuCbIy/v7ud
LggNWKQUhpV0t1/OeStlGDz9h+scIu2upby0H7nLupJlNTb9tqQbRYq3bstxCMbnjVcXJ9oX1cgw
W2mBy62aXgs5jiH5N5AEQOwYNEC/gL++TKUj55JTfG9o9FbCiOjwFdbfWzUDSG/RWFiCqv9633wz
Rj0uzCvi7jFIxu6NF7DXg/IgZtbqj+goTgaYpil/tiqYIpaTy4MjA3OV/S8mr5RIBCNRxxpFN+ak
Tb0AAjzy257seRb0x/xXPQwvX6o4uYrYIVYMfKO6vAgDteqyCX/hT3kJM1Pnp9jG5i2QX1r6LyZY
tXvmoO34zlHTRY1ANxiFBPKhaCIbygFvUpKNLfyna2UnFwJ905DGtBwUP3lPN8bBNihO+bbKJkLr
C2+ID+628vUbBKB67UnrwmxJRAEil5n+y3qNJ4AY0tPA+Sf5GcdtIbb8XlufLcTuNiUBKtIWwvR/
YfnOpF1vD9vgIKzq4Jcq7tiGmjv2yE+B6GkZTLpIImEBpsEn7GW3WhqjqwdjxmTg8nW5A59Du66t
HAOeJsviO1qE2wNAW6xttx6akcP3PhTVOyyLQ7eZU8Xi5GMqwuvsH+OJ4xdy1wfQtMjYdq3TIsDE
nn5DZaQXtneh4DQ0Ueo2JOZb+m7MY47Jy2IxMcSbGgFWZ5w5+c6TRQGrg0r6oG+nKWtRlKJ7roun
uLZMUMbZWIe9va9+w2XuJSwdKd1CHJZIvlx7Zy0b7aTFxQDUaaWel5IuRzB31Nvimak2uYqlNLZD
RGHezYoc/hlZS1GuhvARjkMLVQmulIet8sMqKyMOUc53fWf4p5wl3Nf5Mogaq1jmbLnRzomd69Nq
N3aAUnAhtvDyiH3orJXudHBP20MsS7b05OyEdFBtW9xhhO2S655aBpo57cqXuVHynJQl3u58UrXN
SNkprsB9dg7AlH33LxWMGU9/wcS0ilKCaaZYtUol4rAtJbRsGwC/G5nxJuhOw18oo1cr0FAQtA8i
OdT1wDRV0acqfJC7T9LOKm3nBAqdwaCC/0MGIAZBYQAU/NHqavtElACN1BiY4Pej3VMeS/dfXQsx
jAlynM7mwwrN4N3ifDF3Df0Y7LSWgzs5qeXS9ZhjDKHcksaasfRtxn1pFf2tsZyqC6uLH3Z+NKcv
iMebA4t34tYCi/gxgDI4jZ+tGgq9Jj/1myriOtbGHLNCHWPDlhVp7qPivw7ZO1MpgnqZoW21034w
O4HgoYXs9T1A8g3LmLVyKJlvrFHhVLPsZsXXwhbBAuACrncfo8LY9F0t0iOc+hhOVxIXvHgVqhs/
VCf/BbsReaQwjAlF3wg9G5UyheUxM4K2rqd8F+tQ7/Zik9glkpmwmO+UWlpsD76oCEcz8jBW5Qmc
FvVLm8Q6IKS7zQwZofE8AjLpHYXUaECt7UZsL6POnmxhsCVuXGqgQGnDCe5AiJ4lVwIR+JZyOD4C
G2LLF4ydbAej2TOY0JBReEB7+ygYGKqosjjabOAHIAG/Hi4xwocLQFOunEf3KzcgwDsALic932ne
QPxh+AoCIG6UGC/FBhlhIZ+Hkt58CXowlcBZahBON0tibCj7qkuDhHQOq+OaXfwenM/w0k2VOHs5
6RQEKRP/dogET0iCKv3UM4odbFWntqPUhANTmICoikQaLBJWwI7AfvlDRFWOsLiVEro53tGUYNPa
HuMOUDue+OnvT9qWURdiLsAx9s9RuVUbaCGbhHK3i5kUgmYzWCWPl+rCwHP/zvo8E5p6fqukoIpq
DCv8Z8tSDJ5C20ltsdm4k335Xm+v7BDvmRKUPoLtJWhRsc6RvUgl5SgFg7FT4QaQfVACz11KeFEP
D7n8xuRMUHzrnw7wYdmvOXoZGeoBPlSTPLvGi89n3ic72z9O/yB8GUFSEnTLRZUvBDwyNfTlhLZw
LW+qQZgcFqEPx4N+bafOx7Wh5cH60ucRotVPiDhPEeho8H2Rb5FccMLzwyTAo2410z6K5OCPBdr7
yBKyT7KUpuRia/MTJDzKI3CewIuTugjHUrp786R6sF1eXGf4v+Id/1kRtn9zBq7gsxPRpX+771br
YuYcvDVB87tjkJxvDAr0wGhB4BRVzkLR8AlKRL2/gvcLuNeGNbPtF3Y9ry/v6b/xH0JWvWCQUSRx
OjJQ5UmMwxqbwv1MPJKbXACJOVA7Bn8CJmQaR1w8AISFv+uoHekTbJjjywLD8PVgd/rMdGBhQovC
Gz1GUsG+nHm7RPfC+xA5QOfCTSvqSdWh42mMsBAjagAx8PvCG43MtnWDF3d/3Q3WE95T2iwunH1/
nG40zanEk/kO1F/y+Cp5zXsrdG4wtS7KiAqdeZrQ7urpY7UocIq3xi9ER3ZnhZaXThnvc/yom4dH
JFndallAl/V3tPJNynPS7n+2bqPKOUm5a1wYG5TXBu1uiyN7cLLxwLqxyhYNdPcjK8YO2hczgaGO
CA9bRo5CyNAxlBYGoo8MfhzrLbg/6LZQ9yQmjxZXZAwQpiDULLhEBv0xEnrTuD09fx1O0BiFuHtG
ZPZI9SRr7/jgFfK8W1TWX663dVDb1ICMKenq2Xu+hqDTP4dcvY0JpQe9Toz0ds4B8SZCuiuRFZ+4
V/hbk3ab1aou2UKk33ZODoOfD0gSjZQRzWgK5KndRfPSNNla/s7PhKeNp+gslpvUT+NVUnkyKCxD
FpaOp9kteqSZTtOiZuvu3zJIJL/iZymnj1fuv1brVoSgTLB5YsJRlHabCqIMsiRWUjX++NKSYnjv
jzecR9cEIr/rU7GIsXWWzEEiSIIBxZiQwRvpcOhlsmkVqRulVL1zgo9ovkg1s8KEpH1WJHA24IF9
bg3IOJ8XoTK3jhx+AaoEbhxFyl5xLNgOeo1RcWrFf3KLC/uKJKWkG0LS5eR+6tN1qIH3Zo6ZEVi1
ggyBcSktrMNA+jGDCO1yFOq+6TsaxxPfh5EplmIwUvyku4m36HDmmrsmWXD12cTcwjg0LUSctsIE
nyS0WsDOFvvf0S65n8Ram+gB8hN8hiOpdVvriU45ndopaFdURvEixSuUqpTimf6lOlyLVpVjzvxH
FNVpa1goC6gwZA0JjCGLNAZnCg9tABZjmNrrVJpVZ2k6wobfGZUgSMKIBPnuu/zWlL1vkwCy9TKi
r24vIUSvzgaOiJsVctH81Zyicocsk+h4n3AnRPTtA1K+OG2EUMi2tX0r7l0xc7LODTtC5DPnb5su
CtplZorQBJnFtl9ttiRKgEC/L28HI1+PPHMDgC5gBQCe06NvGrf3VASdK9JBfJhuNRJ2sPXpRA9k
UEC6nXOIuDWeF34nnWTO9G9eqzvolqMByw5Mb0CNQuRxRPPKTqEH3OJhEWq/PV6OQ2iPqURmz05/
0FuTr09sSJEV0C5FdtDZLC2CH0aVOhCcOgfjaxfOtPYnsU9rXmiXvts57VAYSFEIqLPQL25t5NRU
hCYsob1RDmmm9jY7qtyox+iJCFvSaknoI+/8iRdP3yAi+L3lF3zKdD261jYVD/yHDggMIo/P21pQ
y/OqJ1+VoHbROqOkjVbgH4X9aOOJeztJFu6sRJbvvbwG73UcDO4SrUjxdg2YP6wLTjdgyW72olh0
f9pXgAiN4kKOtpIE30bMogZs/zovXL7IqVzPV4fc2Vz5Cd2dMKEqYlGh1qvXvnAD2aY1fTZM5Fp9
x1F/DKTGsbh9TP3Q5mborvbIBPoF479IZ2hIc40rJab+oAWEoSS5w9Dy0wSNBQnZaiawPXkwVv9P
aArpCHnJ18qrWG+Hd2rByHB4aDudaCiGFwLvaLkVJh+og1jEWHxYgsgidSdxYPVg/LSkyqLbstWg
ngK5duz72wGUOwMRID+AQta19v4Apn971uk+TL/qrW2O583H85+fq4NtevnvDmPO190I8MM2apAC
Z00qEnNWSJ/vLdagjf6QewENxCfk8uxmjRB6YV00RQIsBI/WFz9hwzUuXGIZOnylSgZ9XcdtosIx
1Huirs3Xdb3z27F8IN2MCV0At/gaB+B0ehUsnzmH0IqeDcWR/XxkQcJPB0moqZ4IdlZ9VbjOgNUy
bt9E69sLrX/obZubcoFtyWTZJdn9SvQ5ilWct6nSMQbJnE/CS80HfRXHv9/+W5lpOkQcYUlD/Gxv
ARurzTBTHwPXv2ymIcz/fZxWgjCPJ7xJgbbi8YYZJE7Pml1e6JXi2mTFQhwtR2lqIDQtCAr6SuCr
skkDOlk6P/+PNesvJdRgMEF8wWfUXQ895E2niK0NIHBJAwvah1QxApXPTtBMSZD4k6uwm+s19GEN
xlu9O2kWO5yMTi24X+GucIJ0wsCplELvpPZ8boCYNbDRRQBYIF4JFPti+SSciVf7w60VWfiaPdCr
FSfsPcVVTT8PG1tIWLEeg67gXuBq6X1kv28HLpwXC1TIs4NEB4Cgj0ledY4PJ5iC2zQZ3NCw/ZQM
RSKfBtdKcVAh5y8GcwWC6/NrwnW9WmREyq2U490M8PtnNR64kVPmvIl4PFWS04ytChF+W8q70ViP
76mkShJmJitSrFjWqZ73hHm1xlj4gEsCtoxgL8rFMDiNqpyAXQ8BjvKtQBhRLS2C3qkFwKIJn36D
dY4e0zxRhPRk8yF0ILBhdFsRf2K9K/OfaysEl+kGAioPFCzeQB1HskUVmrAs08l9J951MOTP662d
OTrosUmKFwJ3gbllmLzNwozUvwOd7D6dXGCW2svT9xqDTl6C+46RTd/AIQfDUtAd94rxVPy7Vwz9
fS7IyU1ElyLBsv1ZFZDCWPeW7Qga70SPs+RHSbt4ZyuoH4YH4iub1H3lsIGS+3ql9NQlDhXQENUn
BmBGNx8tQdHpVTH8K7RW2eifUmJp5ERqWIyW1YPba+LjHl9bsgjStcc1F7nwWQaRr4dhLqCKip0X
BSlc6/Ipo5uhim23uGL15Wf+RLdX6HDVFoNUZFccplPG7xWAAzZtdWUD/BLHCjrGQJitRvCfUAFi
owQq6qWVqJjaKYl/Y0d3e6OujcNPcs+AhrFiYpOa9Jiyw+ZHGc5Uf9Sa3iGusZoY3GXeXidztWmv
G6I5P6X/jD/k9KbFdrs6WHktAAqGR1+CqZEUCndtQjr5HhiR6RfV7B369BWMoLghLfsNty0Jiu+R
uINz5AiCMocU8kWOmyZs97tUpEiucGHgzhHgqmgK+KrNu2mhqcuOHHH4u5S1/fbiKOitfd/AX60q
wwNuZ2OYW2hunEh1Bsf5hXzTJrG2jOomRtKf757uvXKpmuVVTdxOhwakwImO0bLXYce4EzA2EXH/
2qfpEMqw+cuctfM5cduTAgSoUVIBrwTmD3Ell0HSwKHEaZmHoAVUnub9G8pBam10UhfX6B7E6FhG
iodCh8/ixjcA1r/gNQbymR9q3nygRjA9lFjU6X0lEKzLY85wWcH5dumb+X66F93Zh0PmofWJUgxW
AvhjKYXo24fVRaMHggpRDUPHeo8cuufkOMouvVgyO9Y9OrnhLTZIusIvfA/1MYhoAFHK8uSkT2Eq
mHb8ON2GL1wYHoaEmnhbvZw76jQScpfTj+RWTxuiYadBCFXshH7ba6mog+vB3cM1VQ9N5NIZTczx
TNH9B250LuxuTgBXvnSyf0zqg+onYXOhWA8Ox8BxJEY8/bMsE4c08HCacRcf6xS2Ay12yg/OP8BJ
2MVhdWqFdfHGom4uiTpcy28/TmH/yjaxIXrL7vUwPpyxyWaMhQlgVgFo92TKyrWy6DdaxOIGmobH
hGj5DBNFX9FoeRZEVuSbz9GZ2WQ/mlA5MTBOTcxpfhv7eFgxBH0pmUxJWnMk78eb1fKb+/g96sPk
JJUYCpqBLxwBCXw50UdBtRhAYw8ud4JZF/fY8bWHP7xA2b0OCfwSrpKBLq33v5aWsNds1ADJdMy8
LeBGKnPbwdFuNHz5EEB3bSMpVFWS+hRGAfxAhqVnMyGMYN79MA+TBrQITPW96xv5DVbFMJyln90v
IP/w5pq53/HiKI8YCT3izV936wiP3+wO3SXKbAlqVE0gTaxwRk8NtD5gE01837opczi7G/vjUACR
SaTTtjkf9lY5knU7HeixxN1D//MkjoGpwaWMZDr4dVL43FODjLKMRUalzWKWf4u5x9L8HnvQwsNS
5/jFuyBLTZ3qwFTszMVhEXszOv0s52PbqjhjdUFZfmWheIa1lwDFOCqlwVFFiV1GCLdC8iGckWui
/21C7THO+mFLa+D+Tcm1lv0NOLXxCrflwXYGeua8t8ME2TDufosf/cVzojJKdfxCM+0QoWlJqPge
XBL9XcmrjGAIT2eRAIBrdGnpDQjZ9wzjI/zvemaQ5wayszxB99HKuDQmuQyYKIkteBgq7kYh1Hha
YhLAOZijbQyJgwNEEBzxjz+abEVV6R0PWBgMyv3bMXe6wS0eUhj3k90T1/S5iQbx3ePPVeyPn0WW
i0LAJ/3GT8BuTCH9nES6QObnSUxy1qIc2mjEI9uMvYPQu8MQEs7zh5NJTFPwxoFr5DRPUcQK3HL3
d6tyWHoXaAlHdYHQN3FWD5WdTrDV5VgRlojfS6vZrsOvbXx7c4jozup6lid1r9dD5Gfk6reb6bzX
P9fD7I1uy7hOfeRfzZtddxM9+vVPC4WAxfWGWvgTLCT00d3rJ9DC2YoYjG/hgkoyq+AVavx4FyWb
5Ahm4YfrX0ZulRzIvz4fM7dNnmP/mRuTCH90WV5c2i4oWxE4Z5OKOMOZ+9eOg4XTheRb+fMOCFCb
h0iWBcEPtQehJn9YiynxYIliIJ0VBTSl9BWxYI385963VzdC1g4EFGh06A8+gcnjZMlnlfeJTd+U
Z8PRnPT1BP/pjheKZreGZfNNV2ppFRphKTWlZFK2j8Ne2gl3yVOqEiVs5jKughkZboEaAM++3iHO
CRW+4ReG8kikzVY8ZT2Ijs/CPfe7kByvcTAbxaTwiUMJjkUHP/Pu8aScafjkEQnodqPoTu0Zxqga
VaFJz2E1dyVR9I21C4w6H15fW9kG08gvdE1eiZJqdlx33YpgCCwf61FuHAmHzcOgRc02phmyrPt4
+6IQjWUEgsioaOuJKlVyINBX4GaA5qN6OZ2lJG93GBdNThKxw/uWlIY+lCDh5r15DkHxotlv0DMk
wnGc+p6o7urPw0mGAX30FUn6x74PCKRqYE3XCzrnfpUt2fqQrSoigV4yQKGOjeCLFi8Eh+JAM1Ym
sqUeoZORhCTLNm4uRT8h9vrHfVFFm2wWuSCEvpMRzChF1RdmnZVWsY7Pv5/IKFy5enK1rnq1mJj1
tyuSGmqnBOUB90WRrTFtlfGn0KIM2tBczHLEEQb7rhVEfi1cfAc3+bcuSl3ns8YDIApU9xUX9tM9
yqDwsESyeE/CU01Cl/jJWhzIq2glrYDZ+O+1HV905Nuja8TcGP7vyUGVxgDG/LW3ERHhhbbhUQWt
/GPJqJq8fyZ2H8dVMF6inpfGvTy59TarKZT4/sRmp1LorljNcy4IGZ0uA31yeY8EJG4S3M81QAWc
T3N+j7EToRyuyBwMK37FCnssFBbPFVA0k6Tg0BMzRH5m/qauA15D/tCCD4KPohLRHlxQTiluy9LE
KL4H0i/orWI4uR9WoUcjPl1h+bKuWND3atFXcpVzp3f/YRZqAqi6gbBxM7OFA4l4z+3OBGCcR1a8
6P16qdW5ZDLmBOCNWaZkwjV7U60oPn1Ccmmx2U3J9dXkw3WamLsy/1ZGcfvew/AqM8ms2ND1XA6K
vx7+eUCraRdowxxjIEnjx8iUmmZnmLW037U+20WhSMOHr3lPxgshT5fGgYgnrNV0Aur3Tt3Hqcbt
44uHQNs6TbYGbk4b6muxV0/P0Pj32pd9GOHmuEx08UiuWJ2utF90LOepuivKefqv06CeD/gAaMFS
71+iv7Pmrsb8CT/wrWm7P6lMukAkLGYD+WrCY8zOggxsaKrxi8SM7XrwwuH8ZKPv2B0f8wJXTM0I
DU73De3rNmQ7LkENEaknpnGigN47GtjKDn2QSjSJ30CrtDbwbuBLEQo2mctyIIUTcHQ3KToCLHXq
VaqxZ6dFThfFJ2xoH8+pLsp71fnOxN3rvsschpVMA0teW15ho76yBnaUEDY3OeaCe9JC3hE7x7Ih
KUaPoOyPpK724VnUuCdg0Eh6qEsSyk6IoNUHyjC7tKwE1w6POwdfaYGWBNO+lIdhamw1azcZB4BO
QKo/Ybeooeza2oi033MKbK+z0SU70f3DGAKNEFDWqzmmmFedH+51IKp3xqnGsQtTMsarTlN5HqYt
fhDmlB/6mYggh8i5G2Yo078FyfAGhdi/2nMiAHerp+eCUIsTBRJAJJ2PNgV1pVIRiockSrzpOf1i
vQJHt2Ga+WFTbWgwbujGDONTGFtU0Bj9At0dN6o86UcapEH0xgnqyNTum9i2BlzJ5rbNteZKIlX4
ihXKzBjpLj5gP34sm7Qb974WfGC+vkZU2pYuqMmQUlTqWTdZWAPHXIIg3NSZlkDltbwxESVmSjpD
sPQ3f2uu3uJJZXD6+QIZ0R0TI8bXhk0EgU7j9yZL0fiojANM/sxOLrdbU2IcivyAFr+6QslV3MWj
zrM4yX1nT8I5cIqBXGft1FT4AUW7a5vit6IWXR+KUaHvI85numpSSUFdwM7DhFBC/MSBXiuXBwgZ
H5wgGoTzDAj6cm+ZLJ30wSUxrWJ2U7rR2EscrWTH668SQ8yDHUtB0SDJDTJJhx5Lny1+QflyCJUQ
bHL6KaXIsdNjAVnpZa1incNqRDF6NL5EebAcIY6g+jg/PhBokvfw7cbU5W7/KAJPACDC+EgdV3kU
ZFBERQzM657xqxxIl/anPAaTzL5SjNbL6n9qTzOovJvRfKg33E1fnnLx8QyF1hfXdGKSxe3h6ul1
vSP2XVZnUY3GWNSan0ID2/1G6mcMpa8EhTEvUa+OAOoA3vufy/0CbEG5pRspul4ijGK8M1GoH5EW
ITIyrH1Ag1q/CMBWivhTOzh7TvfJEDfrlUOF5FopXu4dGLXgS05mga+Ant2xC5vjFuX9EIc37kVx
hHZ/mWwERUHXhZlIQqdxvhgZwF55Dv/lSXmCSCw4r2OFQ+FqvL1TKZftDVyJW01n1khzr5mqllxW
ZZFVc7p8Gl9mXOmEMK3vjKkPscPFyCvCVgnuxJFv2b0zyinRW+hWcqTEI/U83a4NBwq3DJxLw51V
3zlA9uQRC6kREqW5uSXwgc9Fb+tt6HtNyEGw5jzhR8Rs/KKwyx4kOqFx45Kqg5dIiikBsYTtaRyy
BRhP0Toynl/bL9jhZSfjLDyX1tkKKIZn6ZXSwsTPi7T4ebYdc4myJef+aUEqwgYys0cmdhgG0n2/
UoXgiE+uDtHORCFiT03BWH3cJTj3kzmIpokBYTZTaFdvn3epVWpBjlascfBdlM2gOVW40ABJLnLM
SwBLfIHGdC+NVnSn0VF1FfwYCmtkNGYtn8nNfVVTw9/yujDWN5wyhX5Bo+syytfLQ2/aoU0y2Wlx
HWVf1Q1uYk9jnFN8nhas68XPTQ/kY9ByQZ30debPPn144/cCDl52y5Nvs1x6Z009nsxmRJ/GfTRn
kKQf663YJb4pv8jgZI8F5RfyVPlzc4tgVb9WN7+AN2iANDHFcEkPRoORpHGTsvl67JnYt9R7C7QY
XAftlb5diLD6TYEcwW0dUec2kMdsugo+u3PBNwdnhi/WFbFXFSGQ37Jco/JRPA22AuvNDxnu8eyr
BOmtsDGULMkVliDKbVHp008YvaB70J+lJA4Rj8WO74DTlXPanOkrkwismB7TEJI7PtPTVpHgt5WR
xMo2aTA4JK/Pg4luxbbMRNhxJGgu/D8hFCn/a3Y5v9IBRAdpxgxAJVEIzBUuVna1+DUdEBBMy4g1
/PwmvxdP088EmaGrrXZZBEohCoas8LdBSC39Jq9BEix9OrwCViP6QZMv58zLCe4uEnQtHiZZBsoW
rLCSXDk1FIklSIza3tKigrqPzQU/tY4h8d/t3+xqugRZV60HzWgcLVtr1rgwlnm1suZu56TpYTRs
naINfsc5GNaFpaXupv5gHASHoKcxhIkx9ZHY4NWcFWG2ca8QBp8TAaimwGIMzy/1ppXbob/qyhK+
uvSgEQ2Vbl4B3/QusUnVECQXtVuG1g6OzRrCowRjrEgxiyMWqavW6QQ4P5IzQkgs+cB8Ttp6ftxw
0C8JU4VLVmr+z8IjJwa0oaz3SVATY/dCjNyiAdltBWcy7vLI9rfeVSWeGziAduzghrmuxX1o+Vte
V+9OB4gdunMkp35OUtgj7cRZr4RzYIJk4SHdQBap4QOr/aYv9oXVPw6CVU9avg3+N/6vCwYGC44z
rJJv3AOSSlyHdpDlwUrXpP4V5ePgkpC/TnzKKqM4hH8xYXVHJKE8LFgV3kHrpohfj/rBtYy2+a7+
ZILe3WsKnLb5qKk+/S4BMD8fM1/P2mTtSNjyeUyCyVT2lUbvYBw1BMLRFiFW26PksIPv4oO3b92Y
xbknV+qePdJ12QbokQb8NQvHeuae9IVvyqh6VIDwE2QIhlgZTTXOahlhzYcyVQIbqmOnXuGULHEW
otEbvjI+Ven/TtNE7DfKBrQD++lo5Wzmoc7tsSeYN9YpCmskTkAg28RzzNQNzo7abQLNMdNfdm2C
qYTWjZ0vSpryNa3enrYN/kCejuObkQSqy/QYEPC23p1l76zvdf0vYwKHzDuuzb6xPOLLu9VxoBUK
pmktkZcWwN4hcmnK4LBExiD/lFPyyZ3Piq5K27PvBA77KEULHfPUFe1DQ4WHLaUP39zhCHKMEDMw
xCCtCf1cAZdjWAzFUbQg2LIBdK3CyxZo9BuHotpUuVBez83tDeiYOoJq3/fKxsnjDOcN1a1aS9K/
MgURElibfGVD1RE7+p7M7iknGwJjAtfkMfVFhhuUfsqwfD48RGVU3ubN1u5Gx+js3ZDhNb2atQtr
QGup1u6w6bYq2o0Bq4pKF0TLJIYuf/mg7xTBsqpcUMK5Og0hf42t2PMv6MFHSTSpZZ401jj98b2b
HNoxYYQ5+FrnLIKLCOv7OLHPtzQA0Zxu7ZkqaYdMia+E4wXcUB34fRof/LhzFavBgHL9HHExaILU
5OJE7gY5PpBuWsCF96oc6IkRPa/J+whRwaXStIoQKOZOPBQPSAZKGVn+7uzf9A9pGL5FAzkLjEXy
3AbrDTqSpWN7W6Va2QT8PAPlvQdugcjQa8DTDDwnCVPEKaCU0DKx5ETlbdC79OYGfTVpT7bKiybS
70xdo4NfE5c8+phYVLE1R1a4q0Jklr7FyEO2Rm82wr0v2XI/f0mnrF0B34DQIcO0y7SjtCiaXano
7vzUH1X/FYarCfGwvMc8bzdEKQvbWPtaAoeJZWBOU+yY46vhKRABBYohpYFyt+x4FuyvmKhjY6h1
gN6HSIPGqL3+g9UWP8w68K1+UuxqVOnk+GHzYJR7mzgazikaYfxpT9+R/WYmvEuDGzmwGqDbRdbU
278NxA3zq0D6gjGsYxGpeezJfLqQruU7qr1QjBOMTZSmadPieCqPK93KlFEWTRd/VwD80j6fXzO2
nnPli+0OGDcYMUNjpBwzOQ7Tbu+ixV33MUCeuxW5hkFzWPM1YcsrMBlyMfU+9yA/+ZxyCbaiEQw4
3fwmBG3mG6nDpa9o6Tnd74Dye51GgjGSHZ7Fctu444RvMWtZqwwFc3xX6KxXNjmzzLJmcFJRjzFg
mVmZK0d6pO2yPRhuZZiOrSCmH/AiE0doHSuwJdaE9GY8CiLjumUfQr02H2iB69x+37UGhuGnCjdW
y2FP5zvxLGB5QMQe0p1/FRywpj5NAkTvPFrGYmhqewUF49xRYjK7C6BXGrPcFSN9kB+xk0hPscCA
5T2JlwkKyU4/4SOTjF+G2rtpuvaahSjvIFtbZp0mJ5myQWyx2LQZeCioy7MILqLB6GsuuVWgEhpE
Etgk9Snxy2LQ6BPnA/pd2QvYskqn2c7avia9dqiyRkK++g4QF+0+mq+A7t/focR7cKriyB1IYd9v
gOA4ccur4ARR99w1FPf9B9XHU6iyWZrF0pBLZLf2LkgVbiQ34cRYbwmtv0xkbFhUEwS3qXNRjRJT
zZwzaPRIXqzQ1Bsg/eIcjV7tBglafd0s+ukBCHpE+RLjTRPy4Zj+dCKic7AdIQS6/Qf/jA/2cUPS
nUTG9B/9s7gIt63cQCZNdCBNzED4AIw5ZZ3eQP0d5ijcpWbN93g0t6X7xgtmvVwTTGe+4dhGgQeZ
c5Q3RMzxkQ57nveP5xjVa0Xxq17Sygn3Pdx0ckdzsyKeh6aL6IRejc/HjyfkoYW0nrEKeVwNYGgU
xc+4kgauCz6VcD228PrJ48T2VEEmbiwx041IQcAQvpT/4UeeVhRwWSA2fIuIrBN/wNAO9i/B//FS
mxm3mylm3zB8YsqIS5IFQznQQ1QHpQJ528G4I247NKG1UGJDY/3Q3OPBVlO/oKiMtiKd7J7j+PLk
vnWAveY9mg8gzHdvcEkMAZls/5etrrpB5z1zdhJel0lTxDmLLJEsYNdbGAH1D/uisxbvDJsODn6u
2kfV6juvk3uMNOzrdMDbi6xCY+I9KIy4sCTroBWwJYJjE91GyXeFoTb2NnzHq2v+gDv0DQThrz5y
+bFUCV4bayECpOSD1rz4uoUOloFhZUQGi/IZghGf7UNqQ6Ic4sSWtnFrLHXEVkjQ788rXhhEl1qc
WF0dhvbF/g7kpcsgcFYgvkdy/c6fSUktd/0mekl7FUwQ6e08LQs+cCxmViaDxCJ3kNU4qze7QXmc
Gl8TiQOHos8HesZr3HCnpofCI2QVXyrzjBG2ZqVN9cCMRGCUuYyUNQUljFj6OuhKRaYI8alIy+l4
JnvX5loKpZG7XkcT7+/p5YDAdb1IEHMTE3bcDGq4S9S7B2LIdRnIynOwS8qctRi9XUEjm853UQ2S
prqAWWM+fexaZFkFu0E4KYQN9i9xL7AuSfS2aQLSlH3YM/EjPyJxIvG4VDDJzJ7vgh0qgOZYgcf0
Ckbkmu/u78z5yJ5iMKhp55MXZ14a+YLyqWm/G4awfTLtZKgzeNbzPJAHMq6jWUjM8kUQiytDFjC2
+1K/vJUkb7FA7muVmzkvSaNppw1uRsWQbSZCBf8SoW7vw+DHmRlkU0y2YvHsz2z0FKZ4dbX7z9WF
82CtB9bWL33t43t7Ilo8MX18vKWCzDOOHgh8undQA/oOV+BNtbFONSNlyIz0TKiH9VLL18Ft27FS
eMlqdXhEYLJ9vqT1NOlRj0Ysb5Qt2RLqWauKklU3q+GH2YnJnfcPpTls5QA1DbNBblom5pknSayz
ue2JAHoj9wVFgfVdDBG8GsRDHKLjf+FbJ4mYM/kFJEnHjP/o80pNyVhMgTt9uTdFgZXTSVKzMP45
uSU0LqveBiJP6e4CJVXiABlg9ZcX8RCAt4vBWtnONyr9Wj4VE4vDxeF2/Xqbpm27TJoDgDXYdrdZ
RQ2Q1WbqPO4+69G4u57Uw0wM4x6CIB050ThPs5bKC4QRCiJkmWy3Kiegag3M4BZN9TmY0D2/3shj
LJHk3MO+fgIJ/+QxaTb2tkOREI+h8k7Qbo3ClT2+0/36CEc71/zBYHTNJFxpHiHoD53mrOwuzmfb
Rpf0Qsggv42DlsGv42svjW5U9f081GB6NAjCa4Y9FetmSBI3o90tC2i+8IGdcmJdqYAYdr+dShIA
fM5c5GuP3v4MjSRrlwHym2SavoBIWi9sr1SnpwWPGK7nGGjZhCuYiyBVWbJ+vLxbWBaSeNrK3QMu
7tTzHoWQVw3JoxTGf/tqA426CPjr8Rld6qbkVpY8usax74lVEl3pcw+s9c3+ai+0ai7NK/+J2rjq
iYUTQKmzzx5vRkOSD4+mGiMLYp8e/rTEiZ51q5vze0lhGflN9w/XTaLVSNqoX6/F3Hg4TJqGE6Bw
k0vVyGfTMAbwwuW960+wpXHekuagVFQ9bxLQnxbSxBg9ku0Wha2dd7DsUC9pbGGmXL8232jaP58B
rjIA6RUmPQwsKWcEs1yZWzu9DU5FpsBgCphTbplJxSFmtYSL8o5WIzHeottdrxf2oBTXvi8WxSvg
NC0c53LWa3E51FaY3jyz/7vkzIt9JgVs/28WF2qpf/9YuxrS9B+fLurEJiKUOs2KsIlb47vgOZdB
m2u/va1M34rO2YiYWxlZSZuCxd5+6QkYVlhJaeH3DsWhm+pk0FMl3vO0atcylhY4YVobiDWCw6MS
yhcZEN2H5iWwXARb3BPVJlXOIHlajrvwws2KOeCCA1DjTbaPWocd7vtROdBgmwbSOcR58lJ9pGTX
IcKbhVVOas2ve0LdvXZggkSL0MXT/eKDBeFJ9S2x9IEV9Nu6ixB+FKRViugZG4kt1wMGb55NP8Da
FYs1g6LLUZuy1UNbqCvFmW8SRdgttLgbt08TT+rgk3ZXYCCfSeIMFfP9PNqoCs2QwkRzKvbtvR80
v2EP4reJjZ90wOKjCohWJuFbvPUL/7UIyJfeAa/unTpkOvYfoAPAIrTmhxbgKc1pelXUy36DTpu1
TOSc4ol3GXsJpwP5RGvdaF6xIXb+v/Xfhf0tTeezpf0476nwDfZuEj/0WKQKH6Uun17emJrBPlCT
WTSVk2GQvvon3u7gcmqkayhrpvzevOJgTaKFbykLJwMvJUC8EXTEBOO0zBkGpSGi4Jct/QKUE7HV
0fvYJLN0MLI2ipAwCFSZ6SqkPMZ4lJmaOryNRkOI8aX0vB+uk0U+zRzOBxfB628fDYY6owA+4ez0
BsjO4j9rX2GZN1FK/p+pkTlcC4cWNOyzBYmLbdN3pAzWODGJZUX8cMSCH5g7ptky5JloKlRzZKq4
D2P2S5aAK9AjS+cNXUaRUTUPZ8YJDv709RfU6PcEaWdOgrKyxJztT4a8aabjvw2GT5AG3BBheRTu
dtH+1k5g6p2sdhTn+96dax1ZQNxezOU6BCVk+9d0l1nGnYnURBoaAJwjudMR9LpwTQKsqMUWJdBh
ifiCEcqQxX2IqihQb7KqyynM2gMIBB2dWAd2AG5F7j/P9H2a5rQEXoWYnvQLS5EMmVPHGXMLW/Wb
BDRtJ18+QEsvTMQJxuy0BVFbk9y+6B0YhQDwEhpzF/4uM2Dgsc7tGuuIUbG7SMnDXf9Ij5bC77ge
LC7u7hTqTtZ4Lw4AZrXjjMdswuCvOXsIMMmhL/0+pr39aoJ78jg2EbaXP7rjl5pZtNjMAjKszko2
AwOWiP/hrmuBKh0z9ZU+JoQp1GjkjfC2acEOmYPXV7ai4cT7PCLuWvOtgZRAHw7hQ+H61MhnafQd
A9XfslgadO4wO4ksi1fyjnfmBxezB59mv19OkRU79tE6LYIDg76Vj1GsnzaZOY2/phQkVgx5yxQh
E2yATkymAcVt+rTWgWw30DPzsFXMqdjcNcXnYrK6cQu94/kyQgP9CF/7TnFghPQXzrU5pOPz4EU1
YrUFSDyyGBXEkOE7lJmGxua+41acZC2HpzNt3Hl4KohQiwqtbDelik1v1PwvyMViOR2G4GOdWcr8
xhS/6Uijb8KOcYq9/VBpjo2QY71IpwEYXhFs6FY+U+SK+A6l9CUbZqy2C0MIu1eLkZReSKZ66UK8
69in6NopiUFAZQaUS1uCE6Uo1tcfr8fkLKI5aZ4Mw0QTgT7OJ7K5Yxm1o9rcpA5OivFjOQzYMXJi
GYf32IcQVqn3nV2fTcMJsPCGxOnbemOMlW5xiuJtMKAw+Gk5Jem+w3/89mJSRQ4mhhYl5axdwOYT
LkZfBPgSfuxvOWYmXieLY2Zn9qvJlgzKBzrjv1trdxdNiBbNZNK8RK7ff1MhMDQJ+CM4Y04YkxeJ
DS8NVghanB3e2a+sMyrrESDPuLkknGrtfRM5pnWngoEiHvwynykNSo4YdxwUEetHIjMA0v/rH/do
r9kE9lwOi+RFbOq0WWCnflFkHUmTIXMVbmQ+MMxSYA6SfQkrqYiXDbw/4nXSrXQ6zPC76APOczBL
4v6026DBJYZ7AG3l95V8HfQ1OtEOM4tYPqYcpLOBpv5U+r7fx2Ac+S0Jhr9DVKC2j6NlPW3obVOj
b0e0gnsQVJN4n30A/2BERlMvv/eCMD0SqagAvqtMZkYwwTIG4pv6gql+kqiCRRR0NzptX8ghAWdj
C1sRrlN/204zm3XbQ9yQnlh0Y1dBEn6i40A4jigRU1b6zqU9/ggxds2pyGxhDlSDcMqbQ8kS6HRH
VoYp0VPbO2NDtATtTYFBzR85GBmZC4tWGkGk+J0K+oCmG6hNIZ+qr9OEIwf4b4EQzHts5GppTBdT
1LyyPCS/8JEdVzitTO4JkrlYm4seiCx7BA79B2VFMuC/zbi2qAEqS0N/OrmVbqNJztuOoeTexkj+
F5myqZAigMlgscWo2asoBxISQxEhfaGHYr15zvfkH8yvyqjrJhIkCzYFOekMV0u/+jCWyRciJlPg
t/arcHwhFBvGnkVtWFLFNfh044nRTzIulvB2bRuIvkahdqt/WcP/0ynUX9MtEVVdXqFkfUro82/6
oVlPzQlOhgKkSNsnqcmwzfLOy3wTXNCBfbNM6V8J5caN/3zuq45cKwuAOKfMHD1ED2ctDqh2L3jt
U60MzyDwGSdyEIyPZyRn9oIqpAbExUYm/pQr5P3PSQ589PrqAHW1rMZ5f739+abdOgPjB37mwY4L
1JPC6sjvYb+kndqAH+VkXnlIA4piADBXdxRIhZ4WpewrILk//dQLTC7x1LVeF447/ntCP9Nehsou
TddpWPFEM11+CACJe5m/KS01iFMwAEN0LpcLz7HoGcGQAWMcbuAlHv1zgb8e8XwL4JR4fH6MrIAw
GdTydr5WHL2Lbjiu0lzDE64dDNWqaiAedW85iEQM1qULwAezbzZoindoN2kVRLT/fjfpbkjF5FVn
BlttyFi+QhvbnZ+WyR9XJOlGs0K3RMfxgkHe+IUjjb+fJejzl1YmZvsCvR5TGJuOO6sP3vVnqZBA
tokxA9HM4P+cnPyeV8ii462rTzj+CQ+CJ68dmQqZL0v/xKruSsNdQRsTC9CJo/Z+I/hTY01No03B
GC5QhHvQhVCDAESfkVaszWku4ndhZxWAysPewdR/RvsRbq9w6HS/9ZX3FnPH6WJ/dSJk1eb8tUTF
73XsCb68Keb5MMDOHxv5jiZzGFsU90C3xDJNXyB9xmgtOK8rrNHjmHNsmIX5sHbmZ+cHS7Cjq490
1JnFNdQxyI1SPAoEyfPEupVteGwjn7xUdxmPUyamRUHkvEEYgFdHRfy9hz7M1wHcTEKyDXQzZPFD
u+bdCRLgV8YnI6GeONfGr87VHBa6BpXhXZMOoL8tJR/xS+qPRmdYkyrFoSOfeSByf6iLAcuzC2Fz
Mnuig9XcC77J9mTxArI1Atqllhi2B0+mM08YrzeSYMuu8C3vgYkeOJdrWOTUEua1raoHKXGuJaJc
Eg5Gmn2lsInzZKjrZEGMj3wwOz6ncQbJyVk5c+haqDqRZB2wHZjJV8+wWfNQFbTnjm26+U7/t85N
Ypcr4PbNVKaZo70ROPmTDhmtJmUOAw3pxCp0W9vnWc2q/9h96c8qYlh/MTvVaYj2o53q0IMQOznj
/+Izp8Sl1OtDbKICACIvvcj/BF3ZJ2+N2JEfy0tBxUc9SmNZqR1rRU4PIcww7UVLL88acw3LsYX3
Vd6Us+LtaTUw5jJoa36EOApH2oNBhzyCZc2OHWkg880KJZ7nESXwY1iYBxhG/fkk9Iq3+Aka6KrN
lkuhy1xoZho6HIpIVgciijpoObO8pfruZK8YQUMWarq46bSc73E+Nldf/HCPp67lzwq188HOCqkc
jR+QBMJIepLk5IVzqAaFNfyUV18+qddWH0nKnpgC1Q1wlFvl1eZ6q1bO0fiWuxCCbkKI6JIcmg67
jIi5OCAZlcneWjxxHczVX/pcnCP2YTgSboK5JZSyMI2LYXIPuvdcw5jW/Ty7VApykpd3ojQBwE14
K1KPm8+II08N5DBQIPBsToSuuHU0FRAY7Qib+KAxcCkxFFp2T60w8lsAQ0lh/7iZQv6IuXQdZTQt
/BDaEmRTK+1+WS33RGAYHziTa2O554cohiRJuytFUqKBJwEbU4C8l0A7fy2DfBc8IvOjppgfOepU
GGdLyRezh2wsBbeg1t3lskPP5y+7uWSlWfgJAIBvJaWMW8Dcydq0/Z0ap0RfPgenqSvKdmJKslET
u1tb0XV0IQfa1s9n3UMzS0XEtKhC2yUbTQuLxmTIh7MC4b4e/CPZZcQLYJF7Y1hKiXdLBIcPhQyv
UrA/R/52VU/+/nN45Tv0zUamSPwZYzgbVhorJfZjMLp0+8wCw0mHrvvNAExfiP/C1fYzpbj5RPKD
VxFHYf5y8AZRJ+bbvd3VQ1HaBey+rgCog5cKiMYqvnIOFzayqXT3YYhbfrWm4iYIcYXecssJtAUs
KJUFcZltZsNKOSbwy++u2ETwJSzNAZtjHTZYWobgeyHjSOmyZ6x1ETy0LNjFGZIY86vOJwU2Hzkg
TQeSl/Qd2UwWsR1L/lFE3QoSYIfKhXWjyfz+HYgmG8q4cslhml+UNFIdgEuxyV3GqmF24noTlrr3
DDw9GM2NorZCnwBn7Ux5IONFDq3P2aXD4xH8CZjU/HzcSp3A+lkLGnbfAPRO7YndCRemAXeSSAmH
LEUrlsMqB5qHsrvbq1GH4pYl1IKWmt+O5MDakn+2ITuyV5LBDbRlJ9coOsD3nhLnAjMSqh6sz40P
2YYfkHHLLPABj/X8FU85pmQy6jZ9o4tXIBB1DMdn7gSq+iqMqmFUyJC7W76FLszvXskojj1iQ6gu
VKsN405vVJB0t6Kchd2PSMVvi6snmStIqJ861B/xHzZI41W8VDsi3LpR9Suf/paMF7bAlhna+2FO
cmM2Fe/P7AinnGw+Ezj2G/b3kR04C0sZoQ9mF6oM68xdIrNc50+zIFeTmZRJ0GW7JCJc8XWdFMQr
qXe2aDXLbZ2OF1zEBFN7Mv1DYE3l3d8S2xQcackSR+BfkdvLVFYyj/SsKCJ01WW34X7aoEAhDNL+
IdaORN4CA3lTaORj9JlOd0ghu7fOKyyh0wi+I+Q/e3KwsaDiKmPayzoAsZB331vy6AiNjTpBgrKW
7AWFESBZJpWQqzjy77O8/Uq80P8Nz4x3FSF19LB6HTp2iZR53za8jD1bNQoEJA1608mQ4hHAfoQV
xFqgE40QkFhdvDY16preMi5JCpnDc/1zGdJ+Rkblmq5Ly75CKxJqWXbYCb/cFOVPF8ItNdveveRG
t963+GbQFbaA6Vv6C/ZWlI26FoD6itOPuSOpzhDJwVWPhTVjHOsGt5WEk0L+QsKbI/nkbLy8KMA3
xb0gKgm7g5XJCY+aUA4JKibMRCA4UXogtcFExnecGAxC5AUFIyZOplvuGBXA7mz20kBUYRc/rzYB
OQDsD4vPCnJ28rIm6IATRETRfgngG7lZp2DVhWLWKmh2bmRI402L7cATfng7cdigyHTpzx3Rlc++
rlbbMRfwduKSofhGdpXspTGjGYslc1ORmXOk4l1C5faXomn2VHAlQMKY/6xI6C1cxYVA2iOCZ+YZ
oKU9U3MIYpl/aiaspQso1s1wuPl1bwA4YPwaF91nYTb4QkAXBTA9KcAtiWr9MyKbjaF+G7MhubJ+
/KHPcKbg7bwgwIoRkjayD972Pc+MFHp3tX8+LdL+ULaW513KRsMExxjVxvLPTwcVBC5D1MsFBRWT
aSariDM/eT4L/+BmosGQ/vj1wWZtG2dkEtbZTbr6jsqLHPNLJBVBaD3jxrMu1YkC9szOaZvP6N7H
Oekt0tbXs1/ezgYCEv3NIfv6OMx22rziRt5wDzF1HDGPGAWm8vpK5D1v+u8d6au0qrQvTy/JHnsj
Jlz5G8wjNhZfZcZsr/WdC9z4GOsjXo79I7tiXfwxCHT19nL0LE0Tw3HvKWeoYo1x/+ZqeY+ViJFE
r0+gBS0VJvhB1SgKZL/Wm33GCiy9CDsTHSR1cPyggTGiyd79ZSF5USBQCk8Mv+NkFFYJAzW+usWS
CTuYswG/rfnoDw2YvXka3wuaQz/9nlCfO514+T8M6UD4rMfanB8Htf3FbvYb+GSZ3XfpX2d3MCh5
Ku9VymdSi7a0W1TgjBVbzwi8rpKG9TYA+l09aOP8RGK+til0wcEmxMgY8J88tEEpiDBEo8LI2QW/
8VIHQb2uU+1UvVeBNAd6u/pfo1CwHSXC66CSMMd3hnVakpNhBXI7MKEXCc3ZIuWlNJmi4IOI9Uyh
anz5/XZCvApnZZ3I6Qz3aChK0KFAGp2w79cQkQDazZ3Bo48VzfofLE/Abty+MC2U+vRih/xC+Jej
0qUMOzx1EV94g7xKCngFf6l/BpN9aKGJBgm/fmnU9vSU7GFO45LGtJ1gISqesXrQlhjqpAdqlprE
8ruQ2riUrZBDYTi+rCYRaGcAsXF+5Ccc3ZcDL9B8N+iOfO3F4HXfchskW4zyEapDEmwFJox3g3j3
DFnDIqtKbcPVICMPYtNlEF0wPmeeDWb+9d8/YxMSRLysKnmHIxzPBs2gVVf7fOYT76G4LaDHIgxl
QbDJfneR0cvgO/hcPwj8tHnQicso8iyULyypmaYixpBUoWfT9Kw1MUOsM3zwAMaTrAJhTqIrruls
A3qqHRWkbviyqN+bDDqTGOspC8E1Jo8lUMAFm6DP/Ci3iD6QT2k5XQOI1XtTnKYAvyzCsXOXgq41
amutzSQsdBbPeKPdEdSj4EZyjaser7VQSUqcHE3vcWURbyamTOmesXFKfG0DZX2D0Fh2AwiJW40Z
xouPtQ0tiwAUOCfInGHk0Mo2FQ6cC9lIZezpbw1msvWEDWDIJaJXJeCe6sa1x1SCN0zplZmL73EE
kNrRbRAaXSo6JrUGL9Bt3wHfdW92BohfqMKBEGZ4hO7fOw0UWCsQc2uvEYdQeIQWV53BaDVHkJLA
cdbl5SxBZWG8piuBr/8L3uZsMHbc0SZMi2Dsi5TECerrG/W6e20AJ6lKP7QUsON2tO4c3ayqOBzm
Fwt14otQJO57aLFeXn3j0IBPU6ZRDqlICDc2JCHqI6iQXYI3BBTXhwJq7d9YwBuTk4fWDJafOm/Y
tYPWFBsbGFAyfkVLVQKoJCy3VwbwjMcHHk+YH2tTfo4LOEl55ivCmPDRsVIiTnOd+1KLbFKs4IwT
l+1Qi/PLvgehvaoxo27XysfqB/Xrqya6XBkoQVydMLPg9KJplywdRKEblLiV7WBW9AYAPvfHSRbP
TicAQasuj8YAtRT6CgqcU9KRck6ZEa8l8RKSai/WOCC11IircuUPaHOs8ISWnbMgU/fLZbFpKBZv
3ExY9Kp27fUm0Rf05L3xbXlcQAFmt9dt6Jv8MjVFZG9YhUL8qnMeOJk8yfw6WIV/1WF3T5qn+9DL
DRqzlptnAURy3uR7JSs8gAOWnTgweALqpisJzSdIvPFtXXFLu+hCf1rB54mCpC0EWKPvDDj8isew
9TZw2QEn9FNGsUJ6MEhyGf/9rtGrQAbDkUe7KhV6s9LvqE2fH9z8QklREs+yzeTgFLLIcyA0uJ1K
/GbX41Jp1nIN5X+Zz2TNo7xqE2rUGA6W/WSdqZQcVf2eZLtONn3drCNJBc6W+WcLgQtGDG5hU3gt
gSkfWSw9n01G0paiIjTFZjVBbqokhMIG+EU8nLFeo5HqDKU07u6ujC5V6WFk69gZrge+C5cTC0xA
gwl7yaBeelnZQ3/6DS0UaieEBNJ+CvNa5PLziUnmV/PFmY+N0YB4YZCRvc/s4xFPctoZmdQ4bLTm
B/yVWKzRtEL6G7c7CouuPoGQU4AoajE9E54EGwwGYCjm1yI5moM0W8tRWePAnAM3Mb1j2IDjDIFQ
owmCLT2Lw53CU47EcydsqE0CfS04o26qb9PZGRUSyVlq5zDllvVqCgI5TbVX9VH26vtziFFPC6Xm
8lAxg/+0DZES7zcV/tOwU37nazos7cPhSUHqFs00sf4tUDhfHidhIYEe8XGbLKsrRgYVDrQyVWu2
HCl7mn6BqU0J0zJDxVR02Hh8bHXQXn2aBPOX+o4gyxYmZl9f4I01aYbgLGC8pfiW914FLuDeVRPs
AbzlNRdSu9qv87kA1kyb2QyryRhQKfmNs0jD/ALkyaiDD5IWhqLQyxPBYVZ0v2Jc77Gk5g2/nhIR
zH8u+uJL60DT24DvaI9XzACmpFGkr6myK+2hFXYlhRaYKcM1VJemGLdwVeUzdqnmyN6s7+ImRM3Q
/NXbw7C/bxRVOEn3BEdi6D1Wnq7IHKroQqK67JUvxJYHvk2E0ZXmhxXDjGmN3DUL6AWn07Rj3oZY
PIgGVlbzFA/OfL+Wou92RGz8KjulOubjh1mmJ5rLzTuYdfaYTnfAmFdTzOppzK2C+UphLf1Ou+F8
BR4pccdYws6LM03x//hcJrSP0f9cHVE8U+LaV5Hhd4wGjF4rUwWs5cMRpSORmgilc2fFDacajjqC
3maR6NHMXWHT2sg097aP5KWuGxMCU0eAlHcXdcDOXizG/Igo6+bwLeamXNCD7qNLN0uR8FJhKz3p
sfhV+PCedoID9bOGuGkNdleW7AWWrWowdlFXEGI13JNZhtbnPV9ZPH4ba9MZOI4iODLljY3jcepQ
mNWrzOE/EVNws7G4q23rHqsGhk3//Eiw2vtPD2PSNmHG4aDSBUYH3/Vi5I2+Cjm0njdn1i9kZDs8
DENoUmyccufUNqPT+olluJr5TcaZ4gv5U/nwq7FNQtDJaZEhXkz1BwAGiI+aNeNQCjebt1d83VKK
/AVTJFqMcEVLgMu2LXsSAC95QKWVLXgLSbfNRLafr8em9Rat4IX4/hhGqRG6MZBqesnUVxAtC8S2
SFCSLJcYKa7twd6Y4v+7rsbBtzuwZLR+qtp6u1K8RnyiLKfDJHdSWAKXdALMLia4nLEEVaIPHAxj
3nepozNUDBxUmsP9QDZhoMHybiXQsU0NEfpUY6K7+rgNRThhX1rgZ8O3FQWOpWOCBrHcUV2n+Jvw
se8i9yngWrbfiPcs9/MsD3BPqMFXBMB316u+fmIujuhQufxNFY2ye/lwpbOqOHZY+xu5f76W+2bn
pVMPDfF4qktrImQj4qtb0zuygZfYoJGiwHTnCy9/wMoLC4fzweX/peqXn7081ChIh3Ae/k309/WS
O5K23n9xs7PvUssLGNo5v/7b1stbXBqGs+4f0vOeDRYSjNKBW5XzraCLIWpeVC0UZNaR7WACY9ts
vJc4XMh6JG8YavaEq6c9+RiMDUpjIMQDWSUnwlkqS6VlRx59iV6Wkf7sFQIzaB5w/SonKRwpyBgq
YZhzE7/rnceaOUZPzfwDYs9MOWH04PSDcv08JWCf/oh5KujPgcJPC0m54IbEULD2PxcuFqxEODqt
fHCsy2HG6yZHMdMQfxj50QxE9dP8LG2Csm0A/A0Z97ZjATPuLjWuGZHGdCRmITFVrnt6zWxCVq0j
TkrywqUfYYBiJ0mH2PL0uiyw5ythhiYiilpIYtZmwCQOdYyTPWWFjA2sNAVvD/e51nm759JcLenV
vrQtCGI2WC94fLmyp/vUMvPtRgUiJECDRgJw09xxRbC+sZWNqtY7+uDFNwhk3zOIbb2mG1KMwBHq
p9w+m4soMyBick0k7ciGmw5zh4+TnQLZCcy0gpLqXuAOffflpBva3bVPHk5Cx4nyE2hx+MM2S9qa
w0zAH5d0UN5nE2hy0d87STGYym2XPo3DwzImWXqKDziHIVtzxXyEj6jOnBlQT42o5A0xtAjFBRew
5h6aqdEArOZykcvqX9FvdMew6dRSVw+Z3izxrFGnKq8FrFOXdn3iqIbK4Eg6URwY/oy9uZv8gXMA
PFvEHlovCMsV3TSRpdZu5utsa9t5+eHnbWVeZ2WKn3h+Gf+tYA+zsNVpJsfAYHL+OPeCup+QpfYr
rom1mgGl+kaY763WYHhdCaJvum+JWgigah0C4wslV00RL+7+ehGFye5HwOI35rl+M1Jpgm5rDP94
omDYcokm0nl2gHT9IShjsZibujKgzURO2oK2hGtekrq/5b16c460RmnjJuOKOJ5Z6aMJ8JhhAnHi
+p5xuvMNaka4KHdUElc0RO390jCCMs6mW1EFG7rfb3z9pKb0vpAz06SYBFiVDtYFjACxOLzyo46g
crhIsGCydzdojaEfbhdAEUyP3A3sLC/xn5sMEwcyPESn5/6v6hj99gCi9QGQD7xou98KFBc5lhl7
KyWLPZ7L3Z7YuiKO+sInGq5BfINy/WYB0xt0Q1xIKzJeyLRazLYpgniDXjplg1ksV2S14MKLveq/
LmKoPfeh/vLX/+QNNHI3l7TON8I+PECh8kkF13pJPtadfzRcculRvmuBqB0nRBgwP1Zyv0GY9GDs
aldkb6nUqfbJn8gHxoIqYf2LjV30+CBJK7l8bfv645oj0SQLVxQOkyw/wDlslCszX+cTt2NSqfEG
Lo+GBBgxgZWgsjLBpGVELNHN5Vpf/xfbvG/PaA32xAEqqqxVIX0k5Q0fbdXZtXfYaWkEDG6Haf8D
AAE+KIwwW6m57F11IOOidxyPm/0p38zIZg+AL7+6sxmv2c+gnc9oERheiAN8wXTCzpl9fNYO4h9S
4k7JHIsNwgdgZ6ACeHdkRmAASYhSKJ22sAtirH2Uc2WKxUiEqsc0VGgUapViQu2vWsBaiRbTafie
wils6WvjR3Ag65ANpwuXqpZw/5WS7Hh06uk6Zg4RY/DieGBpyZayKKZBLlpM+NZEvSIA0ovSoWJu
c1oZ5LAbHvOXwHNqkT/sdSesJnT+sUQXAhXEG2bdlvyjIZuOuJs4QO0NDTC3oQndpo5K5+hhRsXd
wFDznZ8/PPxREQB+wweGl7cicgWMviKc5YOLRyn0vWRe9MzhAgB9nmewI0Td0MKunojWUiEadIs0
cX47/LLkgBG2ahAEWX7DLDggaJmlN/++mmtn3lgtjejovrvRDy3kEvMNfEeynA488X6jZPsQqNJ9
cQhmqVXxRcul9FoXpjp4037JB0/JpmlblmjyV3bdiCZchz6Z4X0C/gDUOmZSZHqnrTUhglWQ21tL
qUUbgn/yvpzS/ks7mMPIaHYH7BH1bgwWnyty2huImhnF9PsiPFySql9BTRbQI7IRDrZWXNgvjqrQ
RCNJM6GUDG5wxkDkBqYOv0yeMX0QRzEcisxsiErNtEz55RlWyK79znNvOMZGA6yAElWisdKTW5qY
2TKshnmRmXaI1jZqi0gCDNETl2CK5xWv5sc4iS59BCz60KB+xy/uKtz7As8Qm5yHL4UQyW8Z3IuA
8dvFICdlqyTrNMAqlfMQFHi/NhVOCR255hFyJVb+oT0VSPkQAKlB9JGg8iJyitp6KHxwpuVC0o/m
Mf8QDfB59BUMA+myDveo4R7lIYQYHZfV2zRga+qpaOYQCiV1ALEAr4dPZ3JAEMmpnc17UtUd560O
SICvYyF0BirIZWNXF6AgdUrc+g66oul98rOLRC13JBdF5pg2AgHVlRdr1AtDXK4Qjj5PlxiGva8j
2+8NUzhfoDtnVvNN8x5x5kr2viaIpPrsPJyJB23dnCuTFaGUjdix48D+YRMseXP2nBZts0Hvxaba
O4cffwrl9o0bwbwpYwtp4jBNRHfhPwvyhmgVZnWOI1lIxJAxoaPZ/nJF2B7MSZQyv/rHh1BFHpLu
JOInMTrhoLlxTmJp4Dycw6vCFE/XN6krwl07SFDuZSxoAz+KTBbs7tbHS7ayBp+KgxHeCB/bFpFi
QL2HFpj7V+SZavtVBP8IARjw6UYfB3RuqmtkBNTsxkis1IUEVM8bPCpKvGiE7VCwmADDdKGKVRfq
CEjqq18J13ikVE8Vden22awC4v+0ICRm45tEkZuDuQlTduq6wQyhkiiTF8AIgIqtBIKtz3YUS3RA
rjRgv/dpWYL18ZJA3eDJbvpDLbWC7tGhO6wro4YjvDTquzwKsgGWILoCBpWRq9fQx43z8+IvXbcw
04NV9cR6Qr+nOVcAqQn4bUS9BNjBNC4vivEUPkpPKyQeXk+cQB8xx/nppcHnC4rISFOvM1aREIaC
a9xJbXKQHoWXHFFW6r0OAL/l9JyZ+nKWxmCJRaDtRvRActbBm3mlbR+ehM6yWnJLStz6ItExCHPj
VksVVLCtUGNZrz4jIbGDviIAOHPKuRZ5ZrbdvBP5393gt2LlqH6RT8FYttawtBWik7Q/g7gb8H9a
yApZW04x7da55fMGcDEnUoRkOxIZzEwaNv7TIwHbtiED4WQXoPs8Xn3hNS6SfETbZ35m0aMrYLgU
1VnsggnKpxKbJiswwLMNmmbG7qkzMPlOgIwy8g1e1C4JpwW0Dx+5iOPfzK+I8d+AabacYWEvGpGM
W/+5ELRBnwl5H+CMfM0GouiBHM5MTaHCv6AExDbqHZrJJTYj5i6HbtTvgdYAiO0A01COGtkf0FME
37kwKs6ZTwC463upn8AsUrHAdS3AimzKQU5Ixw57d2/FtLYDIJvIM5BWEEp1NlU7ALKCfEpIaBju
KlKgwjV+WY6sDTFCcXQJWkLzvoY9SzuwYKnKpmHSZTvmYrRzBFCjE9N5VLLSS8JMCf4cglCbC+kO
GB4cdTA5VyEQ8VmOYvd8bvSBZUFycEtBguAq7COjtCLM0SvZQDH60Y5s2TJ3G5fyQjG+HOrKwskN
H8Txkvi4hb30pOM7qpoo2usm6iTkx0auu1+DwXlDW312nyWPJxKeT/vYcHrP6/i6Y6k81VfPDS6n
WwxoLySN4HLteRDiGZur9v85WIrhI3v2HtSfc+0Wkn6O6qIAmfpsKZJB+Tq2lBoIkRTzRhUI8oY5
IEkMBm8XbteSQs2wWC86l4ZoCblSxpzh4UyYet3qUSCJ0fbggEwzLlQrTzLhVh5YHgL1JbQRZBXm
LQYW/BjanHK+5/U8JgT7533igyjiDfvs8eCKtH+q/MoVeb6VpHDc+MD4XktvTOP/mNz1ymREba0/
AAbTYjwj7udJ9UTzD83/Dp+Qy21t+3c2zJzror/1sYJq0FRVweqcS0AUwUEFGzkOTM2VqqLzaLOM
kBolgEGUoFA7I5iEOkdtMDHA955ajEs0KDFBWUEKsGQkTy1ktU1mrZO+Qm3jP7SyPIPSGlKsatyq
2OvaxQLEqBOX80MsC1XZebpSsX+CgsSCznn5cdm1TY1D2Dle4gx3ghCMmDKMcM8AZ2ZMrF0vAXr9
7C/OYWMpvzhoHfj16DzeS4hPpDvvSYMekKcWN3tSlm0nOtU0UblkPcGSLB5GhFIKeBPmeU6zdq+K
l6C/veFRk44VjfRBig60H2q62twjsqsq+fub4mFS8KvcBU8gGy011xWjgIavKblqrwVu1D+jKQcM
ofIpD+XJwX6uX9n0JBkuel/OIjpyU8qvbICFIBpL90IEBpVcA/9rLEJhiVgjmlFmriwe9qeXgzaN
k4I7i2yLNHWSxlZgJj6w8kM3Rcb67Mfikx8kW25/z4d1RqJv2xpdA2UVDqKEJw9Pwax/G04veD/c
Y4XnwTRgUKTy4jBG0hDSA+SaCVuKgu6UzYOajq/bTzHo46Vv7OfiL39tFhOMRRmR5B8zWGgOnZoW
t8EGhR0FNfVvQD9UITj869ocxKL94LkIcQtcraqIksLszILCXSXJLJlU7TfJiiP3ExbA+3jAiga8
b8pLpC8380CxiPpMGATU8dptXLzzGOzs89MhZ5eeqtrgXDzxR6z5W3G0r3jjzzj3sYjYJAQc77F+
ny6MEATz7qlfj6Qbg1tMhl7WJG8D6fLsGE5bPFF8r+LRBOCwOoUnRzQNzm3DB414IyA1XL3ky/3G
e3w7krNPq9N9cVzLLSUBntTTsx8aF1PnVjnYhBLoKGuPmojvCHzclDlGfIT4IXybdYlAAa3xl1Zk
9ehNbJJ6FcUCO/HdmfrbaovOkEuzNCKogIAaAgjZQCYQHEt8qJzm1j9j3Tw56QYI0ZhEjgsxlYjF
Ng8E+g4FpoiNDWkILs6I/DI84v+G47uJ0158Z4/781EVhGuy2YOirkpt7VyWIYiExbGYLWSrI10a
mgfCtjJx3WD57gjTXA4WEYFaaJU2YbPsPIkx1jbzPEx0XMjtGQlO6KXYtr7TGn54fB5SLvTHPJmA
jdMdV9MN5uaKzQV6K1DmpTIdHeGIcy/uGUsztd4yWvDUfkiCbZNXUBLkLMgqHHDibiO3urJGUCPk
4iUl0VU4fdPoaZ0vjfxFBe/QjnjYnH7qjT3q731lUarKShPv4KFsO1Ex6Vq/UkNJNKHo9W9amZrl
io6x5NuI/Uan0N5uGN8fyAFtX3A/Cwp9EktnINOXyMVmStCHmgHXtBHE1mUTjNQvd8Nzzy5m/zTk
0IS3N5gqR+bKYzmieNSMe2hL9ve3ioC0SbG52kAmbdL/djY2FdPip1/twg9d21XdG0/ozH1fhxA5
aIY5aP5jn2YCZo4YpNj7zV8kqy0G09GXzOW6qVQCB2oVF3caQJ2fVGi9/GMAVk/pPhnKA253SBpu
5coA8iu5tPnC1Wp/A+I+bJoc4fL9w5jZQoMy/VxzzetqBHi+Xb9EdANiZvJL7gdQe0y8vW23ubLO
62SQ3DYaI0a7hRIjZmQcFbt29X440r/zlkKMMfPSntRpVtJnaiNO9VEOfejJEnspQcjhUqMi9515
+qu+DfbjAmet69b5z5vygc+IsXtXB6Qyp1o4Ix0HeVZZWtNQ5SrxSVic0yN5JXfRap8ylvP2kXtw
bKq9Ei5NL0xRVzaC7xxJfJNkYySIU+FoRCNzCLrvXTs3Dl3FQ2L2mTQ5jk+LydxnEdCgk4EGTO47
7H9ItDI3YBzNnkHfgOwOvlHbcqG51N9VX5nQbMLfS9FBbPC9fkDIpdnkxZj4gUPdCiql+hP1BE71
+0qhaM2WhcvoIk0S1zN7hjfbQAvQh/IuqSv7D+XTaCnMtsZ7mzz3M2l9Rn8FX0KnA3oa+R6hnnWS
2rPxmOWEmPz9IoxLV3GQBr9XvTu6dzp55sCtb2CcMRehChaPIiNz64hoLIFKO5zmy82d1oBCD0Ou
2WSxMB4+CK24CpdAI4eRuIdnTzeDWt6LUc+Cdajq9V6qL8VJMfDso+fsxev3+MowPG8flPx7sm+z
1hTLAXqQGbZYVo2ZglbydeTyP83WvV7aa4ns2CIWe2RK8D3lV2s6YElulyY4MN3eqbw//DuZfJnR
qzcYhgXlGCrxe77M+RgfDVflRGwyjvRVMxSKD35j9FADEdF68Vv5OrJxeIS1RIpqxUrbhfNzBlJC
B0DalJYxjnvUxybqTK1QgfemyM40HUtAdPtLXB6Yk+/e0uUSu8gKDyZFXlDmuGfoLGzSqIx3ILRj
qyieJrfuW8h4k/03LGDHeKbmfEJa21od+PEcXqPJXjTA9X5RTQFSKc1HVSCHWA46+ekBjGpCQS70
scAxA2301AJ1cVjnBXr1Gzg9g9ArxwWqgd5h+mh4GBMrc8gJimp6OzCn/HFq9WrLqa4GG4xkEN4m
G3/nChanzZ1LqS3K2DyOc0I8sTkt+NI479mU6pdxl8wYZP8Dtd4fdRE7I8ih+hISCZX1DVMCFbTj
iQYS4cKDqsuzRqeA8FWyVhRk3IzffS19MAUR7xk3xIU8WyU1ST32ydxlhBMRtRhm+SldoorKtGR1
hZHSklCIOMWs+4qQ3XDgBT18qInxuXyD1MyHvBCf4GLkm3xHoXL3uN727nhk9td5t1nkW1RctnW5
Y4jMyCgpJDdoPGSs+RCiPkdr9SKVA2qXWNqcJIhmL4IZzZA6xHDV0OX3XFHenWLa1WDT8O5YvSaP
vBRYaDUXEwTl+CFl28IhYIN7zEsw8dggbvv4aoXM3Kj8V5B1rOx8NTif0CVNt0OjHNWMoB2Gz6OD
syYEwMZc3NKfAchOJjHu3bz5Kd//PaVjVo5Tf2cw/2ooCGQatBcMBGshm2J/jde2INNDC1kgCS9Z
eggiSpJtzywsnPMkI6pGUIIiOhRkR7bEI3+ynoUC6bGSz+L+yNgGNN7ViR8a+Gj0WKxpsObUr53K
kk9XRMLa4sop6qKhD+tBMeoiBjDZYHIT3o3eivwbH5oAjnEPDqE9idiOa7Ib6WuUJ7Rwc4fHWkwu
hNBMfPeD/N8X0iyTZ+AffGobBYLngpmvHgdDOUL1RGLDhFdfj+7hiKVcRHKTm+suJb2BcFPRmH/x
VkinssGMh1zvK3TBDcsR1DF9hGWPeMITNsESLNIDN3rSffcBI264pHAcKP4BeOgu7V/gPRgbHQMc
dtt3kae/CVDh0ReaSM0txdgwkuN9KpgvUsEuA2C6pSNN/IuEwxOCX5AfID/qlwq+txUCLfvpxlJ7
ly9LeleeUDkBIn/poznUexpwQZXqr7SvMYDP/uXn/dxyA+yJGoz0s23PwqwnOP6tshuTXaQnd6AP
f1BaO+71bhiQgJj3YDyFD561m8SwOzJvdbKw2i3S/UMwIJRzmAkT0ZYyqxfte0vwsRRivUaXCBlH
fNfrkY+0/jhVILogBc89CYD1ZV7N35+lY5hkYQf6x0RVh42vGxTgBij7QPKij7Lswv7E0pXF9/T1
cX70Qd31MPYW7xyoc1pLJy+cGYYYmc8KZRE5Kdy5HLZtfXhD+2Iyxkc9efX4hcyI9t/yc3fnuWgC
iz5KAEw1cHUupQSoQYd4tlWBoCZZoKVJltI2H/Mk8vs0Nrb/S7saLyBaBhqGkJTY41zr0IND+6ii
Pw1G2jeg6MidjXtrjTrkdblFLSVToKP7TgalWps7ZIe4bgCtZAn9im3OsglQiZBCA5mbYImc0xl7
eA3RwtQNpCJ4gRZpeVEqirkymvY2bJ1xYVh0FcNxKOW9JyHIIvFkpiuLpX0jZFBYHhPLJXkH6RXN
djVSvaJTY2TNHYXR0OZXn7OnuL7yExEiSrgIDum53nNIYPeiE9JVHuXG3BWYbiAlYcZ9Rsguk8FB
MDYRfvXJM+lPaXXErMrQMXOymgZilxbIiOMgK0rNaqvrJGCfgvk5OTF/57lGoJFL9PzLfh2JukCz
cj1UsoGhs6ASsJFnweVhBYnFPIz6LX4QWYHegYTDyTXdkdbke5jtab/zjmOGsYDH0In5rI+siyop
HX3Yn4VP3tmdsjBwC80zKiOjialH/3fnwwaFLQNbQDogKrLqcgM7NO6+xX1XD/IiOj+b49ctTNLC
vbmPIo9h8pJyloqcpNQgM5u5oIgqg7yfmMAjgXGQPXT7BfXyy38E7Jmr/qzrm/QkPBvR3XPt3TnJ
ImywXZfM4Bd7mH9zt2MzaDzWo2s1miag2xnsle7khQ5kOKzPp9DQ5JY4Ngm1nsty8/A5BaUhxFUp
d2ZQOC4Fo5ECwQ3pSnf1egXSrSvMrFfoU4YpiLl3JX4EXs9MhXCQ3ZMDOcf90LedG0IHiC27UqYQ
hSHH7Bpo7egvYME6ofiNt7vIEL2X3E0+XYA+uNZUZsV+UF649LLqn0A1oNuMzqpYiHIgGJp+CirQ
Lx2Sdvlx0TLj/7/VtbfxS5nlAK15ocedcP6sDYgumYuJpVO6/3/lF4LWpeMKWVQLe1VPnbS75sko
zGLzIepV6aazjDqg/RvFGqcYxv83SU5IdQM0IpAHpoUpJpeEQ1nHReBi4g1h7zCwqpchobpAIFBU
EAUQVhxsBUM6wtYnYTbI9ZLNa4owCagRd6Z48oEhY21yRjdabf8TBI9CBFW9zSlIb/cjszlskJ7b
z2RzFglJ+aRpvZzfO35393pd0D9VU8afSSKilXw/mmjV4o+N9u+REMzxw2xTSfMMBB0lPiANwuzN
a6E8jQ0ydNgIh0ULqUs0gmvKMVVkADoIxX2pzbF7pGmS/o1UQEiqrSi0a2rXHP7omQMW55JoyTFO
T+sqNnNUyEwKyJcWKwVBR8GWlhnuf7o9fwIhKW+AL3u2J09AE3gzBOsm1pCJtphwx6kQh27As4IU
qZ0uY4+YcM91pDlTSPdkxQAytvfGHelQTga5jtVmLlqA9jCkKLEDmVCSG2RZO+q8CB8DR2TppLG3
X0JPQcTow2t4E2nOVOe942L37ySUJV0/t7FpLDt+EeSKIX4yfC43HDJ+IC42Zy31tGzW9J4eu1tO
ESHuPPuhJt0UDIeNSVxyxz4CgdLHvVige95WWgqN3BGlwhqI2rWdb+Op3YYJpBE0BsfNRUqPHL/v
piqJVxsTzNq1TEvm8famERwzGUagKm/+VJhsTOzLpLzeirDtqkPVwwtwNbQERVCKKaxjapShQeqM
HN3/hR3UQOxwsa81HATPRQIHAGkohGae2jiCW5vH9f1OpitrpBI/9iRN9MYNoF9cOq21/XjuhUKA
hTNNzvA0SQDBzoicjGqGaD3bu5VH/AZX6SiWAblRd3WN+5Fyec4tBVGoDiyNf7iPJtytukrnjDBB
zZJO5o+9ozroMG56uDWqzOslSpfbOVuTRLtuG66pltqtmEN8iL+qHj8RVlgbujMkGojdGP+7+mvR
C+lwk9nJsK5Q5DWLhNYUqW9+4GM+0sfrJ4QMhMUD1BekxhbwJqYXdtjLN3AdK1fHB5PsRhsjPWqv
uqCMK/mb1ffR9jrVY/re9aIR3ejGjXUS3DuKwOuoz/zYKo0+UpEoV3anm3hOFDJvyQRbSAZegugw
8Fb0jgRXvH1ob17w4/XmsK2BUoO15s9BNso0AfsIZI1GObb4lZeHmCxVaTqYMnUsLT0Ay7pFrYix
PPgbe6sih75IGjgbOJApEHScsahgMEG1wKso5Vbpaldq8WCPOttSYGbFKq3HW2NORr/PoXPXKdKn
iDBFh5t7JyyY8vy1o13EA6tLhjq86NLFTPhfQ06kF/17lrF0I9ZbJEcNgQjVivryj1e5AUekDzY+
9ISsmNGhfGtgBnS9MjFE2zIyh9FU1qyluAc6opcwwAQH5onfth0kUQfg34Plq8wpVORs8rTlbQWU
cxv11QtOJ2Y2jKvwALgUso+vyI6TYyw2aDxdDn7wWS47ebvfmAt38sLs0RhrisgloanAgif7DA+4
DJVh0VzxWBKP9T3nSipvMCiXzOOsu4nZ+psE8bkMe8WOqryjW+6os3d2tENjssVk5A9Pv2ce84ab
n+G9BYBx49uNizS9s61KOZYAPx1zsoyhVTQiKj1DpcMVLcZdmht2fONjma/Fk4SBEf6OqegHLWYl
tHaOtDj+QhmvC9+hUf2ZbSSJDTtaOJ+I4s8e/NY6q3vuCJzhsZ2yGERzHMq45B8px7cQVr14huQa
STOfTFCEj3BhsIGc5+enRvo17m2fZLEYdeWtlqloV0BKAKwW+1Rp7C5k95+WWBaqFCKXStKBhd62
9mJmLcr6SxvyAXnE2XLJNR3ovPc31jA6NIrGhR6/S4EYTmERS5nN+WdPhsPrt8i2bfuQnjzxUx7d
IRAxGIiFJL8F4q9bISqgbR4vqOSlAK2gxaL/ncYDye43ok9/Epyu9Ur+OI7UVsptXKm00hkNdILI
vpBtXKUFR/PJ7ZvKZht+roEeyDFhtjrmqdPqPqWQ4M7owf3L3F18zpU5/lPf9jXt3vwH9IApEu5c
xE0XdiMgoON+Rgm1aTe3WA3ho3gREFzOm0Oau9LbEbbxLIRwTgnZTmKmYUHSwG2WUJKl/INXNcS5
15J8LvCQtv1kg3MQBI6W3U3V6mrTBPcMHWvOBbJ1Jpk3RVcJpekGHKNCy9DfqrOM4ke5FBonTdJz
jujrpIC+1tb8nxej3ZnWcctJoFMGs+Ugr1Ah0EpzmITngORd6eFvk5Z8jvIvMSHfEejpoKYMU8xA
HQgQUNLOGgnNHhokji+120L0nvau2hwSg3S48OaXz9dCg2sDQN+j4wbIo0U6bd+CpYFMZIWkTvPv
+YTV0Bpe7V0LkOXGf4KoU13ej+QYuo36MlpN72bCcp71KZbB3dVPgfB1zcUf4Dd1FeP8ajG/IKfQ
Ag4tbsFNOmWyGtG+ELwSPRmLLeH7KLBDTdBN7IZt+C+tYva9E1b+P/VIRYPugXwkBV1M8acq5Q+D
pgwQMPEs7nIlgJ4EzuDAPbUvrURtrzk3eJpgqJNe9ckPr6jksVvgCgxGHRrh3LaaNfPyyVGSpgST
gTnjKfHVkbiuOxOhRsXa2hClvRJgn1LI+llcDP97htJqn9PW71pVVrLVMnEW4f5aIHsq1+B0M3Aj
mUYsXT+oGi0UjjMjkRnYpi8V9SCFq2/Fo1rNtmbavJCSpAXoyf3biQLPHbIqgiqY0P618SQkomje
1NhC2NU98msZh3SsZzrHZIoFYEd5RDTQkC5fPpl1IH/XG9CS6qUlJtEPHwtXQg08GIa6k3Sx39MO
c7LSb3/jpWlaHj6vymqH4RZMBO9qvGCigE+LGJ8cRu3Oe5fSOQHY8qOFkOPcCU7tDIDLlBwPdETu
BScn/Ndm/B3BOoMoFDV+dMaKMtxSEQ7RslZy/zDZACfdQyhmaw5+Y0exEwgtccylyePw0zAlpHLN
BY43MIM8cO2QISZ7zVrE4Vg0A/7GFMB4qclSRzZTwkKE6egIXddIhJIDXdREKeJsUI8IG6UtJpCe
oK2yzKaorUADMyEic+It6jCitp9u9RwVXc3gQj4C53lcKEa5z2tO9mz4gHrKClUeKhVGin+QEPFW
dblhZxqXzuqdBmCLc61RjSu8Io4okgWoOQiSRFbz906g5Ul4LaCc1BOt1LfWuU7ZpGslZs1p+uLl
MyTxVKjAx/sJ2pGw8YKUtYNkHtL9G+5I8pF3FDto5KJn0y3izsAQ+byfMB7Xi/A0VJCxfJk8CYXL
0ZeKj8Ni4sHPjfpGtql2+T5kdrRPtzyD3UK9hMB2e7A9BfMLMnsUC7QSbwzMnf3rwZxmtWPyyWP2
aZeYFrrSw1tbRWjHp4yeAHDPB3g1hb5w/CDaQ8JFPKzhjFHv7hiy5Lag1n/ysA72MxRYz2KrXna1
pQ3Hghn/nnxPMEaqgXOc42OT0j5Oy0m0M4NsqIKxTo4MJCHkqiDtVWu75DTAvKqrUL3QPJB1jM14
nnTPm6IXjgI7K8nPJnxpiKra1/lBZF5N5JSq/IEfxTGo1xIUF8j6OsdJAvsKTjqKn52UTEe3Uw/F
Uku8Urn3shoKkV2hmiR7mu12shYV3BjGouX6kwwT+guJWoWD2L2G1UqtORrllvfnCqviphHGPgct
FqDLW75tFQa/aAFuH2xAY1sV0tCnANv14gD0XWWJWRsWLKGHRYQEeMEJNKdvNtmu3xWuixS9zlom
pp52atuKzD+AfiqQUyCFqMUUm8Obf3uMMst/bDRAGpMiWS329RsL8pyMIsqlPBw5OqXpAsDbqY/7
UIKHS73hmSmN3W555QPAAALYxzzkmr80E0mjEXXKc59xNR/R2POJUi4PDtnM8GNU7cAMt3kQR1tM
r8yjyjGSdYLugtSyt0SHYhzw0QYQdPDF7466Bg2B/wWwUoesSElOK7BfpDcO5UvT4YP0s6N9BW88
hpqxci4yNM+NikaaeRUB1AvtxBjyNPKBUIRvMD4WexCSiDgcO18gB/HggNnH7PWtjM2r7ogohajc
ojXJmW7TRwXoWXH/gE/yMwl9gaEMljTwiIrt0RHup2Io+IBqKRFiuw9EusKNROJsMwrAGHd92n9J
qiDQMA2tGLTmQhsW3SfJwgD/+GhWNcHa8FYBhokhC+fTeP8VpuDOLndbeVF11PB8L0nDNt0WEIP/
ProkeaDIPtvuzhmgN1vKITVecxcLv0jP3gjE2iJ9OzDmjMuIGTBuzX1rDPeCrlhOwunkF9FWwZP7
it8s8XTBY2mEynUhMR1LCbidJOaRnM7uNs20/OIyayzdCMGamfOwksXiVbgr7Z1hXmnLb2nh6TdP
AqObg+t1mrIK1/C9Ynvt7B8jP1e/2QoAL/4AIM7aR2EeS1H+3/Quc8qEOLcEqUB0FNVKuJgnAXtX
Ayjt2W6BxNd1yIsC2XoAgWTiUvkCLNURBLgwddKfkCGih0dgjXO2TQQ907XlPFy1so1qC7FVULPd
kZLoX/ISM+TwjaTdEFZz1HmzED14kTIOpM++FcmTUvAsJiU3Ixxv8Sdkl1NjCdxIPs6RibMtkA8a
C+GMgWtI2OTKyvFgxeSoyFZVgX4mIXpfMEXB7bSX/a6WDqe4LwZLkt9X9nselPzAAzMSGxPEHllS
jNAABry8AI/9Hq7nBXQKgs67l2ymp+wbAjOfkJCcsMAvVRreIGuxCa9Dk09o1qNndCpBhwaYGWhV
hqzDpgQ/8ZcjUgKhPHrxgTDINgoDS+4LT75n0MvJgoLUbpYhHzqnV5Qk9ORxmSQKIp5HGB+FA/AY
nMw+vCavw6A0acPQW7jLuFdQT5flSHFoo17s14fQWALBbKor+nH+jAeg/US5YxI2EV5lXVO0QLGA
6csRJ9DKo8Afe13+kUSILlQNwKgL81I9L/vyPP15bZoCGp0e8Nlg7wJueX9AbNrv15r9Q9K6i99x
B5oLkIA0iorX7ZB5h/F62JLASkL9tQ6UDNlY5tEJo7OmwfGYE06y/+CkmPhEqrktscBKpbGs8wvr
ay8R4osh8od8+rP6TOER12icoSbzlZStqAsYWr98qXVvsjI46uV6OamORb7A6mCKkcVTe2DuLIkn
DdnUdtsmrMkICQkQYQAuYJgzO5l+I9PFrhJ2+ElbT8WVcoE8TwhBVQqT6mQ/7a1R956lDh+NCB6K
U52rTOMqABvf6++4GuK/6L+j9IMBDqKcBtxpgsGOfFLkdqz3T+BUwj310rZZ+QLEBy3lSiFkQv9u
yIFqS07fyolWvxoLp8t/tNFsZ8fhz71IECAuiGJUlN0W8QhjvyNhV4rXkU7YRG5tmVD6ZuWjXBt3
gWAcxaP5WVQgvj7lebV47saqIzBLZmtfIDJAxBYmypkBLE9OMheb7af7ououbKmFSbBkZ1V41Pzl
hpAVXcL6YnGED1rvUhU7/4DnHWZ7AlTOM9ax38KbQ7X8zHmYy7ndLvACnWK1iiXHNqqcPIylhySe
h7NA+NWvjm84vHphaA23HAo4YJgKJFy1a83vC9QMSebtAVyr66HyfOTx+x97jk062rcbEblaC+fi
yoTjb8buP/3f3UFGMxpcUCSEqiH6hDOqjBpMmZVeC9CzoIf8gTGwBdFa3i8IwuLy0nXKlwMAIqqG
/nV9QtjNacQHcHQBSoynqfKPJQo1PvhPUBWh/zXCUam4rpczcak1bRU5YP4AbXaSQ1j9psQPy+wO
UPv7sk/zSuf+y70JoWgPhZctyCdMbx5kcr9JGv55b1kM/pomEmziYPCEciSK/mLTjTtbz20+yxvs
T24RWjwq4kB0bvERl5hE951DB2zs2+jdGlJ5ajMiFj+SQUiNHzWyb9WKenKqEvyX8XbJS4uhaRj/
vpS0lUs9FvkmalOEi5feOHPpX73pKLrdJxoPj/TsTkc+ijIPhAppSDO9L4gCsuXuLK41KIJ35N73
r/F1Bv2SfQy8kquhOwuqeSx8McB2+9pIdi1zR0PV2wo5GgQYxg0sSIlyX1xbbD+j24sIXzlQjz2G
EwntvhQ5M/eJPMvoXRjoF7MWo5uDmws9O68wi+nFUAmij+Ksv12+1B8YqRWHK0Y42a3MU9kDEIy+
vg+Mmi31QiqMTVsgksTCcTPloyBNMXV3rpS6JJZFUZa6YxuNLKIBWCcC5nHcWixz3BMS7NTsvvJn
/bmB15ZwNaKqbg8Gn5lAwAu8maE1EkhxvqseF66P3QCldQ1Z2AVFrJrUr+D4FuE7bQ8rHAWE7RgS
tZgDhKIQ0wmSdeP4Tvn4Te7V1DZwJvD7AwMgNVDXXgukYGBKglHHCRAer/He/GwgUkWEzcNFtg1z
MNbc+1wk2jTG1zOplqaz9Iw1LXAwbgW8KAQ1hJHomXral9XKfRzZxfC3ayqby8vHD0Uv3lUO1VeZ
NhuLyqgIV0ZhQonpzn5fYINvomWm/96/0bUGRL7spRHPOQttTsuiSHvDzrpnbvgpCiyAYmj8jukZ
kxK9ltC3mpNjiYwU1CJp0h9kTaoOgddGApIw6OglJP9u4f/TGHcCHse6/tSbxKBIdd3XPy7SxbH6
PNOb67yUq4Pg3QGv25/s3ZyOnL7HxvTHmH1ufIC34GbR56tD5qtDkvV1FwLtO6+3hlOvYg9ve6GJ
GZJqmjmknS1EH5aggyfBbd27DxISVqq+Whe8BQrYSO+0XSY/fBRCCqua+w0XbCI0ZuN8CWkZAXMW
yDCz7hXd1HLsbG+ZsPIKzvichYTjzeHh9Plt5U+EqL0g4xrSA5/ubyZWLssuBoECFPy1HMHfIr8i
prEFHUoy9FatGn10igItd/g1M+Nsxmcw1/vmLFeMSFhgr9Bb+EzdhGNlYzthiKIcYOaI8embulwd
tASgcLaD6VEqh0pjQNeUIlaNpLjKKSo07CHJ0zsdrTPqt/vgQDOhyqs28+fuUp8yD/sWILR19TZb
J5JJuQuZ04Ns9prkxkIrmqaV9/oOF0/ZKzh2HZYHWswrVF9dVdwz8ghocNuips2SsGpNxoz9o7xv
U23/DfQtaJcbjA2jBR+n1NO1TWZ+3v2Bpg8Vj/YBwzoagm00Eu6jz0WxCglZmudKWy2zItdjPgAZ
MzO5le+jqADoIQk83lbYuKcvhyZo9DFF5/45jPIsEYIEDMjDkIH++GD2ig8opTxkQXWuBb+D+Cmz
WJnd6qcK+35KIgHRwi+kxacyE63WgO7+nMO3g9qxtRwsSuGAr3OQ10/PkUQNi2g+A7Z/lZsFw+M6
UlMacQx+cBq1g3y652ulAj4g/Fm1sIEucTfixBiKBkkcNiuX2tIP9Eap6YJ373Lnbr3z9q/V1FaM
HAMvKlrHFg6wE9t0aN79CC21rya+01Bn/mc2C3wnJZ60cjVSYXpDDWyGZZVj8nhieQl/jN7Nw+gD
TMNlG6ixfwDdfJkvs6Ct4fZ5enFv2qfM7tHWrX/IALvisMLKPkA3fYJnB2Gz6knVZZr9vOUdlbzd
vMdHlBF77X8S1+t04T2hG4H1IeXsPwoOFARH5DzBna31mLyGdjDTWv8Wyu8qDjTxyCW3z5o4+eBp
B1wClADUq99Ret9tx419hBtpDVa0EF13P2u1yFh6ag1Z48PemJSPxZltwJZNFRxmAImdtgsvjqZb
xK0rZ5iMONphM/s6Rcg1NgMI4Us9tcb+dQr6hOZ1kO2WZFtxqio2gR161f9w3t3ndrJvhWeO83x4
H57d/l3PDvNoZEx/DFaW+RPas+RsPVMR5Sbt9tcahV7oXwzVpPsxKtcXLjfkC4powcZd0yEtWPiY
d8zYw0NBcPov7NhJm9Pjb9+3UTT/S0sUQX+YbC/z8w2/rPpAOZaCOxzSwt54d88L+ai8WZABtaOy
9Fp1iPqIU6skcutu8PWusyufmKSRDtlog4uV4Rt7iw9O/+0WMya7hy4gLj093K4oX8BFnNtzj0mC
rmyQvnwMbpfKMfLE9dqr4xR3YP5aGKwAnG3EwCeqaqecqFabUoaZfiPx3/v28uyXC5DCsX+Tcy0n
x6FH9j6Uqj8zbOGpmjOLKILPAyf7AnZfKs0Za58x/osOYGtaUnij+G0c6ZOf08NFgn1mes+IMpKH
piCoVrPbBQef+4UFuYvY03H8a+0loG3Qb5dfi5QnLf1RkNXo6K0DNi5ILHPBthV86THSG5MgOSnE
yr9EJsP4o8F5flfjJRnavGFR2GnIQbN1Bm4IdbP736rf/PDYbQKqKzr1rX6/HeRQs3clPFM0AQQA
wAIdRBi/fM5VD1QDshP9YypPUQbdezUfZtItDz0r6hfPOuzkRMjN1iJvgCBWSP12Y4b4IoNoyh3i
X1SAUMcaiEqE8nhc9Vbp81yM2JaFUkbwUN4p8qHkDC5zEnqgWgpxQ9M92sUhiWkVcOM/06B9Ucbv
4kzECwoRjNmREF06ZSP4BGlpNBBqbANLjCMAw0fCxLRIkXXU1nWqHLTG4jz5n235wC+c63QJXauT
v6rEkC10UQ3STOpvgOAOPyEv1+04NsCPNjXopIz7fJfZSa7DFNNlKf6H+chJFHG2gg4z5ebd2CUE
ewK2fBebtSlTxdDjeMp51XxvGpxGfb7mgommX5xNEte1NMKflg1Ri0/uPusILUcFMo97qMEhmCqJ
0MlJC2oXlcUv8uccNA2JnkPRPJGt1+O3OYz1yf4OPJ+ofsWdCr3PruO3CtbxIKqdJB2xku4EKYbu
3a8lgcTscOdVP20k9WIbfjgQa6wHkUI9EfKztoBEQ9Vkjd7hK3UHC37qRHMJvf6s7Uf4o3Stlx4q
3q4QfBFGhO8xjujHHGI2SVr6lMfVEIZRPpKsZFFV7qd/9hHmZatgF9t1m7hl8Zbwz0X6dT7Aw8TY
3xyZXisT0iyyjxO/eQtbfBy1QDVsfBqI+FvLqPm1UKvst9Sa1dKyVCmLYggOW5PHvByoBD1OHpox
5l8RWc3FoNWPbk/Iin86bFOWsQA1ghwaMDojWgNOk2pwCkHmvJHN/zmNCQYN3bxvyDliPwLi5pdc
gf2ku3xGuGBUbxyjjvsWjPeCCptQAhOR4E0OIOoPPaCZjToASVR0hD6oClIFCZEuT0Gz/FZrG/BX
TbMJ+zcrfvcbk4vP5dG7xGGpwZfxYBJl7nZAZFTb8nK/0X5f+msNjpOv89WBOWTPg+PxOPqd5P6I
7yoVjS0skSJwNEMUd0ttAVip9uIwKGtisNESYAgR8hyo6cxsH2Zis/ZjjQLtINEBa2Frrc7Wd6TA
+nTVhVga0L3qbz1kdpMNPDhePnnSTvOX6DSTfl6t3eyHkx6M1x5RElenhmdcBUHMHdpwHoSzLdXl
XxnDDOzB6qgyfAtahgRcqlYlNVQPS0cR6yzvhM1AZle0FzkYF/svsxRWmw1jpqzJlxxgGpdOyZG2
QD8kvTWOGwtheWIVkvTzdVcmVgZSqpvmWJDHEq5s+i7fHXgCF/xOLY4udg0tcWwerWPY8M0wrW9j
InWfne/k0iZ2mh6XQz5byXrLZnQfEe3vq9wHww2m8cnod9g9gCPALnXAJDruAcOgRh7iUSK0vW1C
31ZINSAV0f1oJT7onpsooptXuFQYOT8zGkYojpdoLwsnNtIwPWN1Zw9CWbmxoBZ5HmY0H1QuKllr
K64YOsuoODMpYhrCsO/3d5ZzYa1lnInR7FzZ/lCXCf4IVxLMTEwqFszeUW2gWj3Cc3Uev0fyLEHd
VtRd+JEGDNCWUYvfPc5qzpfBSGvOUD61Dk9pOv4yxkeYpdt+7E5DNkSApNQMFQ4zOEsZu1nxln72
jsQ1R2o8U3gsimw0RicmfWSZaFA2VK/hX4UrHHXZh4eAKr4kod1vwXBxIfj9RDBK2NvbQdAIBOce
X7jCnY/XTQRfRpGHJy6l73BQka4GljrP0IaqyuZ/N2MXeUQK/KsTbNd53c6NBeL56AkQ91jzVig1
fDe7pX3HxGiRAC5EFHPMniCX9AAPKh4u7ChkJ2tMJxDIR4Mmd1c4lTMEuQpxjRydQoVXQrLcb8Z9
IlzhlM0cKOl1/ls5N9UXt+0Vd+Mj0+hIPKLVRJHPrI+yEEJPm6y13asgHf45E6WylfM3B5Cs3bTB
zDzZHDWciTgapB2UiDYlRC0AQQ+LRUgyjeT3LlStGcUoeuHWu5ESxd9pegDbkJ4fWqsyYUUXGdLM
6HscvlnyIoeojCYBMg2Z2svpjEiUFutncCb9FAv1zx20WbQ6u5TUR1rtnE4b/ZmDLQrTOZ0LXr0D
SnRUpkixKmScx0PRNdB9ljiV7m2e/X7b3sPbXlkg6Em0P6KtBMMUQjdKgiZicXwzCBx6Rku5CLHt
0gkOB6s1vvyqxQmYTsro3AtA6V1SVzVht7Y65mGnrAWZrxVmpLlJ+UXbrrnuCGJWaLN6IR0RlAro
oSBQ1DfyKenpse9x0GU8MWf4H8tqXADPjg5WXwSd4N7xz0766KSwA09XAnm2A8hrTeuRsmnZESyP
qujTgtbBSJEGglaHy916/2sjNuPk/d6Bim8BsBT1craCxTs0MH4w2OhZF3afYoXIpnOD0/jDSwnf
z2CC5sgU2jmRYvBGw1MD1S2xdS7FjKs+rW3YcEt/9No61kRfq7/aaHoETF/RvSRf4nUJQGgx35he
Y1U6LfS17kX28OhLItq6/32i943gsYxTWmBgr2+Fe8YfYKW07WAXb4CLxpYVc/I3YbML+AeyzLS3
GwADMb4ng2dDoGchldQprrz4pUAc8fA9tafWO/ozUD52AuHSeBacxRwbtHV3l19aoKUuNuEjnduC
M/A2Ot9RzEHBmHvil/pf8E2QDJBvlWhanlm0PfMmAOp3S0PL2/hM55KHMsqtIug0IneQFygNO3Mw
8wAeVsi3A+3cUx5ZvJgLmyW7dvYQ8Z1bZGijhELfeUf/U2NKUcCGNF7i7hUN5CeNudNl6v8FVgLk
kzZoksPgviZyZblY/wOsVXLVrnNSRQVx2sN8VRPoAgVEzXcBP+JUak+Qygg2ldYBjUFpLlxMjr56
ZE4VZwO+7lGQaXv42kq6aTijfpYM0Sp6C0ntPBPwZ5OIF7YWAQIlC2LQ6Dk/vJfsCSS/+p4qNBhq
eKdHjsdKz7Jbh00f4PvZuAPXs7f1CBFAuiSUM/iouwdGKrol4l8rPxk6+odA34dZiRJntoNV9+NY
ld2e9CgH4PU1FXGHt9RN0RivjL8Hr2grepVuifZeHFXQ4E3//u/xKAIF2kgzURC7ISeGJPmGQKeY
K4uWsH0SD/1XMYVe+vtjivInVKE1MHbl9AicgaWz+n+57npsPZdD3bRksM1DrD/GngJdX6h9IK1S
UOzq+/OsZBlFUJcLR/ldD6CjExHxqvYy3haJpaYfVagHdwjPHW+nm4/NSRr7KJWoDF0Mbk8GY0Hn
nDjkkFkGrKptZTsdYqlEif42vnfvZw8JdV6WvF0b+v2DsnoE4i+W05uKf8wu5nRSyeWPMna89b5M
fwW2Jjqlo78JVk0OXKXD+oOpemMtpPUZXzzlN3H9LQk4E7T0iqLKfD2ghMH97SBj/kQiNDA3Bl2a
SrtSExR3F35m0j8GtUE0d/QEJ/R9zbbr/aUoY70GYMAslJcIjgPVbW8A7Oq4u7EFEQbWyi4R5xQy
yTTLckTaKhhBb/gGhAUuDCVRt7X8W8C80gnWTGePdQhcXjSo9Xw0cPu5BOeswJJJ03tYDhka/qLh
tgfN/SV3AClQ0aa7G3yqJBrE3yj71y7L1TJMw+yyZSseYHYV4VDJRoupp7tbApWwfWCTj5zeQRW2
M1r+YNACB2pRBWfUeylobjp9JbrLINyrZwTbnUFszCFKe8lodJIhp6DRfIB2zUuo5R1nOtpmT3eS
Hr8FyYtuQenU/1i7rxK2Rc/of3KbRzTIfild4BHLiXkeNLggA22RhmMRTcE9tx+eeYuTVwpPLLiO
4bgutCwycwwgLJTIkT3E05kCfZr0TbHwHoAkxMwLxDILUPFRiNWz7bKF4Ev4ApK72xCxCAkqWFIt
J2keSDq9Czx8HG7MdjLw8NqRzxRD7aaVhDO4fv3cIGZiixu87D3/u1r1S5pL+ge4rAsHu2bSdx+b
r5U4AUS6Y2wttjpJTp0PzfY7LuHKDxMjAkX/kYhTFQ+HD00bFY2ZmcjshMUgVqzVsPqRPwnevpPD
Qe51813t5FJh+jR5fnbG0+OEWpmGbguTTsBNMRSD1+nF30T72sfz4mEgoXF0Nvbsa2Wt9e2umTjl
Gtp3QMjjr4U0Uj2xY7tyJJXAWjdIq5C9DpabFtyGges3ScEMGsy3qnyBAARfQVY/hyxKrUb+l+gK
pmgUKnAhLe+/mj0rMcR4nDtEO1lZ6y5Kbr8HAAKtyVaT21ePPAUABIBdPpTWxwoWePocqQFh47Qm
D4mEFkaJzqb0NrVKgB51wRNqhf1/zgHAcGQZw3PetCsMTt0eksbvLR4Di1ujE+rPAitI4RDrnz+5
D43tc6Ql8mK6pLqi2UH/co6hZl2KTRNhRX45oUi/Z8HJqEkIzl8kQO2kYU+vEmtZSpzlrCPzg6g+
Tl6nYv6chnfHTxsUGeWvO0ZZlPELnThqO/tepXCyr/YWi5dq4HPxaSFOk/fzirlGWF3pYVGskhCc
PfJcTu1QQYRRrEQuHukl87fQ4/dyO8dBqpD2MCoYf9UtH9rTOYc9RcKlM8tQZ+NCIXX8Bg6IWNhz
sHeXxoB04LZYk05zlF4O2TWa5xWIG8mvZyixxw/62PRaIm1LPC+iZySgNxfI6oyOooI93LSMJjxo
Dmg+oJrXvVLt+C8L9rxaQPy+h+N4ws9GPeZEKx871zrV2LuG7KGePMOKuAqjKghCZPpTrXgmKkpz
LxYTtRWRBsJh0FYXPQ2GM2ydxHeRKtFfEkMDecFR+gP8SEb5uvm7eRYu1lXcuFDdPPLBLEU40bkX
pP8P0J8PxfDztEBApURcgoM9hyDnmp6QNNAzWQ7pHUNZnMKA7alLjDJnGeRprjMujA4InL6jyzSM
FPdD/aVEnQLwdwi+LR0LmRqKAJzl1pE4/RNB+FNmjVCcKftMbx5EdpZZASGh/ZsZZoDVHVRIqAhy
KMEmiPedBO/QUoBkaZqlEOa30rBoRsU5womD0baWwfZwcG7eISCTdiFdkNkm3XAW1wYOUw5AEe3z
0xlfbfb/DoLPJJYxxwaKelzIj4A0Wt0JzbOV+RAPXCoz0BM8pZFVNraoz1goQUdl3faWqzYuMjil
RkdHqElkfaeTTa85hYqTFHm9ulkSkRTIiaPqIq3jgEqEhtpNryb41xErb6gFr0ZoAHpXg6bSGW/i
aOft0mOHq+3WXg64VejwYEbYTnSSa6yYl9HO5v6zS9/gK5OTv1hl8IOYjch4ab59mflta+SHnxnz
/ChQe1vcUnNrSFjuMAH6d7uR8jeLEL53SAyEj0EjUfZVdxA6w4+CSB4+ji45L0MlJamxm3WgLe6Z
v2EbKigUuNL3Ix0iTo5D6N7Bjp8n1zelAKPq7PHaa8GwSSrjaWhCqAa8wKS2gXqM5SpVSABPh4+r
DD25hbEztPZbiYcw6EUHlK0oXhXG1fhgWwy/rIqff/fN/DO52OAuDn5v83Jpk6S0r+1SHchL2/uH
p6uc23jArKspKhPA9TqdXVbW532Sl7Al+JMzS5zxQFjxNF3yNjuqY0zefIEnOnUeHvgkq9/Qj745
FxD63Io8nQtubKevt80lUFIARLppOkHNk/JfaE3i61SeqcYSSkoQN/biVURF+IPIv9cJHLefaTKU
aRIlB+KqvJl73w/DsUn4+znQrMoCCIf2PUPlyJarzIqZjw6CLJGNbepHeEjisWvsFdQnS2RpZlu7
l1k8ncdl8ccwIDaouo21TwghmSr8WBS0cDk82i/KHJn7XZM0hlu9KXhIu6e3tCq/+0NSNKzBJAQb
FOWFVZsIvEqB1gplD7yEJ1VfPHJC4mgR48XlD7dSxOsU0uJtAnAlX90iuremcwUT/CoTjEN5zgEC
PIhRezZzhVk2r+IPmrSAW35SQN9Zj0cGbEsKVP/f1Ba2dk7rVYUATEK9S8rYZNL2/NAoioFMxIgR
C8hys3Uvs3Gi1TX/BDiikQC9iond35pUA2O77va0v1TV3IthrKG1Lbo65myQg7fdalbjWfToBSCr
STAAbuvkz4D5SMaacjA6h2Ysewv3Nn0Nu+a7bIDaYpD5e7ZNWFWMy0pTxwYaDIWWpHuq7pm1oUpH
Wwjwwx9Vo2x3/Qv01xSoMcV0qR/1Gkg9jK3cPjFhfEDsfle1SsmS8l5eow1NTIv4tVwro2KC0kJf
HYb97UBxRFD2gIWojGK1NVLb5l1XR5HepVL16FBKFT1+MrxDYRZiVw7DiIG269X/CgLDBAs53TTp
q2PZWEbb0HSddXxjYGc8jTGfsukbkacZmbvBEZxDdefNC9uLWdM1v+JAGU4NmNvD63HZA2epfoKg
dT42qS6N4fbbNTVQySCaXftFeqLhHfAAAEg2InL6tbkbaP4EMi815Z+L/RklJEkeFpPipAZ0K3DZ
7pIUjAvmpOS/Eeme5tW3SuL+YT/zrSa9A2LfpIYxI3XJTF88ef7I5PCcoCAFDimmjY3dH9SmiO+Q
q7Fe2kZPWJijW5dGhIJh+w3Y+V0Dt0W6SsznG3vmzRygxKaWH2vAix6MHH0oFTvJfYKeTftWs+V7
FLiWo7o+DcfK49g5W7/gBqK6DcPw2d5AakeFnAdTX15XXGlBHH4iO2KHTXrU+2ZVy4mRAjZZFpdA
wSPpLRp2/k4qefsfOUFG10NCdoYtTqesLw4fk+4UzWtsXFsTPLggnTpOHrWd770JdNu3/i8ybdXR
YsosbiC6pnxILI1JhxWD2gQqP9QYnW0DwEzsFC49vGYAH+04AOjg91DKo019+H7QcL4hPT7XRzum
kSuk+F0SV7+7T2j5kyH1mVIsjbxDGuRiF3CZ5iGHefwmQR0/OeobENELjigd0mHqrXXWHWDsrOot
oYZxrojzpjjaoDXpn0tVnuhKxWGyHFDoGrr72BEoAk39wxYmZKMk263r6x/Rp/fzeimmiZ1PvDL/
2iNH6VwdKMgwmtxmiBtv8VYHjmXnFwGCVOLiTK0ANkVj1gk0PsC9+Ex0Rj11SueaDfMRPfNy1e9z
JYqji/A3teupQwzMRWiq1yG49D97T0IFtgPVUyxZ/Ty4syV4aDWUVcbIK2NpDwvanAzdTEV8HRb1
dNp/dxgLeONNmLrN2RlqvjaS7WBmW4++P6UartouwGpWBPQLNjzxppLNQHeklvgKwq5ZVtHSslGE
7S2EmMUTnLA+75Xj2CF3LM7f+ri86JX35WTU/v/zXQXGwtZbv5lVZszMYu1Kxk9weES2mWI5pIdn
g8YF4hb6e9ljZo5Ek24ZH5k18/L1k1MMd8hC2qXdvnyWV9AjFRF8hsHZI/mhe+H/HaOaFztlfpIQ
Mk929ta6nA9qRmB9Qzz1vGwTK7opb9a7aoTfYur6ZhZs4sjeYDUB6Aq0BT39nex0R25Nf3EZi80D
DyvtoQaq1s9o7Ostqq308u+jlX/gmR4ID37KSiKtiOI4yEJ/fdLCJ2WoEw7+WgSAX5c0GWqT36OG
Hxrb1owycNBeZou7FesGFNSQMXBflGEy8i2ZLBJZyTmrsoOCcTpzVkngA9qAw59WH57SUMDssCIL
jidXYHGNJwSwCMXQ5WRd+Ty2hzMw5+NocqvHS/nzzUgf4IA5/rcIk37mYXBYe5g1B1p6kYdX4hMZ
Kb978dxSD+VpDKR/ojFKA7KBvyXEyUtTzqkS75/CVkBeQQqQepCq6QVhb4rT3o7bCYdExi0H6Zzm
dHXz8u6STyYfe5zto3vLTQS1LnBhzU9vVrj7HklPdg/fkAD4mNFuKyC4aH86xzMv637Uyef5JPwN
F9uwIUun4Am+DMeHiNKjuDrvn2EFwN8tgZ4kpLla2P14Y7VAy1qDCJ6lT4Ad20aib4GFs0/COZcw
Bm9492BSkjoQQxI/g+13dbwsMgXRLr63a/IUJbU3Z1U8W8iB9X7SgGvgYON6kc/N183+dxYZQgF+
dO9/dCx8u69ZruDcGqqRkprtzRn3NFcRKksV3EKsDfcsRtV4rAfrbrjn4a6gXnlK9yqU4Cy6Kq2T
HU1+xk/YS9SahMq+9qsGUV09nSxPTETWmCYXzeoxfqnhFWU2ERV9uVYqG//0ERcwqVfaC7VbxJ+h
qpxmBkwyva54sKTGqpW7wUlF6qtCdnqP86serxlzmp9R0Gryo7l7Kyn1ejMXRZVaRhbmYklOx9EM
JRht39pNLKsoF2lVo3KDmOAuItTcghVAlr0cfiC9g9MhvtDpqj6iB7LeuUVH0JLB5Mumc4lt2wAm
rUAkvUZvsB71ozqRAcQ1X4XtLuVdEpu+RQjEVk/XAIpOAwyuUXqx/1JRGYHygy9B3W0YvwQk9Fdj
x6dq/ygvfgo4edFuCOeowf2RjEQkR7sR9N8sZBTTB4NQxYn1VyYVeN72wwGzxm5btjWfL08PKP0N
n2x2Rbl7sJyCfLdV1p+vp7PaYJiE+0Euqb7zw4wgOj7s0UfGykRDJ8BRijNUycdN5mv/ehPD5/CH
N9pbSb+31hG4uNtIrhIhNoj4usGwjwrfh8RUw4kubGGjGvdAUIzpvBepmLjCKqVNiLYxQsJ9jQue
mRY623bpaLo/FIVTE335/xDyn2VSWWAl3jWdeqFkJmoHOrNUtFXJGFmySi3ifAG8fLFDaGmY7ub9
VKKzZOGusXLsYP5HtOLUq6VzRGt+wnubdgMybhTPcceSnlcnfgbVzulPDtcdAdZ26BbHYCWSFUOE
ZyQhyc9xSl28T1w6d0TrcSrsTpxGx13UxgnwpWRiWzu+vFn/rcnzrlUW3AluNfTNgRhK3oKN+Byt
UgRMLmiZzfmycO7qQgWs9RffSBGjHpsPsHL9bifq3Jd9+kDpAvwlsFId1GPFu47nB9afv0eAzh4F
+2qK2AF830McyIkX1Cu4E6EmOKWiIntOQ5HkHjb+trhhmWkREZ+TwndA3p5+YzPNlJ9AQrPXDwj2
W0bVWEkOK7gw7MjgOnKTNj9rOZwBeT28hqtIvUKjw0tteT3PtxVDgwwvDKL9tv5PLy6uxHYkOuZl
Zei3psILEGxBuRh2dlpTCYfAYDd20/cdLNCx7ou+WKvsv1dNFwc+y6DDey2cTs2PMqUNJ7bkq26/
MIQ6fHrEeo9suAX+HVpxdJQy1z0biKK4nDKsbUkGsUz8Mjp0aXreORFCayglnSt4vvjuEn5b8F8d
jxfQAyPgKsjB4IsNQtjNi5qXwAftZTWr/uDBZq5FydZZEPkuosTrNm0knTQrY6q1Xm0nfomMSzRj
QBLvnHPeQJqPCQ63ZabXyh1u00+mmGAzwrSW+C5QqLjFzabmavsEYyvhQVI5KUYjS+Mx+dzShIt9
XP+JjTQ4TXfoXqr3U/ebr6drCPUOG5TFWtCxAGU0RsJHnTVWFPySLCVUMmteurrVRr2LY8e24705
FCvsDGOdW0rC+wtO/HiLbvl6l2VsBBt3KT1Zx7rLb/2xoTLIrT6RBlJecxoK/8dkHnVIHQ8wk7ug
PxaRB4NUgvNm+h8HlHw/hPaIZNfriQO82sHmMuO79sd1ob8502MUAH+MJ0cJa1XDol0KeJIxg9mr
13Ycsnc0jCKsSAp6SKmT6u2coROxByQc0Ec07faba338ZOryTCkJ74nW/0VBfH/nwsr/QPbUVV2Y
/O5E+TkrnLaHNAPOLSTID6ViJ9VJFkypyf5B3DTzacR39Rnab+ALrz8b2yLdkJ2C3SaMvT3+IMQo
U3I8COxngnM6gkduDZUmda/R3GRcCtslnZZ+X4EJ2isfgXkh7xRFSy2xrPYsT2oR4sg6sYcfa8JI
g7cJj0SHYcrPS3/l8Gl6H8w0PrFwMyxirCxaFlrMA190bIz6cH87JakXFGrEpOXNnPaurZL2UqfG
+RgqZ10g7ki6fcYxgONHrCB4wC24HtxeTdyrPigsTfvktP+qEWWdyqL0KlhcDIdZIDVdP4dOuU4E
fjHyaF757FTxlBleMQnXNRZGjAVOaRZmZzuShz3fud6XEsU/PZDEw8/oNgrKfx5cCMhskpaeTQJr
13Xxcwyxi00cta36rTuApAH7k1kYycs/AvJBotDNkMgbAq6vCc9/RZNi5EEOlRon56F5bT9zKJGY
MVJIvygLYVzztW9zkTEW37kzdxsNaDBd2DjQDZvXpnVHmp3EgQfeFrZHzDJP+1PE/Fc7PvgncAWN
jN5XrqRWXvcJhHOcZcAeLhQFaH5Qwu4df/irgEdmouGw4tytmVVFkZFAd4UiIBq01rVhRpl05EoL
kdg5x66xDSIkpAZoAEzjHbWO7GFq/SNqGRFgX1agu/7gFG1tM/JrlbHIzPMhJ8fni7UrSvjZxi5w
JQed5MINGCO6Sj9+ESkLHhl7c3ZkHZXBvBA4RzZxassGZV6WczIHMcmU7KysNX5Z/evbxIwlmXPZ
zlDQp4xJq6gG2lx6IFpMEhhb6dB5EQSWR/SWrlk8BwG5z2YlNZJGweiCJoTTNBPJbkjTgNUUCDvM
GHRVtsr34qu4lgtv01QG76ixB+QF1YjO/VGEPYMSj2CKDifmMxF98smee94pqapkvRAXoEj6QZF/
G7+/AVBsl6shC/V9mwJKTMnFSDVaNsiQEgeHqfeECtNxy3GqwixFguYVox2xVYZWbofA58jXfjzH
L8hunvk0mVJnm37fOKMBdDC2l/6yQ5IIUcalZX7aa5vjn3DuVBrV3X7aL1BGnQ5EyMtmOk384zFz
sOnjmWdgXkIHAYDH4Ng09X68w6x8csAWuXey4OUzFuy+voX/OLcsRvLFZXGyVP0B1lZCIIZu3C6K
eo3Q7nWAhsAtzov2TejjclxE+xyr3piErYupb5mrkfG5xSLtGxZqL+kQAJj6s0VI1BokjrLGsmfD
HrXj2jRxmziFEkW7VhgPPfb6G3FSzSt1hSgsOSKULWA+P4Hegw43uDYxCxSy+abevyVnfTb3HOTc
//RDUuJimKRlb7aWijyEnO1WzP1eVVSaSzi+caePZk8i7BB6v0npmb/VEqNDU0kMUST0IPGMAonk
pC+Sm+itD8jHIXNXauKQrX9rsI6vR7F6I8bAGC4ruO1MFVy4vt5LZcUH6L8qs4591czPFzcl8dgX
tBxy2aNXmLMysPn4Q/PZ18YBPgViPDPJi6pjtK5GdCZWEMWriEebQxzlR/Yydwe04OSgRNrtAmjT
eTot+Wto4mBgrSdbf1OyCzvcz7JSiGST5QHvARVxDA/YTN7hRjuG0Yac/7lE3AHRUjqofIoCp/tX
O5jF/Q+zEMudSYKNWZVr9lm9WtPQ7ewmRoZGSAwqIHXsQDHWCn3FLy9YGRiqiwnco+E6Kytst62f
uGkCnD8v1+k9gMZuvMJ6zsDPsZk+b0TMujlUnErcqYLPgp+FQplliCmn4aquq+cPKbQVAxG0RmAn
IljcdorhMfjVLay1GDgCGz+QFloEvEdIMkySy+NOt+J5BzOND4D/W7KHxYIEFOI0JpX53sOYLYpw
tFwA+FikgK4mTfq05yQo7sUKTwC0KiNBRDE+qzBxia+KrB9+j9L2yh5mogHlqfpWmWSNIIjeV9fK
VR12P8IoNAHSOI5balNBSLWy6MJ6LG9YagBTBiu4QkiEbaB0lUk0wktrE60PuvZxAkHDr6CKTcnZ
dTkRsGa4HaX3SJkGNDl2nBTnBHzQUfdSVtS/v/08j1wx8ZqqOTfYGqRp1n9XpI8XQhElT8loXR5/
Kfc3t10hItA4zALFztb5p/69CBpLiuiD7dmM6iUu823EWKkWqRELM3yU4cYnzIGUzQa5TMBwtR25
b54/Qgi/mhRq79vNUGQT2JXC0wmbLJevOwhBYNj1ylTlbOhldfCOGP5BWpuk8GvqDFfSiwStGq2P
Tt5AvU5eXVAYjNiAZuvCN2thpJdD5WJd8H/nU46w1yY6GWWj4QsFTscAeDx3rByXJxwFXSI0iUM7
edjhlzDvbAlKgZCbnEaGJFCtbj+nZ/Wwlv+37wpkwjICtZa94mSCnZZWu7TIU5mTiX4K9PoCf2nV
HSaCjYZSuErow3Rb2hgSRK9WClz0m9EFPy8A4SzOmoy+G7GzmAYNUtg0bwC7Bk4nG0KGm/HPFg80
kkf/kGI4nUfi8FjHU4LxrprvUou/KlTKtxGrGOWxhEYO0YyN2xs2ZmeOjPvhPxhbc4WozUET77W9
aQIKjF/IiWo2HD7YTdBOt9AobHPCjbZ7gr90jBqja+yQPleTgeBnqYavvbU+eXEn0vRRbaAnqrr/
lqLQoqvLDthjhm8e+fgCYwtGe4h5GFTw1vbpgjTNZdEY3KDNp/T0Q6/1U36kSl3jlfNy3ipyr+/D
PftEIbSPgTJziPu+OGzePKJwUjXFY1ZHiJjXPekiyqXNpGHHFhDvlxd8B3yjVqrxeSr3tHc9u7MT
ana6OBLYrXeWZwQQmL3wOVX8+svou8z8BWei/+l7VDCZD6OSSJrDOL/NtA+lXiRvxG2qeklqkery
yOY5izN8TEAN0kkivzFyqACb9a2bUbtnngpmzes7IloeClKURwKsYROyA1EF/CJlYLBRJy9xjOVo
EqKRZOrxPgwiCNIzQYqrjSU7wyaRBCpmsUruA2Pibl54kenYd+1t13pHmmGQAvXtHwos/5pNKf2H
VpqTcr9h/9PwWUVY7h1gkpRWXYunEBWeCto4m7o2YVK0da1kcA3iFeeJIEZftqVuw3vlDbT4gXFW
M14e2aluR6IdTXlKy5T/WkC2nRVEiQDYS9N/04viL1ewr0VtlG8SkacTqyKQ0iLRWpkBKG7kf7uJ
TMF43NG1HVwG+h6MSXNhlXgTGzcl03PLb45UqRXC1ijVuHHWsfQC8NxBMg1Rte4PnSLeVns4opWA
sAdTESUglC4U/8TVQXGWNEY/fro6WyNrYF69JvNSrbVSXIRhTFWvmr2WieQ3WhjLeBK6Rw3XO8/j
LBYLDYE6qU7Xhdz/7K/8MwElazgO7Vu9a6U9GeBYBMpXsYSuJLXTGTQ9TCzToDnftZ/0XimpA4+s
oa5HMt7bdxKDMFuxjKgZSRKHbK/qlnZakhmYrdKj+WRmUn1fUXdrZBsan76QR0e2bKEZ3jXfyCbS
l5e1ArqGhIx13Ub3274WOYF75DZl0potaJscgdaqodklBZK4tcnnNvu50dI4Z+Ya/XNjF7Wllqy2
ge2U6PBd9QDMsiloBZQbRy+pK3kio/Tl1/B81dl1CWEDfAYcMcgPEGvhgok++QZ79qBrkK/J34HI
QMEdIdcfxtn3JLV9mZ4wjLKaNPO6Zeo97Qq9zu/znt9dyvFI+N7wrg9jXZn48Td7aLFWZfXXQarb
dk2k8TL4+rfp8GfnC/Xf9IfXRINzwzHWm3SB025GplfHndiLSKXH3Ga1XRhvF/JQ4Yre4kqVOXth
RbzOfJ7B5p4BerY/XC9D7YII7fWq/nk5N2ezohVjdxFkTloXmAVXpQZFGAbhGx6Xf9ia4e8SZqz1
djmrktJXMb34ZdD+VnLFhhfGkWjEKVcT03/ecOf2QA+G8ieKE4cHy1uyEaLQ7QwnoHsaYSvMGIws
CJgLwPh0cREXhIQujzDh74WU7lY0sG6SwdJ4FGtajPASQskIpLTv/6tnJXsH9wLz0rTBAbotRcnL
7D2b2TKLCMreGLoBTaeGAzLXO9tX/uh5Joqr5RKFKNMOzoB2nnV97Xa47GnKhphmBrjxnBrGNgZ3
NBGYT4ULo5wm3sE2DJt64dpGBeOlNk6YdDhl3SOyRqMvxbxjtASe/7dAUylnFVvmB+MTtKHNVQm+
KeXctafDqK/npYEHXDoIPU3cSnQsZIaQk7XsCOo9iMyPgoV2t4ximmtj6NcNWpjYYE4C2oVORTDu
nYOECMObF052f2bhOG6wHSIXiaeToMocdRZDoXPepjR1iFKqX76Qx0eu/RQGyBW4LAJeP+S8zlZr
bLBkrs8yDkxUV8aSSDR3IuZPaUJp+rYHdwj9gYjYsX60Gmj1F6sZShlbJkwuicmDqOpMmO3SxVgw
CeYBWUfruK3Eac1d6zPx501cYmvX9ScI+tXvLUL48VDUUlpjJX1OIKWMudx0F4ONhuhSRB2qC35b
irrfK/jAN0x4FwzrLpcxDx5XmNjVDBao8PMVmW+bT0kilttCEZGUCmBpGmR26yS8z6jIZJuMhYYs
NgxuoWP41GoaGiN5Wph4Y5yPd6VE6mloe5DKl940DhqzrSAOKhKm6vR3lxnU0ucVF5hm/ek1oxqe
5ar4hvVjgC43IYPq3Fmcv711eVXNBhyyzWXuaXGRuRGzLaYMYEnaJ1BrawgSrzZFPcPoHcbqIQBm
VcErn2T0gSXbgq4U5E8y/N//4hbIHeR6pFc3RWF5bS9TiYF4hnTNEWytwggL9n9h5RcAp6Uib0di
LbFTPhPKUsfETHklD+NHHIFDNPjsPQTtaO7CSZhfyoGZC1sRCfHkbU1uL1z0yX3/CSLxoMR2Qdtp
78vF1LkTSuhqXvdIGWAUJzTDNWc/0QQOlEbIawSuZZ3BGoTJO0Ri0cjOtjCBwz00phE+wOP8Tjm4
VTayK8r8PsxtdFsSP+vCYNMTVGpkFgx8KdSX7HNRC6o5f0iKJpFDrvZiVFr0140a6TyXciCIYxEd
6pE1m5kRMv62CCdlw1T7Vok5TIv1kL+X/bZq/nFrwby3ePgZTPAs9ytDQ0ia+yfJiejokmhjkwc9
IR2nmVbd93FILw7KQrgTlG7LKi4BQFpWoMcrnGLU1J3e4ylgtpg2kwGhLBVcnLSX8xUidcYcntnF
Di4jYHChM4JxkrvbE5GYj/d5bgzzEDotuUPL7pv0SHDF/7Mkt6AbnR3IDgUsPgjTiWWisQtmi8X2
ccZOL4zI5lJlK4QgpSY8PS208ka063yQtfSR/zBuf6TwboPwYbb7B3shCr19oS5fTTzwzWuuBhtJ
TwO5b5jHjRnTmEGNg5rJZbx657RBELp9tsP9D78ORaj9MCd/QWatzXavDRCALciZKnBOkZwBP5i2
gRN3v71oqvANx7Ltg3p2ajtDPV6qpMUStS+Mzu7tvCY0wDMDDicILW++II8XA8HPaj7B2cwGQ8RX
2HPHp4G5YV0r58s4fP//dkzhWTrbaHmeoLGziPpCpueOEWcYqQadSrJqjyHhZEDgWiDe3RRv2d42
AuDp39Gsoa0k0SH7M3h0zK8VekNgrKidlrnnqnFckmS7G3Qv/5bG3222megglTeArxx9C+gAzJ3z
gr8hOGe8LuS96DbpIn4UfSVnED8ubEFieu56Z14uqe2EL1fQG/X8qAP9CD6PPHJzL2M+sa6o+5Cj
K2U65/jBbp7lyPMohCeP60QxyQNxFkksT3fcaS+D2kZwe5VB1QosH0wmGpqOlNp4u6hMZB/9IjtL
PTerfh8oQnvM2lm1cRZLebHvc0haD0U5kWzVkfyCKistspc2z1zw8Vn1DRgTZBKN3DJQay92n+KP
YkM7HyJHSbqKorNMgGdxvGpzI/L73T2fyr++mN5SkQ+toJ2vC7fGE+A1qMdk+282nhTyIzA+DsLh
DL3pxPQjFpVByNjL6TdYvf7LOCyU+z78bKd3k+hYdT62Txe3oZRjGwOe56iaVkI0OoYSw12hvepL
j9ojzAoTE4uBxGpqeB+EqxBFfqnJp/Xv33ntawYejzevRGnqofV5GW7kO9ZFVyG5xmYFMEE89oiq
SY/SLDSd4Cd6y0H17IIccMkVUaAUyomXj5c7UyfnHod51vSk5uDFKtAucXImy4D3LyNrjGpRF0qt
Fu2asX7418SBuMI36SVyhNrUfLnz4tQlW1Gm/h7sfozZsHoK1BSUcgFgsyjt1RDnbbIxWgzCMmvp
ckUagsgV90wYKB6Xq1QhqkyQrR8/CehYI8ndN1tdWtqj3qHz3O6ubIi+96bmJ/Q/Vqbs0LLVrzkQ
WDgK4R00BqF2lKF1klD0Mh5q1CPfAo94/0klGzI/mTOSs9odhDTC+ykLLGFRQ2fZCHy60nbQ8QGr
0ZL72ONAFcOj0Tw+YlRfEbVkDkyef3dQA1bI8bIWv70EpIDhi4J+Zsq6EkEgJA1kF0Wc2QXzvS1u
oXuro+o72QtsydGHh0+UUF+RD63gPDDGw+racPonoi/KJGjyCnxhQV4XYZdI8oPNsUvgiOlqfmFx
8WJZcp0fKSv8sCyMsTsIoxglz4LsN2zsZ923foSI3Mg8f1K90t58hoXJtuf5DUY+NsgESnU/zyAS
/azSkdjOeWEIINP4vtQfee3bvo8k4Fxe3e5PM7jhBWio6S6bBXa4cXnez/N3S/5hIB4fcV5kfc/m
WaR5+JXmSvnAnA/gcVy1dN0+AqdJxLfIfT8+3oyj0ITLD4Tkc90Ce9UZrSkuvlrB5kR6WBIJDmng
8FREagZ4AMfFyMREQ3Js6mWgC9IzaCE6x3sgGkyx4ZOvb228gnnDToMAcUL/5dGvoL+XawREfca1
WP2Z5hjL3V4VMWtixWXLxMl6B1b07Ha67LigkIbs10utcsEerv+HBoJbfBAfDxTWcw81b9QI28bG
lmtS2M1Uy/jRiv1TF0u943yHsIhyZy0RVkawnlVh67fmeiYvc2dIa2ZZySggqrW8ntm1hIAqGso/
wFuO/rhJ8ASW7p4p36Cy6znfcx7z7Jch5JqXfr84NfDspr2eIjg/qnsq6ov8iJuk8B1WGoTEnxp/
Jdz6yvaPc1AwA4RBS66ewInNqy77rpXRhw8dBsEs0PmBXeZBYBeEy7T02Wb6FexqE5l7nNYWkHdB
vlxYTSdEzm+6iFAdJVM9Mx+X3eJgplFkDu5op6iM+pHzlo2WNKMojz46LfMgxD0UNWIoT+wGGw/i
o0EpfMXZjC7vsCdAurYRCzo96gyNAEtaA0Nz6H4jAzEcrDcSh5BBCWwiZIb1eHKCG9+3hYqhYHuq
FlHEgbpC0Omf4S/suyK8sbDc8xR6snS1zr2fQBrxco71mNZLrUPwFi/wJEhInE1p7xig1FTl8Esh
nTquROLpmpuQ+cbr6kcfPldBveM3vVy2HP+fzoknsdVRyv+nYPGyYfVUlJv6Eef1N6Igfc0Uoe7D
IgreQG1E1ayEHwH+7zaDix1Wb7sb5t4WVo+g+D8nB0bN1CsfLs7l5e9huxGP1gLJlRjaJnIHEt1j
CWcSiYKE8gHLdNx+5DGPRHwv8y6S0SSb0Ad6MXr5NnUacTuEmNEch7ki+aYhwDZ3L2IO1+ditnn9
axUWBBylh4HxwAEmtCAUz/XO4/Nl7wxyt97DTs8ocObj5qCnaMEaGr4fK4qxX70527rYyu4ZHtkV
zkV+FwILwq2hYxSQ6JAcaGjPkxvlYaUGB7lhSVES6po9f1HxeaX9sOOR4e96TNivZ3K0a5DEUISS
X1TV0JQ5MjsEahB5a3HD9ODEgjh7fMdrVfh0G3/I6Zi2mmTOXJ76mKNcIjozfKkVmW8p33w9Jldd
ZvRbfyv4CWvaS2ytsSVBNae4H4To/n6oIsGBQDAjE06/IVvmTOAkQhjgNqYgMrvDZvTpoXkYP+Rw
kb7E2u1gK0hv0p/UTAjR5sfTRP6MnANpSRjHtikXzXY+t+F5WKJ0tcvFsSpmgZVvwRkJEwtQHswR
PVKQ1TCfSHaeamkGpPySY+oS2allvqL9deWctwkFlrOP6Ry9DEC7MvUo8mVT/zfKRFdfeM2spApS
QNQ+ZPhwqNSfqUWaxCH4xb46w/PM3tMpdC8iGMLSL97TYhqXpmzLiuUbQQt4ndtRGMQGx5SjsXwj
6uOdTsQvcKuMEVwG9af7hVCi0oOpdqRdPPZNMl+YvcQ43PUUG0p4ItFZekogt+9gm8lJi1Ya3dsV
L90or94yYEgF4rtCP78qRG8FyGl81d67S56SYphgt3aP4A20aCUtarA7MWF4/imtiffj9Ta+K/aB
T+oqyoQCxn+l30c+HNRQ4/9QdcUbCMEkPCWhrZl3TE8zoFzP7LBE8TG7PNQPa9plTGoP4U8rsSU+
Z1cVshA2KXdCH6M3lPApAIKUxUxz5LwagY9Dan2j5FtXd9ywqA4VhuHCWnVvGBbko5Br06z+NnUb
r4zqCwyo0TBSaMlIC5th/jstMAKKOniNNgIsYCge+AFWHM+JwYsJoMAev06A/mjFuC1wlY0ZCPjd
CQxgz6Zj2uwwlNu9DJjRUWhZcHpGzAGAREPMfjR0EIrVGrebLIfbL8+c78JVFFKzL9nP66FCwym5
qWwt/mlhpBkdK3lvKQnKmCs8gRe9qvn/2JqJcWrUtvURQE+iYTa2ykO/JGVRtStX3aZt69JOx4eP
+Qi7uPEPKF6ZkUPfPDPakJocgcmCApq4iXLm7v83oSdRLTINaNRtbjnbFnSjtL1Bzfp/ig5UBp5k
6uylQSUUPD+afNubvBMEwltxsdH/x/igTYArz8/wckORX74qk5zeBnDriW1B1QLcrQGelzSyTd1R
LMw5OyB8jKbcB+W1+ufcQKHbhDtXMkgbTpUaC6Ff6nof9xNShhpyrkTan84iOByRIZddw66iUePM
BUEKKcFgTue3iV9+3EhWriQ2HLCdYZmfoujQoWYPlQP/HVhZ+LfxPqOQyYZrCk1VDg19mNhISfsA
YXs4wg3UMfOjQvVmoWeD+5FGa3fpMEr9gYpu7DbDHsCHdY6Y2IdhZ5XA31jwbzk0Z96Ha+tXs9WO
6XiGYB4Om3ExgKjftRwB8SGugTTDVotGTsvcxPAuuQVq9eeKlSXdjH3l1ODMWnXaFJZSAUHbGs1A
BTkw9y1zHAsmi08oBp2rBuCqyF1RimVcBCnyOeD7VD7V8/UJSeJp6QMyvuWJm78UCLRrolSo4qqx
LwKmKzeAnZpfeUSjJsqn3SZRIuytMPcwz7IgAbhqd8kCK7z0dsVc6g9oTBgFX7Uz5TkxsmbUNk2P
4/BYaNSvCo6khGaSDwrbYfGdi0wuT+5AGp9g/lYMXu9hFNk+OmNoOPD1XeaPNuUXRMY/MWjCi4Sd
viM9kOpqWD4z1LP6tEpGXf7yYY6LVazHhColXRwXCXah3PA8nIz4zpNi6DJjzEAcyzfmNO7ydQSk
msHbwqnT69lkVdbdLO5YuVznc3kpAoIU2yAnY5FMS4Xt6MdZJhQxYkJhnVCTTD1sDEwpU58jPB1G
LnjuCh0226HuUkbeApguqm5i8DTnARr7qEhLlPqYhIdcuV/BJ/xD+6Ese/RnEU9j1n0SRjnAk2x4
g2lpTPoQpxiSHz3HfOp0wZjC78tGbPlVzFhSM2NKugdS/VFSw3jv+UO3OLobKot7u4rPpTKB0cKk
YfOyj448K9roXAKtYuKlAFobL5S6Hp57MRAVA1vc4bBHcUaldMYukF7uDtHTk6VqQOeM0zsxcLC/
GEQzFmPZI2tsTFkCYQeHsVLaNDjUY/aH5MgnCVOIXGIdDPWFelYuV8Tmv1c/WDjXv6sFTCec+l19
rcJVQoQGDkW0aGj3iWlgDyrpfEyWttAaNzU28ixSvMjaiLdVEopgI9nJD4T2JGPMr1+wkGlAV+s9
i5WHV6hTnKzLXaOaamjqZUmwDvgqbIuKExZZl0FQl3vSKfpdfgCBlZgdeHExD4sdt04b1qjCEBjF
PfKhy/qsIEPbuB9AvB519qAwa51gseB7D+omEfjBMoNjIctENBQ60j9yIuLxdgNyIiWmXkXp6QPl
i9XyZONKxtOV4o9psrmDdHjWykvGZ0J5YEdKjChw59beMi3biS44CVQlBLDLKaALhvryiTuH1piK
ag/xH6lfEt3AoqwYLREZUkTcWfipu30IUp1Wx3SXz+s2K7mPzI17JOv5DM/niXRP70gojn81XvCB
0wrQOm3Ra1R0KzZqYVxx1sTzB1tJXwpkqPFYJlOLa7n6bxVyet1vM7g6SdfYK06JYfK66zcNDgt1
141RxenP3tQYaZMXMBLsUyh360do7mtfBxHWHI2FYS+dLSzEHSt2nCR3tRj0Zv31sWykrBiNdN17
D0ce3LfZXEK/dR+gaIusMVdaGY2VfTacgIB/Aqr1d6S6Z7JvpiLOcQwX0Pih02Z1dU89rCmdvMZD
k4PtAhq9meZw5UrcUhY4DKpbEGX+E9l4hP8s8+ADPEe4E7aoS/MK/Cqg/+LUwRJdZyNS4YxOiPJ4
85YMVppeGZLPcmTxuziQ+SUk3HnY/5KCGnLglIx309WT7qPU9c3Mo3ruNSG9g63hMWAoOPk2CAa5
DTAx5iq2klzpwqNe4dkc1UIo5fCG26K8gccEH3VNK58dw1Se4wlg3+QCkOaoZCeIUGnCc3FALSEF
xFVwSbzCHxjayPDRROl4efs00E1ejPzj0XlEGWi7X+rH9/mlEm1jz9uslVMSjbLofDnoFeKIywPX
6P84RFoooMr15v8/CHGrTOV9/HdjbyJwLLCAZCEqIR1H9Jfl3lNIzCkxbKm68y+97fSv1mPD4pwn
oYJTp9Io1Pwrh4Lvg0fxt/ibDfuS3J7zDcjzpNUbO4y/kb6sLlZSPwfRjr6zg9XX1yxhagC4Zhdp
ezecKye/3ezCL72/wZBKgrUEw+XL3JlXq5YZ88LeUBmEfEcREV6AxpZJyqibHewCn8alAsS0pSTx
Oh3RfnXt3p5ppOcvjhpcB/111tAJZxaTk4+FDzXyEGU8RMY/p8Vxasqr0DjdKBzaB4BuIw1s/Aqm
vawMW+HXNbWszVgbeo2yzc70EOexBtIqZEcKOXmxmKItyWqa/5amDKY9pKxMhZK/HiR0a2/C7+Bs
LRXXYveIpTxwq/ewc8N7Y8MXTyuvlzkacGG4ET+QVKD8+QqCs8h1UH41xVeohhojT7MJ8n+YgwI3
Ay693Q17+iuD3sFXB2wP8tS4gpVNOhErk3sw+lU7ZttLAlDvyndSd+YjJPBrvuzGGxLC51CdRbl7
hL5xV1Sq1vS0xN1Jia6LNV75D0Pxijh3GM5s0fwd4yZriUibGWUeFYckX5MhZjSQbM9ivRcxnkuR
CxxTu5wE4Xqc90+GcJqlo1HVSTzFU1ONLzOMVwin8QtLj3Y5vQ2vGBMJeXGiS0vETuSJoBxwYqws
rO0Pg/N4MujQ/2duDJXHQgaVMyJFxDpZiUrY7AvuhkELbZxuM02RttAS+ij6Qpw9Rh1rLN+F4Tix
1NLGgqzJw23ENhpoDVmFE5da1YZPXgmZvi1mTPtTGIYFIHTKUemZJl9fH8dG4HzdUXH/zn1B34Bu
Mfvs5GYkt/y7UXHOdLj0R3wk7RpKsUXTnsXvJCZiRiAy44zKDIzcuywkFmrSV5P0qLKIFD0F2KUI
DAOBvZcw+HD8FZYS/3Tw/wKu4C3u3gobBQaxSOHAeWDyksPBgpNqCTHMglg40L6qTT4Ri3lhLr2v
Acra874EFivuckvHRUmrDiPNlwEPfXlJ9us2O8qN5DciPvK6cc0sAUr2N7Ui7k8yrt1lyisu+QRE
0fNZXk8hXgSnX7P9fjpCGV1rqFjsl4xXjXX3r3EfmamHJ8I4Gg9nkQY5d3r/qJ4v0dTvqRdq9V7T
Q6reXeXj4QrTTA3khVYJMgNi26OgTpSIBlQcoN9hvztMIMVYM0QUXpC0yhHGdA6UKdloCJ7HOpWe
rpEQOqVYb5FnXDpSsEhFLumErpgzKN0nHyVE9TxUeuSHD3htxM39PJuuvoiVw3dPEpIIPPjrBcKr
RGiMPVgKf2J/L3LNAyxD6g/nrCgUE97wu+lLZMgMKp8r9OHhz9I/l3HVTp8YJjdT01g6neMUeJ6P
01QiU1XCf1AkwLNzClFWeA9y0y7Ekll/fsO272eVbsz/bnnWfCEr1qU2HCqWL1Oge+0xQh1lrr9c
lL4fH53S8RYe15MVBt/vePI1INmshPo4UdEy5OTRyQyrLqK99NTJMwp97ZYHau+WGwIb0Cwk81rA
W/9wznV92OXQ6b3kTXMMVB4XViebdRTNN1+3W1PGcEowk2IDyqGTpFj63TC0OO/XpSkvbbIbjLMR
0S7iNmzJzv8AE11hgA/HywMgTS4PpGRxNlU0RM7JNqMy5L6Vd6B4IV6Rdhc8kLaErgBnSPF4Vmcd
pzF1xvZyw3q7cJJ6xDDurTxiHIPAPYOyl0BFe9YrhnUL1/7/z+yCuoXPdGCfb6h5niUPI1UPNree
1EF//DxREowAr6JWlh75+QJB1jBaiWrN5ITZT0BQLxF7mgCPX6Ax7yKfx5q87clHE0Hypu1o7G2+
nGCJpMA4B77xigREzIKlck/fRfzAHckA0gjxYNsbeuTgdSa5BMbtIRvP8RFCx7SiKlNRgMdKy8RK
ehx3q7JPh5+zvker0TF6K9XFnbv1O5Qi+0BUP0lgCIZUQWOtX6pEynIgwZ+DA2Yd7+zTjQ1tgUzh
R7xiHKq2fq/Q4jca1guC+1u8AHGsJL07Cy7hjUfdlzPb405mf3D220ticUuxR9mVRa5I5Anllusd
jBFuueG91fA0mbEeHM2pmdw/KKWWV/qn/LsgS/QAI9BLvoPRtepc6vjbAmkCX08K8xJupATYIB1C
hF4hu7Wt0NxHbX40LRDJIJEsZBGPPfC/KN373PNg13y2kRkEpsvMCAgT134I4wNvay4hEdQof/m1
ONrk3aUFIatAQE8saDApI/eLMXsTm2szO0QUE08xhOzIxnxI0gwJ482963GF0EzP7JwvlT/T1Gg1
E1lpdUrD8NKCK46nO4Iqup9PNq1G3mxOeItnz+++h1euqLKHNlLJ0Vgeadr9XSX+xS9796D/rfZ0
8p9KCOutut7iNluQhnZd7jcZ9dCKz+1ukKcNuHtqqaEj/sjGa2yOSvzV/c6bU1PPCTLf1O0tUzal
6bY0Rx/NtJzhzopk2u2gZDcFGNkj1aCg0EZFUdIOZlTL2t3gJr4I1XYfmaPBel9QR0T/Zkqxjgv7
2+WW6LWdyhGoizxSy5lgGyjYsZXj6Jp97si8gzJyit334kWggQ/iMmbbDsc1P6YoXVWaAE4A6bzx
rDdRmo0w2ej0s17eQ/AO6TcOLeG03zS5wFKRK4JDZ+4Jc7rc032B/sBKAjxHglQU/VnnalIIPaev
i0QSwdAUq+9CKrCmFEcUN2h4G7CZkkwgCm4PsocQvfMg9l0FJ1vJe6dt8H8PJ2onsComyDrR24GA
VIbvRhKly/FBiSCBsBvbaaYZ6rSicrJ+lpAEo/lPNj2DB1pGCBLQZGQki96STueaEdh484Eqidkm
h828GQmYMVR3jpmVFkMn+Labshj+pfIgdmuypyl3BCaLEb++SsIQ3LObUR3RIdxPbMBkg9h2CEOH
LLMvCHAD7EqYmPVR8THpuW/ETQFC4/emodir/kPl/AgfMZpL/ohjKnvgCpYdeXRlucOlhyFVQqEd
satohbvLX7JlxndlmIkFPiUOo1ZsX08ccI67jhcRay5w8/qyjy2eSdsD5qvawZwN3mEZZMtmw9hs
8bD+q8YZ3xckf+KUTt2iK67iEwsG5dCNOD71irJK5S98nCO8QHKlypeewgBbQZkvH7ptJQwyHnsW
BJpNs52ukVilRjaCyCJg2h9ymScM4zFl37f2nt8xYqOtMzSdZgwmcL2SzlV4Rb3GfFW3jiX+IyDW
UcnlFdqp/q7Px37zNQI/+9og/Ymb7X8Uank1THURdfrAU0x5JSDeUoajVBphpkjLM9/8APa3zIxe
KALvOugkEwsz/R2JbYk4K/r4EP3uHoGtOhvtBILQJl0umYnEFxJKzTGtGGabZCqWNanjm634apez
0GWESp+q+NukMFAZSzBHS9+SkHpdkSNnw+SCIQ98uPXc9TVk7Bo2BYLX/m82F7azZY3OtssZpvg5
Xqut8il6qoNWlxQKHBiKg85pfYI1zQORNyG1gxbYaWEYRzcZygn9cEzQAn3mPmUbMlwc3ZdSyjOK
a8JNkDXkanxM8zW9VXYf7D7cdUnhcmUr3+3SdbevKvZvMZeUQfh6dzP90qgHnb3UBIEwvgYq9hyU
LSze1oQMPV+rP3cgmv/FgxCBNPtdcR5tHkdNeasuWz0HUty3u/sz+Pgy86pYltmenYGJ2peQDloj
ACPdXxR29O5GD4QQDrcXg6NZ7ox4H0fe6q+duro0ImpbjY2XhZz470ExG/I01xmlM7AW4Co900Pp
XRI0NbWKf6moWnvopm5xyHBaInptUFohfncKW1csAHoV2BhSIBG5tDx7UItqwyx15GJXPnhizMXz
KrFzzQvKNoD+R+8OWlhUOAtJZvtSlYRO7g7E4EUNoz9LZBnbFVJ9KevXdk5REp0c/9kNdKtUkIhJ
jWQJwQHv6ux3VOJXRQUIJNq/1+8H7OkiLIJU6Evv8fHvv1PQW0AyJofuwSPlb0Psv1+t6hSQ13RR
frAaydtor7PSC5aavtuEAMm3YAarlcxR33l/i9cjcyZo1c+UTxP9Deo8chHSbjndL29cj17QzfXh
YLLaqnmyAP/EVRbr0Uy/4498/jOqbc8cioyr4O0OnhSjQYKbx9ogb0WhI0vavoGnlqqpzgwdul78
CripSz2G/1B3QOBHvwOZ1vZGhnlRKp2jRFH68eshc3SJyC+WfaAT2FaZdJ835uuJrzlybZHbYFJR
N3Iy9xbWkOCJ54OGi73rldqLpvWFPE2SfHJvigE2ox02L7LQQK9Tj54MTO4qq83IM5uCAZSgZ168
a451maEDu/4wCNjAh5FFbG2G4UoKk3NWCJx8I5RfrY+e/DTi3+gqOM8GsXI/p3biE6KseXuN3YLK
eghw2n82HrjJwXRg9AKaWvTnDuri4Lyn8Ou2HHJpjr8zPPH0imqclbek5vI9lr34Htg4WddzSPlJ
Jrm4sarzI21fMspDzpopHDW8apAT3VgtqjwBV2Gce2BjSIkBiTf4mCmwH/2Es+8mXm8k16IJMI5h
SAJOBahxIb+JvflMf/DSYcBnOUvvjpo4e2pZRzDgLpPkTKSNRx2OQ/0GEzSpfi/hf3X7IJ3oOjZD
QZQSbtBqi6Uycfa4SHs42uMCoCVgBC4fvqQnAI56sYWtUw5tzCcbb2Dy6LltXtrDwVGhn9d74KLG
Auo00oNPbOeJ1wY05O3kO1XFlbUJQUOaBCcmbAK9QNNyG0hZw1GcW4/aItuS/U9qaeUJkNrw3VJS
sYR7RoXFEWDorN4oyxB5VNN7OLrMQanT2qdIncKdvdNxdcHyKko5k8KgrgMCIJ9Cziow/pJJYOd6
0liac19BP+/1n+Ri+70XJguS/LTrYbh1tH+SaTPJMj3j8zc4P9BcGqnJXOQZbaZ6O3Tc8VL8hPp9
sdOuyr+HgOlLUNjIx3K5O/5KiMSThos4DEVUND+aoZ7tvNGk61K78EINRgMALCO2niUkfnIAzY+h
DAXCEGI3KcF2AS9t7bLMbkDeSFDhifi9O7hFZlsFYEeoChnbtnrHYuJf9OW62n8fHCgSe1kjgUyZ
WXe1ewFcOVRtDvbQo0sU+pharXsjwiWkR9ys7hHu2xqLxZXpSePpP+BK0rTBvOAiagJcbiNUSOC0
s2IbGMDS6Sulr3H/FiTsWvyX4DX3tom0TOAnBWoNKvqj0LON7dsJ8XV1SXpbxvejZ7mBC7VZezow
B1MMtS9NMrQStjN/oD34v26BrjRKu6mycdIu9+/A9krFa/0helpGVcqfDIKV70w7NNO2k+3ZQjUw
d5EKfsG/VBNGHc3T3YQWG0qBOUWal+gEhMvQGK2l3570RQIKUe9fuPSuADN0e50zIQDQsdx6ymZZ
d+6rmYxl3IqlLpqLzMJR4RTb21iX96m724YkEPxc/EZbiUq/3Ekw+VLQHOUdH9b8TiiGux2v+dGk
xQ5KNBIanmdeTjRJQE1YttXFhHxK3z4Bod3ZDcKqXlc848sZK3vQYAzl0k0y4PJq5ZVIDZ4H5F3r
FVdb5whGqHn2kOVbcKnAPKMX6fzYypq1mitb8W4ow0tavWK/Tu4WUOpXG2kjUSaiZkvhYeWq+GNi
/YVHoXQeAHhCTHATkztUfxYJbi4dtfjUL+G+krlbojr1miXxW3t8KhNHz6r2PiVwQwCuzkG+ssF8
3gFGFSCnhh1qjCbmHaWkeqwWqjWk3drt3wC3Ut4tWWWbIBOEm2G9bOizGePONRNE8Z27tUFboWaQ
IihEoniejPY4cv7/Mu3NTE0u1IFDP8ITqyxH6UsGDXRvA6zjIOa8f4lA5OiJwMov0MFTHZRNwahv
4XP3MFcu1RNYsScK5nORCm3VfsnwMDWq6tSRNTp9+eHXAdM3tyXrH1Oj1PzGJOO3MNUABdVipPsw
GS5pZDsOuWen5rxornolpqZWwmjiGBcS864CRTEIm5N9Kjl0nDmtAcvwP+Ohk1wn8CPpf4HUjd8D
aPpHA8H0F+PXxUwQJlLRVfjfAETVyiUh9s32AqN3LIcYWYy1QWmFlcZgMgNtr7/YZJELMRoSXckx
fUwPIxI5VRuzHhQ5gCHvTH7pAIGPZGvQ1jwdDdLZn3HPvLUeecaWObeENPNO197US8f6Hv9ZSxdd
V4wO7vcQxp0Pp24CLgG9QtPZhppOju8mkr6VniR/onlYH8vqWIqsjNw81QLIlKPN4CZQcHez9eDo
tgFHx7fIAGHLxkU3V+jUou5J/Qts48gs5y4a7ZqH5+wvnnGQ/VI1VqJqZNbQMUlI2YW5p5eeTWgu
T4Hu7RWfZ+aZHf3goW8YU10cesH9wqYBx1b3Txc0PrzV4CaetAWzqKzrdQdljPvc6Ldv9IFy5nqJ
tuYFrA6HNzSQaafMo8i72atNL55R6M7rHwgP9L9sH0GtC8pyBNZ1SP2S1NYGZf2Fe6rPgm2SuYRk
9IXeSWYOxCbUrQVFLe4cnCnJRlO4nHZ7RXx8HQaTo1HolGoRmF1k4eb0S1v7K0giZbG8pgva8ljY
fzbO8lV39FFTV1xEIjTxLwBToWi/OaKTLBewyB/dzYiqzwrRE+X1G0AmtRl/KrlbcXMYgBoUJ9XQ
aUuN3J8Odhi01pJdG3/2zU+vex3zdkiZIWg9oKKk9wdW+XMezoWK5Zzsuw3weSacWAit5It3fosE
KH355xOsvFtgVhyZ/DMRwCg1H5CD/3zzkHkiohQ1mvj/iQli2nwHZE/vCNJoiKj9B6MwQgYuBi3J
E/toA7jCI9ZyYUoiEstgXtXl6Q5Vm8ubFVAwz59q3nRwFaWd7yGuFoLq8zRHgOLnOQ18G4l2M0n7
vaonOo8jpodrfzgkDutA7yKXn16NXORcS3brtrGZOI0kqUYwT+1y5StGNpIdsnsUKMBxdAO9EnrC
VGe8tV2UAgpjdqvVMRlgd8fXCxpgETKZreIy23vAKV281qei//3YgPVFCROXQ+sTpbIZkG1um4VN
TJAKt0BfaNVUYFHQbHJkH8/66pyU6jvahzfQBGXIBGKEh+8qkZhTzjIfY47HRHVwbH2SZPfR9Myy
3fYlFABY6lX0lKe6L7aTiH00gKvA5/lr4wWcsVFifjKiu3jDFNcL/lzdNF2t58m5RCkSESAF7kLz
Rj5Gjp4nNOrKcwjiH9CmTMZOgQOvPPikZl8zt46jEalZZWFK40gkto2QPw8jrSs7F+RP0+nNvRiM
GwByoKhloEV8VpMFcuHgsqIy8mioz4Nj/w/b3JCgToqr1OhZOgxGRY3HHxXgQpMcYH6zwDjX+ujw
hcQ02EgMoI5/sRe6yAR0NsPjq+CSolOKjWwcowCpewCGU5oyEzF9UGAGWIuXO+SoRzLik2xq1xuP
YvIyI0DYoQqGufG3hxEnuuiKqpoRMM6LMk17tHbDoL9pVaF/OiTL//rxTgJm91yiiL6s6JFOM/z+
WgJYiDwhFtQTc4ijdvMMH960ZoBHBOdxuJ7WiSjMpTcVMqh0aDkMT44n9UqNo6PygeFmZpMr0qMc
6dT4KmD0PUYbg5d7BglfFCfx05xX6g+4dALUS76jHmyi2mRwi5VDYHSlu7k2nJ+u1SGLPhtGmDEM
+juMwt5cCXxpb00HxFORl3Exl4u9Ecox6rn9d0Nx/bW3kP7HjaJMHkIYG9dxoeMtt6sZnuBCh6LX
UMspJNiiXTOpFXJfa3+PAV1wvt6G/F4xgWijDsszZxFbqiub8/IVmzoG4b6XdHLc4rVcmjsiQXY/
aEXlHzDFFF9CHFqEW5xECUsFO7bJ1LB9XGPBnAaa6TmM0TrgtI7R8JkB6yOMiYjx0NlvuzL9c4jZ
Frv76QYUhrn8wFSal8CGPxaw8HBGjAbN5Wv/7rCO+qQqsZsKzqOHYAaWFpIIOx6vm7efNM/x+y/o
HeFeSWXHW6js9cPzwXdUjz7Dx20+3Hia7g9Pwz3VJbtaU5uVIWvisaNDKe9D44JjSoYr4If8WN47
cq/6G0jurKcBNVdPwayzjuiH0NiXvUDzqc8HqDavYSRzSiiSFyuGhY5gr/8WNTXySVbzPYx9enLu
VOhLJRtYbuSmiwq/+xKmMfiWpKiwR/INRrERjep9DmGIaTAQyzU5jMGzbzAtUSihKdTlqxA8LYjH
fxbooymPC8DSVLCxTHz6ZPwYqlAKkpIJm3GLQOr0umyuQvDiuzInNSbV0JfZ1WJNV4MmtVxOXd/M
hGV5MuxjVktfbsyFtLS1J1axwBecjiGY2MXAyAI1NPn5Cwz20A8yyRGk65VltHeef6B2r8JB0fNW
RJGM3mWcUjGAxvAFtuMSjwNEd7gB/afETxYf4X6owhNJNxrUtqRb3hqhpQKkf7cRTw+JZNujemb0
fELweevHRGPFuPdOeex8wAM+tU/9Lx/32cT6qynAhR4yVohqERqsPWk4Y5IMNWwrrXLFV9gaehvq
RNXxmBd7aBpQ4R8QfxbtMmir4zb3gooG+JUjmAJmN/9tYn1AltPfL89SPp4k/UdNy0JfYF/ipI0P
XvE33yujt+Ocdr8HVOYNSrpsvg/o6Yw6BMhwPtdjBmfuBzFxbLcAWhLzWv0H6KxFdJjAc09JJAHL
H2ASorRZJcjFI1AXXZZhexLnsF/RxNnZIrayTatcwFLYKEszCF1Q0Jnawwr5jTMeNy59ANxU6c3o
4f32UTYvAfR6EHYfmnTh2ONUU657jT/S1mhEXKaBW53WX4MMKKja1bj7rS/BKizDzOwEXQ1DRZsz
CJazjwlBqfignv19nwznT954EkQeGNcJQix3hfud+vZeNZW9a2J+dXi+4/UoTD4Xw6oMYrQiERvL
z69upvdvvzn//cvovJrH3ZerLzzZJCLaudJCOQdeIeNrt9zw3NScPjKpVvZOUT0eZUF642NxLVoE
AoDEH79wlHQvDt3ywwhgESK1qkyOL9/JkugOeOSqUaoFKNfOUsbaE9uV5ROZjl7o5cOZe9kLosMB
pdoV5WufUEAVAfH0cBDNBrxXBc1lNDegC6El8Kj36qHJJRT1OzHH2MOg2vpxz3aSWYObKF7m6Ema
/+vzCdkEfhRHqDn7DsqjWsMd60n50Z+tQyDT0taJRim9+nLi7YUb1CmOwNmDlnDoh9qSsY3BQfOb
X7+49H+WL9xcDTa51J1mM2KOWbxZiEaWhrDCUTbO81Y/zcXyT6xcOeYRlYzsCg+vbF0QhQF9dSGw
f5VsX2jbCBMe0ron6cvSszW2Qh7grxijHyrisgAUB7aU6Q1/GDsOiULvI0V4M2ezwURSPqM0TD4c
kP9cl3ASubkaN+t3XlIRwCRDSGg7xo+aYTe5ovTakSZFuH3PMF6mz+xoN2Hto8MO8GnJxRbl+Jzm
OrIU2zCFoRAkSpK9LSvVzf4ZfH9vAcjfTKQ+FukF7jJJyGTk0HhdSdImJg77QSSBbjPIqFgVvkVe
SouECHD4ozz9eB0VCKQ1j0ZgleE8oCG8QT5WMLoZkxIYjh0bQ31Eg2f4moqk0//rjrcmbsR9QUoY
kU0eTGtSZ/vA109VLu6iR2lRIZCZHxBrnFhXZWP+mi5qu9mBC3P25Q55PeFmAY/Xs8Bu4z6vyDZc
YjDGfaAM68loHuHeXsd0sPdKSP/13FyqFDjPYZYFx5rN4M27e2ff4A55mxOgcEehrij1Src8OrG8
3ag0NdsnrXFmkmz6jVbCOE3Vd+yca1VqHU+XyUnoGarbrur1On0zC3ZRIKt99Nte5e3xGCslNU1j
rD7w8bPUK/f7Miuuj12zkr3mESRVh87eDXcAuw0jcd10jW0YPmktT+XHApY3I1Grh/xWny2Kr/wN
H5nLEO8fe7/70t2ViGheNIAbGmNHoLeZF6vkxeXuVxS+3/tBY68FgNVobVv8820veZVe4nTj2gbL
gvtGr0jKNL/bFw4cNXoxZVslNoP9kZ9w7HZ1vhrqWyGsxwQbaxlZcaFtD/KXerjhaBZgivJy27S5
6bOuCp/C2SqKwA9NpOTeiMqOhdP3VD6z/Z8/5QFwXjq9dDioxhWSmVFtTI2SXB/HyvYRnbqSl757
q5j5vwMYPJf5g8LQ007QkIMz4p4tILAj3Dk8em9EBJ47lj3ann5KybU1C60Zk+oOFoMLKadWjJTc
h7OjdNFPyxgr/FPR8zXCiDwTFFGT/dDrkYR1IiL0EUJfJZZnCo+ZsnYxrobqPEc2e3BkFugXieip
rO+QMwSBtlMW73g/wRMOrSO88o+y2VxOwJtrHT40PRb6TXUaodeJuKbDr7V5g+QFMC0LcU88d3qZ
G2oIOBHm0DqcsoJXh7aIds+FJmPx3corqmQMdw3Le9CUKXHgItueQMv1zBP2cDpuzzSEe5VLhNdx
Q1oqplrf7wQRkNH1TU70wW5m+IadeEf2npAXB6oLuvBU28fPQkBFCpHb96VD7aAGNm6vazCWlU0k
yx1Dp03UUCdosdnkXPqtvew3LnYB1O8fVigpy800r58dWLJdojcSQJ0LgsrZ8HrCrlQSJvYj7TtT
AVFBldsL433CsZQwBnFzNWU5iEhrZvaDfPeFJM7yTjBPav9XsPvW+u3ZUXvGPrYylKnht/0iS0dz
qCM18inuHHewRaLZ56z/o/xF8X4DHOdeEMjt1FosUqDUl6aIKSFJsnrS3LiNqd9GFcLaaDF8K7+a
YFiREfiqQwfAFNmLeElcrMWj90XSQRke85wSI0wb+ruEXVhftKwumMlIumifBPgQ6lAr3SSFdh6x
//EYwPJwoJO7NzQPbKfFYTDuk2c1n0nu6dRNS9tFhK69mv5kofHP/bqKePPNmLwVNZ4lVwnqodPH
Lv5esyxkPj/9VK/OGrwv5RDbmay/xmU4gnjkH8+1CW5Fr69KaJqffnko1+2x0BAbqDBgl2e7YLWk
5DJx406gyny44cbCwMiKfxBrti1szcxV5CvTjqU2qJCeGb3TqbgfSloFEgzs5c2tQNlmJlBI9KQT
qQ76+2cCohtjwlLwbjgOhWx674kBivGOe0Ac1PpMlGU8I1W2oVJ3fk4WLbulf/Vyhiaj+2zHr8oL
Yc70RCn36zsN49eqQjSxWWilo4S3/YqwtREB0AYVqIwMmI3B/Spare3t2RdBqO+CA7LUCnn9neC9
X1hTejO1nR9QzsAU6urVUk/XCCBmJtnrlUk3e9GtZMQNR2pJchz1otMFbeXuElYN0ZxPIMuNty16
7ePE/JhHuxqYF63xM3tpwvY3bjOzVPTi6zt5XHlqDJfHqTy+HnDOK2twkhsBJ1sDq80w/dcZ3oup
Zr7F2Xc6S3IBeMuyLm5FN9R1Pphbbjzr/zeyjaib8ojp6ilxgaYpcgqEc7/1qW1mzkVPM25K6Sb6
vg83gzwNLLI1ctKpIgWgV71YXJwYjCcgSVv/n6MMJBNnB3r9ZfpEQHrD8gS0LB2yiR0FpSxjwcxl
LrrAII3MdVH8oURrNSaKF1kLQfPU55LOQhObs/gi1431uMxK2n0g9wLr+JbhoVw0mOfI5dGs3yTR
iUy56Q5vbGmVKrH+rM8IxkL1QNrVpnPp+8xR6Vadtgp5UGcRIIh04tLMCupLn5v9YQygyXO7657y
SclbutIHvfD+vXckC/Z1yWjqAMhFWQljwa3hvLs95zCa0cvr4baoz3qbXlC2altZHIqNwgLO/Jtu
GqP6A2xc8RfcTho7haBbzHSpCKPr7fGUXTN28wAlsqYFdzb3ffvwpgQKzZodGQUNA1jeYuE+Mytc
4mypy2d7Wl13JD2WCrIMEDbeYH+jSjSobBVWmqdogG0ypTvnzEVWXvX7wiPC8y/dURJpWfENSmmL
yZbaWQ4vX0WHYnxrc/gC1/5FIb+Q2K0HdVUKNwoHzgphpu1SErxp67pe3sQGn9gienLaEQK10TvH
7T04CWvNGVFXd1ZEWX+DkB+dt5+3YU+wkzA7gSQo33sxv06+v3Dw5ObHnHArpR80vVV0uE1pVuzW
jPOyWB01UZ9Y9Zg1hQnCdSfJwm2muW5eJTS1qR732lmy8dWdYWN8/JgoukvrpE1Aa78LB9MgXtan
7QLTzDDZx6CQUztJpqUYO6o1fCCkRhTYNrp4pSC2YPzl+0Lp5hCwMKtXm2cMjwHl58V2eHATMBgn
YyabP/4zIirv6cOUrEz5gC2c194oUBWUa6fW08EFpXrr+ACDrbqEQgPxw4Wk+Ln8YTDo1R5Fsw3y
4HqKyUGDOay8Jx9ZFJrprV+wUS3FyrHRRVwH3XlfP4kccw/59GvzSxpwpACDXn2MYTddecVlSelv
5hHO+ZlYSzLs7Y8H5b6GDGVkjytsDcWgnt7AXm1itK/zSuEBh0MstIRpvHTKC4Be725NZWVOunKh
oZAD6ntocuBQdjSuyZO6wRTaRMIjZfzjZ72fdVMMgZK1V6rx8pp/2ZBY1lzElb35o6jyVfCRjyj5
hK+tRilmV1LY7k1TS37jFtmomxC42jNev4yaVB68LTrvgvLqfunPRDVhKhT92rhV3RoYQIn9k1cV
5DQUPPXNDq+qLfV3CDEQgK2V2Fdm31rYnh7P5G2eS38wY8xSbKq2tAuNnIm+ko0ARjeT8+nzcADj
0hPr/26/+NHEs/CWNUtJpRwvsU9suHDezwpF8O8bXFIF+lKi9TxsGRmtUGdHLjSZkAgkSZOQ5TpG
9a0PiEMRD7uq89qOsZlgLR5IYafmdP6L/dWz6vkTnbg1nlbPivq4pZl3hHbcOWxsIgUc7jmzRiq9
qT/9u2kv8+VUeGCI5ZRuyPMkv2fB7o6DUGkO2FiS9q+IrW21L8WDwXdSfjoZnQcuOZbsaFgilgfk
3JjefchiNgJ+BiMOi2Ig2GghkoGLHt/w61KLZN+dh8rjEwdt7eH5adUzDmmeTUiusiw/PkUDWSZu
ezhO/SK1p+4NvUG1FOvvtoKEHZicC95rwDy3IMa09Z4hcPj6xDzWDwibL4fYnOcyuG7ruXa27pWK
lVsekUWpOm9dez4Zlljlo9Gnm+YEJ5OxzT/1fKcpVarKUbmTscoNHjXfPvwaqawSBCV66zqV8uih
VJcxEMIRy24B4wEebgp6FxkiQJkUcGKpm69qe5gMPYp0Keyz+jzpv8VSHnG55zfEArQ4j09U8h8n
RaKwhCVU29ZNqVv1cWnGX2Hx7wjH0AHkv6WuEEFPLjkXDp5cChvK3kc44r/ktt1p8VTnBdoiG9Vu
nQZ2f/TW67aisVB7MsMlkBX5GLOnwr/E3xWu5RqhguYC/0PXaZFt+eOeMB7m24QILvfFw8ZgdjGQ
3LgXyVJxCS2lWO75cBWxLTWV8Hq2l99FATJLCWx55621QicJMTPoHHmA4NqpOQccVLRnluTuxGWE
Y+YqrK3BawSwvebjBq0I3TWFyiVjr0C2zD0X0lLr+NfmFxvinlhKTuN95TWVNKq2Gp8ptVSvuEwg
pAi9QwGT4HjYunDaQ7+Gh3aVVxL7eKeWoCu5/ToAIyr/5NAmRlwMtIpLyrHr7f3YXzYmb9ppzQgU
z3Qrl0zj7axvN64gkvG2oADbTO6O1ppSgKB3jY2xpGvRsF4HZ7TpjAF8MSNWIbWSbNl2joHh1AR7
IsM79PT2lhjRwupWqxXKV/O92Irwhtfz4SGgb9HfBuPNi7c+NnolN5iGMbRomP6aXoUS3RN97gmY
VEKGb2dFxAuIpyAA4MQV1o1ofdYW3CzzIcgmyViHrep+0/egKYoFuLB/uDj1NkRsWUu5ReZjv6Sx
pQWsGhDEbqO8VsCHDoLmWpWemj1HpMv0hQljAjH1oGyT6XoFNDIRki8Ft5B9GEB1SjO/FQsKAWI0
1LUQ/7zHjs3FfKnI4AIYc173kIx+T3x4pBOFaXjJDu0cMD+5qAdD4uC6zJef2HpjkGhK4VPDjTiv
mlYZAca/6JzMxUReRrkYk/7LIA/+Ol8rPAkUOAEedk/uCqO01VA/T4uNOskl/xh6kqv68RF7vVuu
ptTI90dkIyWYsSSd9aRazKC1o6wH+DarkhCd4KReG3wTxQVjGe1nz3hpBAol91ZYhYDqUfdYO1JP
cv4aEqFrxNNtX1CvVAnR9gQX1SoERFfYRa245kvm81MksXMScAnJaU/8UqMPz9v8cMnLsvarEyqP
Yzjsy4A6FHtKomMvsjfycpH2XVl6I6yfvSCi/KP1opItRH2GUNNWFitZFNxGMJ8FIRck5dfXZxMo
AUZEOuiEsvR4izKNY60phPb6XRdAHBPqL8yvhKUsD4aiZwKpEq141ZRYBh1HKnRiyCVWVdw6ywL5
UMf7hYJQnsej0jJUno65tUFmnVLYtwBfn6gJuEKz3GQdZcNz4IjSYg7UYy6Jlkmye7qLSkgGlolN
Duq/oMstmnxeNKlWqUUdz5s9EiKxC6Fpnc9s9TqJPeMb0WffimiGK5aIMVTTQ3xvoieywdKeeocI
azkKyPT4jwAR9009ZvGo8FJGeDXN4blHZDumd1yTNBRulMWhrxDxnRiBr17OZWStuQq0ZV09RTAZ
E6Clhl110+az4CxbyvlYIqyLxqhIN6JOwH+BnsHOWDcOpEMcVXA9CDeFkPfYjhbjBiE3wkErlgTj
7Zcr37JRT1TiTVYKvPrI9gVOcnj9ff+IoOH9jmi/agdGNlO1k0jpETy1MQIuyTRqnlQEra4WbUld
tUY/g4EMBzZOH2LdFioTSs0W8hnqsTCqWJelaLbCtu4tDnI1FZ0fuhKNtg9DP/gF4o3A57In5fPB
s25cuNblUu54WV9XuvABN5PcKYJxjEFvbE+M0YiHXVZR62uLgtVBnd52o6iGB9E+3FdxzsWewmLC
ypnVTu4JOq2beaPZESPFHFIQxmMQEZuGXxr8JiW8qigbuGQF6b7MMV9/8isW/ZtCcNIgSGx5jrQC
snDLlSz95u8SRLG54eMq+BedJjvKb93KRICV5DR7tmFrgkWlprB+XOgvxtzBMdO0a4LKSQDLziiK
Fmt21nvAuh2ZGGKw8JjjPkCSPYpvY3nscFZKC1SlVd4ggOqHKayZh3CnvXu7kN+awT80TrKtGAll
KtNFJn0bC3cLuaVd6VJXjf3fh83zNhd+IGW4n+eSXxrMGsXQKRfbwuwr1sRHP+wxW0p5xK4TC9/U
97VXlewy63oZVDLYRxr7t3uO451JVgC8TTYdEn6Y04D8Hms+0FPIbOVgDa+V0NdknUt0RJyZA/zI
ZM3uvtzGtih6hXTDtwFyKLuIRK+wt2TBAuuUgOVnh1eEKMDPDpvja1v/+krKgbYDd9aRBC7u6Rzd
U1l6pJEM2iQ1Jasxgkx/vegB6wpxSTwXvD1FN4cW94PfAzrb/N4RqKZb/5wDL3atQERXTxTF6xqU
uplfmvpAPalm6HXQYBw2eNf4KakmGbfFpFbVMxvI3tLEmDlba31sv3cTQcntJ+Nh/J/bXOOz8HKC
WbsSW5BEzwm8oAN+OVKEeD324jWV2LRSpr7Jk8oSpzEUXFU02fc1rYT//5P7HbSQBWWdqNjhMxSF
r3yNjTez7LH8CMn02zicX/KQBNGd3q834+8eRkVzgMgIc6JgfQOMbyN9W6mXK7P3tybB+EdIeLHk
4hkYTQgcZHTce4ijEeYrsUHa9sbZ0RWWEASh5dM8o+XEMfGMZU1sXlRBTGcL0BLop59uoOj1E+uZ
tpwHIxvVaz8AzB7csazBztufuG/f/xjYo+lPemb+Sqf8d5ambmzSa+KcPEmqXCOb68d7Du6kAj+T
+uXm3gk1s5F4egIo1EnDgqAzsJuYMKY2taWc3+vAIa2A9djDlRXm4QgyGWAR0AGjQAe4a8Q1kp6e
hUu8TNAeBlooHieXOpMnKg0P5zNEHj1FlrbMpN6HTSn5fEA1tOYo6R43KciclAUhHKic7IaCgnTx
at+4j3aIq8KfVPpl0je8UAVx0SiWQPrFfy8kpcniptod5x+CHmCJMtN75k1KXGJY1YHEegHCY0Me
4iIGKUBA+QHli95u5bhrHblgQzToiFx9xGnioDQmseEOWnMsyy/lhsvt4YyYaRHZ6jcEfmwnQanj
BBGvhPJ/4+M25sf2NniPue5cwdJbeeDn+RghQDpJrefYX7ROAWJpeFeeckdODLsQfesD7iDjXfDq
X5MHAOBMyNfDTGZqMtV8m6h4CpPvQu3KyENME+/t3FTKoulkPbovLeRcOq443hiMJqMks6VcDy6V
6abs5vjD96JtNK4nD5lSWPMkeBW4v42zuLi7RN6ghdsHuaipQAaPbPfNmu8Qu5mwzEw9tgdOiZJa
rRTMReFfmFr35CPd7PzPep8FqyJAQlOyJzDJI1QuTohp+ftak7xWlOeRDl297SXKnAwc1WHzYDDu
p2D1//0OKrv7eAi3aOPy8TdIF/v5Yi95GrfRuvXJSJpbXtyfBRr6KbgtMtCUAuHld1eqy6Dp7Dal
B0WLBugiHzxu89gZOQjOIMGPNMuuCROfzTW5JXIZRLYF2GSnb0xwfM7wyUCwbJvPT51Mir09PLJV
YccehQ/sXhDskT5erEwm4hKCpttIggFxMnjDqxR3xwbPGgnlExFDCN9FOzzAdjC85uQWJ8FLnxtR
D7Py5xmTjqAQOvRUWXobINtICkB91KfwPc87woevispddJ4OgHGLqE5QWC8RF6JLt82cvCrEsD5n
OIZtUEHuxiWASObUUlHlc5iRjwITZPtOTZJATwag3J4Y1Fogqvptfqk80XAwiF4D7a5+bAcs5Ehw
FEDKQFGuCyn5rnf+v/nHXDq1RQ1B+13Zb3UPLJcRDiyTLG5+yAqUUC6Pm+sKEEbpRhb1MGnk1zkK
QzeG011iV/noyc51e+oxJ61cIDn/1UVpP3CJUZ6H/jB5TbXZ3sr7L5JpGOrFEcCBrUdaK81A6GBy
k8X9jtpuwmhcsTFLW1+B1q7dwB1wCOJwrzytX6TpJv8WlbkFFji410r+SVxsrgag82C+HuHS5hRM
3ivHzyymqyjF31TiLBME+QtuGwOJ3FZYCRGVu9Ok7MTFtTNXX9YaJUiq9d0pTPHDT6dXxleIfx0T
34TIWcrFzbj2S0lwKTcRnjTAVsWDjleKmabc8BrUXyr55s7MCwunILrtUodq80e1eFSMoleQpX7g
mmy6SPTFzkhyXwCMImbu2EKF5BydER71YBxOKrb6FSPaPdWe/Gs+rJbG/oo3l7A6C/PepPn1rzYX
oAlkQ9kNqLGBie9aHh0cpYoxJ7c/WaJi1ryEKgUZpjr1LSFiyyOJDM92oI/UyXcd1ESqJIQIE2wq
3rDDEyoGFAeefa7iA/zigsiggueS0jYvKBgHMZZmD2LSOEmbqhiL3PSJpuqu0HNI2iCVbRZPrtf2
chHFSlz0BTc+iWCSQgaBbDT+XQ/rly2drmu6s8LsfkZE+oS0gd9Nh05JmfizO80MbVpH3agwWWvL
hmHfBUuTKraBMJB4U4qoziezqzcYKorQEWQ2m9DoMXuIsujAracMWpWthfHSkHOumat1ZOKQ1nED
GAJeIIpeeAge6HV66fJ2/j+/m7he7mFzTnPDS4KjW2OnJ6DZH4n8vNxKH9Sfv7uGK5JZQ+vRGhfu
iehYsCnz2my9K+qrw9KFjA10RZViNeUztb6w79zInCQoM9xV99o1KOGYWzpkS395NBFstG1u0Ogd
M5ajYezQaZxK8/cMOx0qaaxAHk+ZSRqWBGED3my1abUFBPFuWqSIrWySC5oF+L02wBppwzYXii5b
YF39gqrgc0kSReBoZXxEo+VYcPs7Wc9Q1ysZPgpV24usYUY40gSIgPluXziUwQKYMsaE0i+jMo9f
zFB/cAFf5kdlohyJGyMnnF6Gqt2RRsWpXvgcxpYMFdZduYmHOzmgiNX8JHMGYN6vDG+QY2fF6sca
MG2q/1z581yoUMOZmWkjiN7pVFZZfNOFUTcOI8Ou1wRpTGsk36UK47OqSZKL/TpX5IUDmD+4cd00
TVI4OV2v7VLWDmDHDTK5ZFmr6tsElcoL3wk6WRTfv+/QOUBSedmNUq94uBioyLZPAc6xzJKlUsOs
Acw2QMplMAhSIgUaRX7RufhocPsz+1KsJ4Rz5ezQqu8ywULdFg15QX3s4Ph3U2WI/ABonc+QPlFC
zODUTSVuH2+ip/xDJWl15stCyHaJUv479GPM6q6MckUuhfJNs3wT4b1ltTzkrQ2b35skR5RQHIbb
HVb602b/wEypPXo0w3YypgyeZnj6B1i/5dBwVECoDPEc8+EEUyacFXtCGB4ePpBbJaivFLCEhcYY
qYVfYZq7euIIFVmYRn1hNBbvr1ZI8d/RFt+hvSjSTLFKJKPOxzhGgGlpsH0XiWSAb2a2kFzutsOy
0NT7Y1NxHX3ZrTa36lwKmeGO+07xtKLhOOqzU0QjqmpZe0d1lHnCQkqFqawd3e6ZkHs5OysjDW1E
Cton8yaJOXwkr3ufBgFvypMucDHg+dlb6uNcGpPvkp9pA8y/XG3+/A5HndpqS/IPmwuawBH2RKgd
9PKmnFUqUxgSEAPcwgmobdV0iLhVW1u5IvzXzsVoAPrPJgt9z6/hj52IkgQ1bXkRtZsq0wSjB5Wq
cbMjst1jCuzjY3+t4Bl18Dp5unvcZqVzMePqCRniKohyAr1ZW0hCn1XA+ghI4vY4AwTWFnXthBEp
DubfVOKPrEhtw8jhb1sD4r9W0dA7FP+AaZSbMSWjEWoevkSkM3AJXCbSi7zliwHFxv5LiwxhXB6n
d/kWJvRUH1X+7eY3/mtRDJnKJDbAyz0raWK4jHOano4B1DXyZJVZZQMTqvlQ/GRbQUAlMQERDiQa
dDs8b2McSDNPQPRmHRlPkCYDicW9LGda2Z159oJEHEWi1wF/9sI/Uc9s4okJxzTr5/058JIRkbl9
M/HEBUnWrwW/Qwb4NGZGIvbzRfbGZ1NvI4U8dgtz1EvyfTL8/XJ+M7xhGFOwxSLmTZk9szzz6Utc
1CKxDgGu92XPn2Tw9HjbaIu1EEWSY+4mQf6Fee8UFWxHMmxjGXk/XoB7bDKcoxE90R4OV6lu6Ijr
q/3yYwH9L8JJtQWvS7oqwsl8toKfVtrAgeSrh3qw//7ciFRvrSBjx15RXd+ZvOOw5AfLgAIhOouK
py2nBYFuEgQblUK/uUywjNJuL+5Vzs9nuscfrIwLxynnxFaMOQquIHyJcVr1+qZifBUAjwo2GGFn
+qw8Pl4OJ0EPS6tUEzGeBT90FDMs1vtTC9NGD1Ocok1SJWWso6eBdOs01jRvrMMzzK1J7Q2djgQx
B8tWT+AMGvnDrmQmkStSUI+wgoERQNEKscxCuMpvbCySQNCvlVLHFokIisn+bqDNiJMnXaNRMfiU
E5aG6H9QFEHmIB3LPQmBKLU+WFYM3ANNdsRn7vd/vgfF7WiGjmSWpWArx9TtREBl0A7HuT9B5eUb
XaCQ0U0kUHDBsGoRbqHWF7KLtzFZCNohY90995mkaI0OC6mopBU6Gf34kc6WTlSrYHzjwnm4qHes
87d6LHSidkqEcJBiBk+ljA3dpi9ihswka/+XQQXlnTpGzXD2no7fj4zp6HeB09IaDF+3OlRxmrON
ETvAMcj1pC9m+bkoJm4Tk7kbRddpAfRcfwLpKvb2O1dMQtidY58q9nw4FB1nWsHWtNziwtjQQcer
e3fjG7AcT6YlbjBwO7cjk7MYrltSu1QdEYSHS1M2aQfasOQQ8hhGNogU4KRTvTz7rM7ZpPVPGNkA
fqX52VnMOdHb0nkg4EOpEg10HnPU1El1yv2ZcErrr9O5yfMwDZhQl5naaWp2BLIOA68xCKVLxEOM
yVhA48J+6wSzjhUjl9VYysr85jbkCOLEh1FYEhd91tiulVwUpJmTgSrxXs0qchZTWEB69Gzn6Sc7
IsEmiC3mbRcFuJCdgSwvQNsoxt77ASsTeEbtfDGgckYTRb2CLuKtUBxP2EbD2T18zUGu0HlKI9Jv
9wSa132H3y8D5xNfYDfy3lT4LnCKHJ1oGQIr0BwpQ8MiQ5+GTDu+oSLFYwu/H3oHGhPEt0UH1cPu
k0O31b2tzTKAFkH+GFSAxHLZBGGgIi01PWEtpGu5JEcPfvXBPypUyOqAlgBax8Vk4yVvc0Vc/0n3
74QifKLaeHMSY8Bx5FzhA7e3fq0NvSmOIGwrA3ZWbbLhMeaQzRCkIBdLqTnpFNhMlgEQpcdfksoo
nhgnL8dU2ktpM1Q0tg1tZdTrXBgA9EQ+35v6WHjgN19MUuG1mbrBkteKkDPRMCapGu86jyvLnA48
viUgvVszr2K5X7V0WxvFPaTHP8k54slcq/algDq3AaUzXvFYFHkTP45diQNsFSUgEmGR+MyT4AT9
cwLBGuQB17DA1XF94enD+GTd90Dnoa7GvVhQKVquGuMFKpO1Df0TtSR8K0JkrfIosxIaHbFRwb9L
91KPb+Kt4LaXtT/lL+ZtUmefG7q8JJh4FfnblBqi1ovuvynY5BXV0iQLUSvAx4RnpHWqH0T+fgOW
aDJQLw9jgU6Hryn7Qc1r8Lxxe3p2bqEON3cXs24xsxFIO5+LigwU1AUIyi+mpB5/VHaLmw3vmKgj
AGz0/ym08KLT/INHXsZlHF9Xzjhp6UB3f3lD7Lh5tSE+OAfOXEUMYd5xTrrOe40uluDdaRU7AASi
+cPKqLbw+ib9yBIKi6bYfOR3FClHeDArl8m/8nlG9Lg66mAzhxICNW7ub1XnQRlQzOTYY3ZdWNH2
p9iY5AYSuhT1RChoZSQDguI2s4ces+oQL1wl+SlyCQcCsX7iq6hD8tgonx7p37kiNfzSn1LW6fch
LhSjpBpzcJhiSLUd093gDUhYxJjpEoKLvpFh3uti6tlIiXAxq7bpRMeJndcJiMoCMeCGssRQcA+/
Sv00J4o3nfRLPsQWLgHXPKdmDaiZUiiqDBF3Pp3RVIq9DgYeO4pCY+E3rgJ9CcpWiPfq2Nno8Fvm
xwd4DQOo/IhNA9UxiXHYorajICwPhUvAmMWcJTiatKpsQyTOd08ziL9QwHrv8VFwwmTgKU5GfU0L
z9V9R+I2Tf5z1UkdjAZ738Qlg43niOeK7i2TGgDyBzqagpq+I4FRkIWTmnpor/hlnB8CrXMO7bjL
F5h/txvPQN32LS/q4GAO4Z41lvZwUMQXKLhdyV8ht6DG7GFgkZMLMI1SIFqKwW+6I5RuZrjQ1y2x
JBWkFH7PXE82CqXdhUk0if6rMlz8PL8eBVdRCzxhjB46POs81h8HLLkAG5k4JyFipKiYWwJRndX0
2L/fUPUdrHqiCe9I7jdN8TliatppvMIeBiKP5fFWWLFvAUULZIQZCs+dIA2+lGPWujzq5EkoK3QZ
ebqDPEz+TjRMY+L0SV+3pLjgXRT41sUIL2kCN25IDUCOODcVT9HhbWOXMf3jzAEZPIYYIkXFAl8K
uULpA64shhZcCWiA3Mwd+h3zISJzUulAwzwOjHTHhZ1AmerrK4+DaxDDEBhHeYDmbFa0kKFgk4cH
zXYDfh4GIzC5vc1QmbZm4bGUidox0a+olm8n1wMlNQVLNN8OD4JTRLGFJ+dQUrah2iwjuAFAgQ8D
DCr/lXC1c4iCa+msuiLCFZUpBdhyV7LZPHruLQk2DrrxvuX1ttWSKewCID+Ubn/xTCZ37hMcxbGr
ptOj0J9/0r+W2zPOomLK2rlVJaZHz96eSkmnv7a26EhFvrO+7L4oKSFumkb9u7p7ag/WoBuDYghZ
nXXnprBWgGF5WIQDIRrdip0c4umqhl1ZbQDeVLBW046SL3XdvNO4d69i4i6kQoy6kv3i0d9YLo2/
+38Nrx8rbmfhLXGbcLcIWhoWbpQFmlQg4LAjEhy5qJq1iQKgGKQvF9NfebTGgTTc8jWyxZZtuehm
4flY3a7N9SqNuywJhOXi87uNriCvnFghXttrG5aIist7rt6fZ4qpgGqPcDGP7RX4yLKA3fN9uV0l
+sRXoTJsDLaz+idZUKvq4ZsXHx0Km2WkHvohc1vWMq8JB/DnUMokj45q+IR6oTjkzKq+P8oHFPhV
/8g9yg4+vf97HHg7kCtKBLhEBrOjAXmKHbeeyNTM9WDtHPvq3Jop4YqJ13uuepOIfkLBeyvgmg7u
cbjPP3fwqzRpj2FhK4vo8Mg2t21UlKYcrXbN9CucIuKwhF/BZBt6wxuHyOINsPpyCYuLKuLXoD3I
ayuM+RHzKLBgYgxJcw3X6MHcYo9JETq0ZL2pEEWlixrLCSslffH3ktOvwGcQQNVINd35tWLfd9rC
7cWNjEIvhAzZya8X0mDrT8VzwLtW++zSHbWcd+S5BWS79oDPwF5pNdXvshpxzmMokBWyqgKmmGbU
0BIH4RjmkQaKMi83Q5mrJ9oA1s+9U3gZVWNcr7ArK8XuqNiLYo5c6u7NHop/qLtdp3UpM8207Y5E
HM0v90Pz2DbMQsHoh4HMDxCM2pfEwuwOUewhKJTg6qcx9Xqp9B4FpYmtqI6WONM3LzliO5wbhrxK
ROQ209k1E2ODOKInIpoWpZ3qsmAeb6891gcK2T+T80rrsDMPKXFSSFEib4PWhxrVPMwoW4mdAe6e
wSUeMFqIJXEIQ0wKYhwfdu3Xr8/vyUpwzz9h71Dj5GlHG3qg++BOlOELir8M3grx3ge25SVZ6b22
Sq8Fh8gNCEyMqHG9qwVKku/dlwoIj6+oWF49faLNB2bh0r1ALhdllWq8qeLoz681UttXD3MRadRe
G7w3X6OuikrGpvKOeVNzf8PChNoOb3L1JATE2j9W752v+LxhADazvFSEuSC22lMJoBs2pWrU43kc
YgYIrpb42SyrIx1y55K5JmwuHHnyzIHMCpGN497RFR474LAjOB+imQGt3P0q2aXaNdazFGIWzWvy
LIkCh73z5256GKm2bTQFl9ednnhEu18r7SCx4zrnB9N5StFOT718o5/CnGwhEawYoRIUu6eq93mB
L8ZnqrlOG9Gv+J10//XP2Oupd29HdydOLEOlnmY6h9cRAiT8Gjp8vMdafWWDm1z9kJOPmIXZBQOj
pt2TLM6Cz/yUl8uL8CydWSJV3/Hl2myk0z+BsnVdvSFXneajngWehpziN01ZHSJaPCZa2Plq77Mn
c2BgP/MZlAET3nO18Bh2+h0opzX8wSesv4NYWtWZ2MxeudGnBzymODJVShvHiwW34zsvWterlb0W
dYNL2ZoZ7Qn2jN8DE4l1JWXr/UF1BPcH8ufLtR8ajoExvUHn4o9jZOwOESn53XUVprxiWSHNHQzP
MxYGLfouCD/6K1CGH+Ycc9ExFWhx3Y3b9vcLkrBNRF2Gq42GRhkUA1Mz7NrLBnhoPi26kguzwHvL
9va/ZQVMwvai2XZh4qChmWEl/Dgf6JcMmktHMP2HH6WHhSSpFYkTNIK7g7JBcmQ3D0D/Vukwb7fs
1pGNFwwgjtmb6mim7sXt1Plq8PLnO9ilO4cM4xHZhm16jegIONxdh3Ttu7pOt4RRnbKNkHGD+F3s
cWWMZdMFsHmABCHCLAtYwkeuUEhSAhTyQfBscZfNvVdkVlgbkqUrMeGaMZE0jHItRjXOGQPhtPtv
fHHMnwhwmSk0qXIpxlVVcMIPTp3SFzXRpdWH/A0q/VAaKs5t83wNc8tVqwK3hpJeCx5QgvHYwmw9
3Z3Vga/ElylTfgMXhtpaQ+rP4jEVRuNX7FuUdIOEDAqJqwcMOyyExRi+lRpB14/7HqNDPbOG4zyo
39rcNkkLlg+j4fFqtIvWXwPw1fXZ3D5QyLP35iLEuxcrCWJemcbvlTFhbtAeMDM+fRZ2Y0/2bow2
RICOTjN5wYEbKapIyrHQAQdNlK8avzdFi4VXxXu4nTmCNsq344yY5pJUC76WnzjQ2JR5weh1qKzB
rIUEKGFZ2RHeh2/BiyB5n6nAPNIDJdNROA+nIjwKUBEkJ20KXTWZr3pscQFpPAHfwqLJ6FJX5NJ8
4MjTmFJ9p1AYw0AE5sR9DOpYydspH/Fe0FsFCtRjNNnYdOaUZgeIsF2CM7mXarl131yWIhsKde71
guRb5Es1xbN8gv6tcrgrEExcqChuKLA9i8YNlijhG45g5rd7YPWFuc/H13Bw90EVnjTCneUxNKma
/WGXkX2wokVabf1VRNsLFBBSqtn/mDxru6exNI9CKU0u6IywVw5NFEGh3h4coaa5TVGCB2kcT9ym
4jolHPRy23NAJIgOPpk8ObAivDU7r0EbKOBM3rdYJSHhu1eco0pAPnpsPpkktZ7+ODQXnRsRtjiv
iAzZez5k6rolanM+qwk2Q0Y96Vi6u/1VuYtOnDOtyN2g6goZcyd4AsymGI3p+Uyhvt5kjaBq6fwZ
Ytq1Dey6G3GRgyq4gCV5BA02reOx8ixsP481CUxxkK7Jnl+4d/5BZXrzv3ZaKGhTC/iuwpb8FHDX
7RgL+2tzNhHQ7EtE1q3fgSVw2SKMXAf/JG1zEI2PfeAeuX0YRmQ+c8fHKa/JyDt0RqnL4487crbz
DLqp13XYEnpj99zlSOx9dBl3mA3KxtvsjNMX2dmAK4fuOC1Pxmh7lHx9ZuXxmizwkcWnGX+/m7Id
srcf03rRmNWRYIZNiDqapETMug/kzEjMtO1T3boOr7HUuwhBleTWzrQdm1WdTWC9BuzAMD+Oq7Nd
oYN2e8hsJId502auF0RiMWDutdlY4BHqmq7r0cgbEfV7E/rU48DUGu1lJsGtu59+Xmqvgyp1DvF7
VUKO6hZKzHPhagP3LhR4nxBUU+FhnNs6Lkc5u06fJuTJiuATgi2BSdv+gFlU4YjoQmzkDIJ5O09d
hnL9FTiYePiazGKYlIpQLIGU73Ab98MZ1fBlFDt9s4ezy1zvr6bjoH6DfAMIchKvzanakM8VYa1D
eRmtzH/2KzKbQ+USGXp5AWMKziT+e0VsfQQcGrt3yj1KiuR+797AAeJfW2A/ttrc60yws4k3OtpS
28VVjriGgudDSbH0OMV+pkAlAxHonQHMWM/HuzvQf/q3AfSwoy9UCT38pGLcVUwOVm0tpTd5QcD3
FFoLCKeu5+UjVW2CJkjKQCv49NY+nueFOucWmGwXNDoWgUn3oksNxcaajf+StetZ/bQjszz2daMN
JgOJSIZwoziWGUr/8aVdFv+S0DPI+WvTVCIRl0yco/UWMGAlvGthse48HGiDCuCi/rj1mqY1lm6K
TD1ZZDsEI+13P5k+1h9uxI9yE1Dvf2ltHBKB9ZSz/X4musn+Y8OVBm2CkVanvXi8zZL7dK3RthAl
yypds6Qnwe8M1Sa8lde5g56LuA8cqW4Ab8yb2dCmMsHCHKLwZuAMCmxF30uqnm/w+OceGHQ1RS1T
Im1rBZ62uZ5oagwxRxDjblZNgEHPA6B8F/B/FIV25j0CjRgX1SA506Dki/4ejN5x/EsedUZvq1VN
Ok6H1fbu9x4THX34lDDTC2IaKVwUgN0M7MlMM/bZXgz0UpxcX6kdhkJlhGh1dcyUGfK4zCZIP6Po
G6yZCb71uNLwI0YqhkVV1ss5sgxyARynjW1QTcGgAaWGMGPcGkzBhyAVDJSyjYjNOTSDlw1i9law
QYH0WtwPvAhbyxElct7WhWt1B6d8JJzfCKmTVal6HOrHYO+33TeN5ghtumaynPrcvBfLVJ3/nwqO
8hOL7EpNNt+7BrLVWS0KCpO0KU0KUN3xXagBOtLLKdNANnr+82Chfdj7lM2PKLtQZAF5mk7JB+5T
gw7BBe+z9PDPewJ61htG+WCE35l1VmcEd+U8xZrSB+kL/eSIB3xnF0+DBnQhYaFjYnsiN808IqN2
aluhuwTy4A+/WmOz7vzg0a/JWk5MmjEqkCWyiVih4eyrp38mvqvshWQn7B7DkuCPFNW81fHgNFgJ
S8c+UtnRQpLx9xhjemiZJ4qXd2UKOLkzwUV1MSpifyc+TAhr9yCBGgcaY24n0BpiuP11z4rNQ+mb
UerVBMTXlVOaq2NTyKO8kJC3DJpPjkzNGwBqEKpavKsgnPnMkcqijLNgxavgXu4/prDF8oFmbdn7
DGVqTKq3r3Fbtk6IkOoK7VEtM75Bfch6Nahc03fAz3Stl7izSJIp/Vk/nMUuMEJgsPg5Iwdwtn//
8SkzuF35V9Hzg8eUvz3IJwIR2DeqJUHd76gE2Gr70eF/NdjsVQAwr7MWnyf07hfg3ouwZeLQX3U5
yIEGigNkAYa5sohsmXZg/4zHKei2rEgY6o3dh8XpdvGT264aUPsh6C6o6o1bjwodhinInKHKE6lp
ptgSbH6Ieg+/0VZ7ulGrM6ierlwzhpGPdX0g4EbrAV30T3bhY2gjiJtyPXshv/tS3/UamH5+XWYc
q5Y8Kr7RCwC6z6j29oUST1sQNGdgCYFf88Rndpf1mA5rPBhucqJvQs4k95CKXBd3FIRUB3wlEhU8
pTx7QHlYlsZ9zTGPrFEPNS4QT7JKKsmXm8qrOcsdDzJfus1pZuORU/lISyLlOE9maNF6FXzRaboh
VirC8pOppIV9idxEcg2GcGE0ePiS2x5BRxsl3qxnut8cAC49TLsqawr3C0knxvx1Sp4ARB4edck7
arjKUs4VnfSIQNg7XOUDtC92JZvHJeorGjbYW0ghGaVwHAV5WJeVFESu25bhra82iinFTTXsLPKA
ZKDjlGAvPIlSFv1Jx4BoItmhFbg0YWop17UnPw5dMkJRfadq3Yk0cj/y9oqEuIfp7ZsVSxiaHCHT
+VC8P9UyKjq4+pYue5nCcyTNhmhsb+pNPmPoUNX8m3DBi5ZAOHRkJeCu6XLhCq9ZRyX2/4iESCyo
ylRFVJ7C25/A/VMND8vnicvdHTNJfHBR0eh3mind6qAtYp96nxAV8gKlmbxAZZuqigOMatdnP9DL
M5+6XysGkkpOX0rZwAygnVyMKmgWmK2FOKwIorGn+iWV/zMHjxO85pJyPZXRW7ABaIX/tMiTsQ5J
RoO4ZMi2jpGBpcMnqQDravszRfnFzIAvGG5mI0qAodkddxujtNyAoa7uMlmr76DEHGCtrkdBxGtd
sfPfC4K/Bb2rJpZnhxv1ZN0IMJP7vsEQupnJ/7B5hmorjsLd7OH15L5T+exQXZR2OYwtRcu3Btbc
9esom9DDbFIr9dJtd7R0zb78Ql96rVYEnieB6sxuIzrYHssUNbbf8MLyfpkpvJGA0RSu/k7f2Hxw
xZQ8ymupsK0rdssiWfMq2n21QY1zL1FEFEPl+mBoyRixwn9btTKYPFMUSJgwXftvHeiO63oX4Qq1
N8kTqAUhm9S2kqlxei0Na3dNg1A1velLjvYHpt+R6ZJIzAhr0xHm5DL8ixUCOYvTS2xKLFMUQ6R5
3UXNUjrfS22e8jpTlMs8xe1Sybf512Dpg73UmtnBlilqeUmLnwfatnl6mLjqSuqE2Yy/VDIMgTGw
SPoL3k8sHn91kQnvuyGqpU1nZtRMIOW4WStxvrJkWy0ERNegiuS994T0gjPxjuBIJyxFLME5agVS
01znyOkVRDXawwBaKtmf6FPhX4+6pbT/Z+ZW9RIP8IYk3cNKGSDkBO3Oz1Rt5go7GLWhk8TVC8a6
g+RLFpt+uZbtdXiG0f7FsYLJvhq/MmZtDizOi2QbfN1Zstp/ojIOFgKCm8eVU9gSldevxxtwHBCy
/aAGR8wehNfhvxFS0x7cIbFfOrlQ/HdA0jby9R0E1LVbwn5me/UhV5Q+vOaw5gtyJKHDEunsxhaE
t8JVMjy7nANoq7a1waeLywKNgoVpTDe/wlpmBNVFtKC12t8Wo2lOmefVyiFTgGqq3dxEt3nY0heC
tmqq9F+W583oBS2kUz0Snn2UCcy2iR+S6lc5fbiBIDs5qSms1u1KmF0sj+eJDKjSKn13ud+aKiji
CHmQ73+Og6XmRHhjtCeXQnNWsIhdWqsLugozPpgJLVn0iwZ1kJyYNmxhyCTBvKIW5gMIXQJlS/Wq
3TkQlg6EPZ23mRc/DCRCDMSkHbzF84KHx6shTJPQl4RfAt8n782aqDE0rjn8Lm9iZe6GtzATCXsm
+8J6TEg0+8ju5nw1JpuolrGwza/t2hwO78cfUr/22ZfAeMhe4FCyOmnlI928/5HHkm/wpdXIOQvt
MLArjKW59HBVrLW8LL9mr1mInaf4kDaX+t9lwscVBKuxL3/Gw5/CERqcohm45es4lxyzlRjDX97V
vFswwYyBqsCpB50XY3L7dRebnl6ejZEcXATM1Ss62SBlJP2JccyYDm8RFILcf99OTI2NcObNxdeI
7WncE+4DPPm0wAdkQjtxk2NR5AxzNzwBj4ITJm0saFqzUxy0MIeESheTKp+GPabokNCWpwtvBHRI
olwFsubpBAJhrD/PksXVkYSymPzO5gfcdUVdcJL81HuG60/sOnNxGNj5nwnnSLQ0T5w57jYLyfag
UryYn2mDmMCfek25yNuEaLTucldYvokuJ9usVlAlTC+l+elV6Hl0OsSSAUNuYp8pSz1YS9LiHUJm
bcQud7fpBO5N3Nud5YJ29fiVcmlV2g+A6t55mAYuh4wfrRK67LUEbSpRXxqOor9udWQrsENZ6gi1
9JMeqT9ITZCwBdy2EEfu1Z9mRnGzxbVMW0l7h+ymOKbTwARt8k0ADTwhAuzytRF8nRp3YwvOolZh
ebtsfjGVahpdQmjI9BkDfdqFLp86YRxa4cUyPoPVXaTCp1ZwSgHiaAkyFmLly7tOjGt8hUHJBWrk
Fdwr7yZ+kYVdU0pxdmhCD7+5zqO3ES5m797gfRYXSRNyltzqVVv0n9AHgvpY2w7967lVT4hnzKVU
J/jT+1w0Pb91kW0Sg0D+9n+e6eGKRTCkt06hRDTRKMkFKFyxWUVujqSjJDCpcU1sHnj3vpinrD3V
s14PC/T6iyrfVcP01nI6aTs+PIffhwvYWq1gR0R/atNFyafp813DZVc6HnklRYrFiPT2mHXsXIzB
bLYhkog6e6erWNDAKKEXvj2DkMsDg3B/VaKjrbGzHzoW0pxS4cG8EJAl8+Boo8duO8ejYP2ipl1b
EdzClTauuYw2Tmi7hE67WJZXZyMbDJK+gEH7e3mv62NE4V/4LoQzwhbLW2LH3NZnv3dOBktFAzM0
b7+m9D381cS87lspX6IpRZ3z3/Gk9mqqKGys0El06H8Fl9JG42oLoOWUzPRcr33a1CdrPK79J4Ec
zPQG4/asJZtat3d5VNEBca0qKLvy78ndOK8R7CENt4D4+iyYVzUJhD/qBExFkt9Bl6lOFdP02fEs
Mhb8auTRpcEtGZUS72FQ3Ss0Aki9O016tqMRD6KabIr8MISBQ86AJlS+zXkjwpqXRdjzkfWOj1Af
P5O2TT/cHS0T3zSSQqd27l4x9CVbZ+XDjEQyqhG+C1rvwITd9jYpXplk1l7fsmFZpkEwt7bt76NE
O7R5ciVYwiuuVMpSgiZIVCnXhunzZmb9snqB5Upm1qlFNqvZibWjFSLq81Qd923ftW3gke0tx1Up
CtPeXVmysHRnuXgf2f8RaIDElaYLUZtL1AJiZVc3AcsZ/P79pcKI2WMLbSp6U824H7iVL9OSnVto
aukX2mxKdDLzhz2asi42grd5fzgD0JbMT3RiNfJSNJg//01UP1t09qhHJePKk4IyViSwjyxauO1U
sJyVzrkHrxRnmbeJpcwZ4OGY8epPlww4PudXQ1v6AGeQ9dGVI2oS+uDLbo5FdHP5aZ8LHivyNAEk
KOrzYDXFr72U+zCWBmbGHxeeMk2gcg44gyGeQs9aMBmTyyOZF2gzSqb6RUDEeL/2paLadexYNIrE
pMag5e2sm8uA77DAwjOtX4fdLpwFBiT5Byg505OhLIMfFHvIptQ0RSq2Z7FmHJw/pb8UgeZDycKp
uItUijJI5qjEINPkMWnjINb7KeV/Y21GlqydZTTaKztt55Rpr4sJoVr2xKMtfI/zeZx6pGmjilD9
bGfCX0xzUh1osPBwaSO3YKyoOwjUa1uuGA1tr/oPQuPZIc2311RjWFANHRf/bAHQaRi5atweB4lY
DY1dyXFtdLChz+p49ollum/Jb/9JjjM6Dqm8NWrHYqFSPeuOdHF8soMNWho2KlYMomhxFstKsy7X
SJuqlUhddOfQrdNmnZ4/5j5D2ErzBs78xLOJ2Flyt5HUUXkCoCWrjKF93/aKFPE44zTxexga8ndc
ZycS8i/4M9WoXGe11HM5AJfvQg+Uujz/2PAQ/Vy99c6l7+PYC1CX7fIKqHHDX5ZkkUTbZy98C4Oi
f4UwNQ+QA4tQti62k1gf+aIZQtKStr5qt7IVBTAKCGWkWenYULA8OW+/yOzM8vr3F8ZiUEtYyMCZ
koUBnwQun/ouqU6PK66XrIak7aVYCCjnI85c5kTyXcRPkQJwifK8bUBjzI5FqO32R7hdpHivULQ6
aYR3CgOjeDiveCeSj30wmePLRh2VTLNun1OJoQ3tQGX6tnKrmhXYHOJ5oRejgjmLVF+KDzNhUQ2B
sf+GdUsvEMKhGQ4k9arjnMlQQAHYQ6dVcPfZmN2u9hUpUthZD5M7EbY4oAaxbOxx9tjuxv69XYTd
bTHSQikeIcNnshezPDEa5IQW8EP2hwsQXbFQswE2tfjPQAzW9F0sAe6CJD/2DI1+fCWHgBwcGvMS
HXfp4N6Vkgz/KZ10RZUwyqDiMvVLkRpcM0RmxH2lkCLqQrqVbZMqg+Xyy38dg+HE0XXl6yRKX7mz
6b2Fe50YIofE5TFyFPnWS/CIwUsRj/+b7exAyH6xFuqPfYu6c5I5HAkkiNwIvn5iPbS/M2Pj6MU4
rggwSJrQGe44/MkreSwfxbbK54iUksbOAxmW5OvfO1mpyKkn6wGjXpT0gQOzh7rbnWvUa8rSj5ug
EJgYIR8NKY0tNY0KgLi+X8uaHjg6p4ZY7GblsSU+TcId4me1ZkXZfFaB4sBqfOJwcE6+YcCtS10r
Kuw7PjJIR/HN5/+0Os0qJe2yXWAK97mvCsHxvQuTKbY51E6x7xj2kkQiPVm0Nva5urBW2wYBNzJo
NjSiQKzw9qdQwbRGvQJ4lCIPmcgUJDA1NhbWjgJ8TPkrO5DdHf9haXgS6qGAlNEDmkWKJyEA5oot
GY4JYIRkSNa5hW3wMJkZvzqXbKhyd0jnLmRM2AGT3D+hcuVV4xxnxk2+mOPezP6Hsmm5u1yik7jS
jqnW0te5W+Nrze2wJ8V4BKL6UVEEL3DMiE4104hLJeHwP/m6B/TiaFk2C4RYAJB2NZje+2n/CbHJ
wJcxT36cqd1IvJqVlceLODh6kQLBijW3zk3laTmyNf2GrPdCN3Q6ImuWrh33khS1aZuMpl5HL4pk
m46CQ5+FJHT7aq0RUqJABUdKLbf50H9qZVwd1zTPVL4CtZkUSx8+IY909rl/FUy1oERM2Ash30nj
PEfEJWZFzzIrL0od/eJymaEynQ4KjLYsBMahpFo/byW82wgwln+3N+nzXYKb7sx/bMUAwP4WK8z9
Coi/ZdosYiL54OkV8dpn9LH2QVub5VHPQcY12LhOTQhtLdg3az1w+lejP+97Ta29PDxSFnGUDzg+
Fp5SY3PbsDPZmZFUPjGiWWrct8GcawoY5goCXDKgvJw4OjCrvb0G05gDHirYaR37WrxeIhyW1Gup
qPe7EsxYT19yBi7wjVo34j1fagwux44mwKOm7s7/1p5aX3iOU4dWh7QPetQNkfBHJZrJpVG6mjB0
USopJFyIuHIRozaFB8WUtmSOkzwhcbl64HXqa42cdl+b61FuTkKRrt1c2H+PbKqtv9BFuwBXq6Ot
WxL+CUuMF2lXhpzSO5DJENV13cIIpO8LHgY+8ZS/EKG3MFaZYts1FrzMrwPfynNQ2Ka2OrqWagqz
LWFptCySu2aZDHepIgGCHy0UfM1pypJFdhKT45Gf8hvyM0O0yP6TaXWOJVctwzbaCrN6dSRrqNvE
wjZrWFXxX4RNWSpNMqACLAkGFcQGcSCbzdnRGXg48gAuD9DO1I5Q2sQKkFN5nOamqDmQvXv0NrQc
2dbPrUspk7JRX0AAwwO7paXSwH0J6j6FIXeUgY7R0yD7b8AE0t/lf5xh/ACRNwE1x+MUcZp69yFM
4VFpzHUxjOHJtv1osXL7IPRVMQoqovdfDSxc3sGGbR4E2xGaXO2WxEivbEJvN2MlpJAplAm/CJT4
uP05XuhRUudlhbGtY5MfgsmuUZAPfCUw23INiV088qB/bxP1gLzRx9LJcKFR33i+qBz6/IASpfpD
NPAk60RsLaope/IZbgMhO/6foniDg/SmtS9407pCm42GHmWjsaNZn+uxXDsKWGw5/UiaDQ+E7kGD
+Vyb2XGe8cL83FyHPAwKFh1n2LV2Y8laj2YLTfGiMS+xbb6D/9Rqnptd41v6ZDv6UCFod4ziipO3
HWrjmN+t3gvk6ajz4XolBL/nhE8EGijQ7m4QobpMnEErdNsviKnW2V+M2Y0hhH796OmwUamNcT/R
V/2WPNHlL1C7tg+kzdot4G8+mgeKu6BJl/Rd9/hsj3+s8BH1/jh15ZyDXBUl+vsGodaqqP0x3dcZ
uRGslJUR8q74uYYUoXv3oBnxClK91o0MTPu6frtP+Twx7X9Ld+s7Eq15nenV+x8k+rcDfbH0KeDw
Y4HyCDolK7uRLZuDbTl30EaKIwr7Ltyp1GhZS0Z9RkTRXVhA/5T6jqV+SwDnCNNuFUohPzVRJF54
h8flv1pIWxCaH/vD+9cyuyatjzpqlDuYWcsL5SmBkL8brzLHS6lAVDCOON7BvSM6yXpiyH2pAnqf
mFm33xXmOjaDnfdkM5rHcP1v7H5GrhtTZ/wVR1gRDGPb4cK6mrsSlSC7L/d+rKWlWVrrOlV13/k3
Wau3WxiKzAjKEYuCuplnkHsLgkelOMP2t3Z7QKTym23gW7f2L7jGiRQpBrl7/efzOQ79muC5HeWn
7/7uFqnK3DueW9HmOeDHMavr5rsCh2ubmMSG3dgv5yX2TbuC5Mwu/cW7/yDwtk8eex+xUCcu3WcZ
pzgbhuri6hqeT0qihpv7PlnHxH3mzEsyH3R2V2J/9jX3qpmk+nONaGk6WbxBg197nVp8T4xjCawn
NV5JUkIrbNuUovaIb3OTDM+PstA7HVwzoElMsAzspFWqZ2mY5b2GeY9uVytpI/e/jR5Ba5wdRZRG
4AHrdcOpoKnMIiStuTQDv3YVND7jyvkx6p7TKtrYVoVPnb+MBfK2GE/AwsOnhScUeA1iqWqygqJb
OWGTBUb2Cpm8jxmXWgpc+PAtQMakHQ9xIeZ/68SCnloIoJoXjgy2aO6baHXKWMv8wK7q71ptNSLi
O+tei5swGZ3rLN/3unl2fDbuta+z34iEpUr0cY4MPTdZYeJaN2ITw91sx2G8jeCebTEKDSqO2lJn
13G7fUAHCg615tjR++fY/GuGqEGXE2pErGUH9Th8I96VQmTtVshGBbMZIM2R1H9JRZ0e5sSmNHAE
7VgsVBTVaSuYeSYjI4MGYZPKRqjgq8bKKWd9P0ln/jnHXaGR7H+qMM9b1sKIJi+3WU4bURW9W2+x
XtuuEAcI3QZ/Nli4mkfcF+mLa/EEny+venX9d6/Msi2elvAm//2aDH9698c5hsUpuBrSQ6o7UGaA
c7IGFxlOdNLcu7Ywhs8Xu4xg9/mSq2yjW0dNW0QykarAC1JTqTbM0ObqA45iBXDQHT6IIkVspY2M
8UTpJyM+lzHNa7D6dU/b+gaQEWt0i9I9GfAyTCphxBIO0l7pb5Vk55mnsiytlRC2TnB9warpOkc6
tmEp+ccAItEfeYkgBWCqBFbrBaqx/U6lePh0vNXtTrPsIj5fOlMo6bCHGfmR6t59p5bSMkE+VXJm
2GZFrENmZtzEsP+cCYlVv2FNx/VWd+woy2cELyajWVqRcSx2DB8LZnJfamvvYGyj3S/7mA+0hXXF
6gFkuOXpCn5sgtpMlT+k317zIxuOVUB8wyJgSKupb6f8x7bM+HzCQPVIVxc3ACMnBoms94/vHuGB
+3IYksKLamTYE5nEopdfkQ8C03N3mycDriafKbQtGU3ZPhl1o+SbbQgzOdIyN9ns9bSd6ZUelAEZ
32ZcWpAAjKHL0QlS9vBgSULglrnEH9j1jeimDKs8kxBhliBohGDZM6v99Ji4F56Yuq4By1sIGCGz
HcTCBPQcU+9OVV1F9kJGi3uXL5s3hHkvs7f6dd68dhUfXe2hbiWkQvlUPYMck4oXdeNB2L41qNsV
pH0HEVmRJZdOM1cPvSNgLD0Nt8XPlCSnFuauE+lotLIE561cmJ0w7SXADP2Y8OzrN0c3xS1/wUOB
6YBr0BFsofKM0RUTUBJLK/1SKyEXfWS8XVyQxHelLMlNZRg7MD/rxtqzgstqp3ypGw/E72q0n9NQ
boWKi9cfL+UnM8bGZTit8SxaX/9PR7GtWIUO+bKCfqB052WiTy6YGnzRPGr/vtF7EWmyzNLd9gjU
mpyYRNQeV0/56q4xc1bt07WrpSIV2SYzrqwSqPU2jN6CKNzS+syc65J6ptvVCUMXcf8tx+PwHidB
ExtJfBy1k+55NiZMXuYIdhSfO7wjuMt56H5MViCwf1xldDEXMUuluS06DajmlwrrpaMaFqmJirRR
XTOZglnDlacUP+w4tFZp0ZjMig7J7vZvwGBlqO1Ax/ULWZfXZA/+yHtWFeVXNJo2n3o0qO8Xy9vb
nXkd2O2qx00+cFjP5vk/dSeBiQubR1BGU2VFsxKTfP7AXJb5v+T+Ua1mD4jG/dpl2VrimH+e0rpZ
Bkx89PU4aAqOWjB9b46rqXnSYCoGcsywZjekdyNlh5Ee3fLJHBKoQglTfjm7aXVdTF3984NZpDWg
OQsw8H3vi64MK3e7vOU4XSnT0GMe9U2E75f9mOM3kp5hLl0vkA4AaKDtPa8ivOH93+F910D5eB7B
Dg/ElWpPnWSfLQmRDpcJZMBSvus+bL3oIH5T8tqHpvOiL05xq7jYgVL+U75d0drJ7zy2GdJXgVQf
1sLJa1atUXDxCeTi5nozKIECgTrA0DLKF6mXtRai92z2yTB0kJZUqOjZLQ7Vhr2+cbfjm4yQBCao
sot3+eDPjI79Cjwj2CO6Kbq2cxsNd8KnrezX1qWAh7QraFLHKqzt3IamhbPed/WpEpa6kafbahVF
HF/DJ46Ez16eiNLTmuZ9MsGPr/Ojg8l70IqzBTpDM4TqsXfsYw9F/GOzKC2bV/N5uoRMiIyfpSl7
EVd/WKoQ+PWsXopcXGEJQq90+DIQhl+UfJDf/aLWM2R+SDGLXPBbSOuEW6mZi7x9BRsKqjAqKxWw
IUD2JNzmp26crbLb9uj93SxJGEKxk1bgNfoZV1IWLYrKc5xMa5l+4Fu4g8Dowl2l0whjSNIfXUZB
jNT1ij3oI0KgG6z5m/bLV7yyw5uafl9yqSO0waCTfkUAvcnGhTgQEB4d6IfcBMvX+tnELuI2IhH/
9uOv6bMziHrQba4BaiKoCRD2358R96QfvBdwfz3+/HXl28/y6VKNrlHtbYQz/l6myfRAPU2DpZa7
4EqVRz3XIeDbh6KP6X5v/fMQrZXARxSduRev+g2XUEyKqxpNowzw7EjL02JFtJv+GCJNnbATVU9v
KgJWqcrj+OIKaNdhYftfkAz/f0wk3si/7iXD2atEE8n4V6Sm5WqGuvnFb16Eoxt4ZKiJ5aAmxu5m
oaGRP2SImALbKTLC8zqmGQX6oJssCswf2WfMQUAUwWHuKiCDBpsewCt827LQSmdsc883YolsE/ha
rO4TJjMzBWXdW2xRSzNPaXLhx8SktB0aIPfV2ttOiWin3S5J0nNsdr487IAA1ndKxNXiC+yN7dFv
05EC2Iw7Oe2xK+t5rZphdphAJR2rggySglJeUCMStmGFQ/KVahSQC0UZ38TDDvbgNTQYZ+uAdRvu
k07Sv5h1y0W/mi8X7dKW02TzbZTDYfH4XIevnYMFpD9PegmGRO5ZOKXYiYHYQFfICQE0Gcu9t6MY
P8TS298PUqEjA2hG9xviVuEQouKs7BCqk8PQVEgI9M0yvsdVoYgX8j/jb3aJniocd3Mrj6czpH0r
Nu17GWRduFmKU2PmIWioQd5UHDkxSwGxs5FV6sQ1HVtpmoF4z0TsY+xSeQOxri+LaQwBiDzLqydD
z6E8CT1lpvEqKCOQY/FMEuXrs/Ff6WYBCeErYxiqLuNDLFCPxhGgIIHA4me4VVufOpjJZu48AinJ
SOxpdd22+BEUjxeg0D8k9fDdZ8p/zBnsyQc0h+h03Mi1s8v1hYUaWakrZXeva6uvu5rQ95tkxbE5
f6aRrF0bPeG7SdmbgzAky0GB5OEtXzE5PG1tATyIS9kR6OtlEaqvIzt8EMzH6p/+ASjgyCySplT4
WmOvFnlYAmCO6cUgcq8MVxe3IXml7YJM77j3AopZ9J+80Gxua41DH8PxFZlMZxdpzXekMgUAsYo8
sjpYN9i1PpiIufcY040caW+GUs4lyM9AtjVLzbGoq+GEJUIuO6iRJFPTpSy31a1n5UCnWMMJ1JUQ
Hs7mjYV/WBT0AtCNrts5ZkXSNhiwiy1G8YJP8UdMeegcVqahAeqWY4Z1D4qaU0Wg9Cl4jI3oS0FU
sWxm7GDPbor2745XtayeM1sGJRebbwo1dL7wU0huV+UOpT1+UaSxjPD0cDipnXArX9AqrQiCbAlK
y0t+XbpElKFDqUtF1msbjammgB17fCQbBGKeDULfwF1YTw36HsM7Rq9M4ti4/q4KpbhmszfEXoYZ
VMZlksCghLCxDHfcp6Cp5pXUBQNCJU+g+21ulaTecii4apoQ0NQJj8NQiMGSgVOfMtFK1eBBv3Zb
8BEvFWYs7CGHw0XLrenqIUnj4AW8jFC62QywVujH2+5WmXyFSyURAd4K0bnmlmeRERIUL2IKdo/D
VOuhgH4jQpAWXAcLP8XXPbGXYydDqbdLwlmUTaePg7CWzEEwboJ3oyufxDjaQhcwZOy2aOSpx5hW
a7ca4xGFqiptKoe863l63axuDzuMJAawI8ZF4els3on8avc7KjU5jvRNaFSH9cBp9a6rO4yGPunr
Y9OyD6W/+WBizbDAayfJe2cGSR1qw0JM/czJBgltn3gz5k8qxalg/rpECBmzODoXZonuBhSDo+Fg
vopW3PkduOkEzIzC/ThB9A1UwaQdYadOh6+u1dduwV+WCgH5X2t5b0ihlb9TtHRRasv36PftcZo4
Pzc6uoNAdtq5HK0QRyiQ4QodMB0AKz8z/lYxu707Mp4cq0lFit6HShztgTqI+USsBT0Ah1fY98gy
wXAkdqictXpYdbVw4Ee3vb9cbPmd6VgWxqUkaLmTGrdi3H57Wkcs4amMTp9nYV+o1+GTcjsvP080
JSANJYchaxfVgk5/7gUwV64M+dixFySD/oJguNJK2QjKBSBnD3VnQA1htwfPIIF4Vh79uUBglZcb
DpbpU1yVkSAVvsWDU2d6NRXe0feyonpwjabSHM91nku3UKdQm3UFOFQkEjEKrSCa50SAnEMenM+B
c80v8IRvHN1ZrKS35QC8mkMREgUoXSDbe9Nu3zPpRwjntnaCi0idErE1O10fy5C98thvQathg94p
eNsp6dgCwtEk9e6egSCehvZ0csr37KyH/BovZNNNC1knpc2N+DFTxxB2RxbLhQfEoGPhENtEv17Y
Ujf25MM4AX/FaDJBByPPmAi67wWa5zGO7S2JOh00LFzZuwwiT2U7fIFXE9PLJikEY0pJCT2ir0f7
OvonwIvRDLwm7oGct3S47pJFPBU6IUsIk60tJsJTOJTVsxnG30IrDcqhFitEzcuUIEkzYOMRkdUC
pQUdcTcvuO5qOhFPsYTEw7wxBEyuMesrnL4oN0DlI3fGIjDCiOTF4ObwCwA16wyjF6XTeXpajc5m
0ygIHXqnMZbZ6FVEnONERTkUos3Mo1r+Ny2w08BSR/98qA3Hc7HB1xGawvA0xShurNqUqUA/zp17
BKat6/wdZxCm0O0WbQOHhyh1SQUhrse0hrwyTQJqzP0CBe+kh4pUkleHwDhmIlqXmMd9LHXp9Uy/
oGPiKgaEvVJHGsLRdkdgerM1+nySdx33fDn/lCw+JH0/UhJX/UrrumxjHlNdOvqtWuHhIRyh3ofd
HKqGlDkiFREkTBk4hAWGwrd6OnF7C7qmHH9soPXb/oBTfHzrH0B49RiOoMtyJfnXdNfYPlAdr9uE
g6iggpSKpaAihbYnZ0H98Lzn8zyJFxNxz8xtqZYQ49bpeoxRJqOJq1KVsV/uKeD2nBQFzHYu/MBl
yZljd2wgN73svt6g1TYqGYMp5dY2SD4XUmjFxcJNKIfsGkTP5VYUdqapau0+D0VI88xJU/Cx3rpt
7m8inus+5feWz6tVwGFgWcowlHFOEmxb23Q6Xo1fZvvhjvygM9N/hgTw4T7gigsUeAx1+TbpHG/5
O3+o43sfpbuBJzfakx23CqJIi/lwuJFkgHCUdXMjLEjQKjfUdOu3NcUh4wIXZGyDnzpzuDYYLqmF
+TAP9TojR8cG71jBsvLS4oWH4Dv0LBtIeOP+YciWAo0yJ6OS/QuZ7A9TvKDzO6WwE0n8Vwtug4SG
H376biCWXH/daGZvU5pgsVBURxJ/tJVGPVpKNEeWzqFjciEK/3bBPklj7K4cg0LOV6+UNN2tQBl6
exJSDtJY1L8pXs5+DeRVUl5RVE7apF/h+9J97N+I/yRtGMNaaSPJMmm8hBplj3kdaNzWSGKjmJsE
A+tP25Wji045Y4hsrWnkzCpEVfm4yGv7wnC7G36Re6QtPd75O7gbgWfm/BnW+2PeVfkSN84Iuctg
cQmm3yh8Vr/Idycw7J3F+fASphNfTGIS8TZkxyLOW93JZOfCcHmBSA7pwuJE8tGKoUxhmq6sNmmb
w7L+fAAERflUvPoQfDpnMJCp5cVyiYgOp42+V/6nilf4B/jP9LZEJuPutFvmR148Vv+VbHZ2E/Jg
F8kN2PlzJUrSYKEnugtTQpJgk9q04u7gmd9h/qfsupfAMQaRtK4pzD9NDLwsfBdujOY50LRcV+Fj
H7+mldgV6Z2321h0+cTcqnKwlYs8whSPNraD6IPjPwDVORA2TUWYyNVKg+0kcXzd2cWC+jcYCHGA
QB6c5+HC4Awq+bokdmuLGqRylOghKrj+gCaQ9d44DgHVnSumFDZVGfCXVjv5k5O52ISfztZRAoc+
ckkS7aIyU+1uJCKovFl1pRK0qjSeC0YS/YKxEUkm977G2qVLCG0DaYdAsRQO2rVU7/1In7OFuYAf
la0A8y1xu67cK6XWUkfTSOhV6PQB0OnDJA30m5UfEHoI6QAmB3KAUr+5U+7C2Y6BuoVMTJC+qnLY
kXBH11PG1q7cA/hlgc7GltSwymJ4kbsAzi/2SQDdFflzeJPbeT+c9DoKlakjMr08Jit1oqorBXcB
cUxq4CXyuw1jP/0X5Aszf9Sf5SHDsuyH97xwPLyWQQZGw51chPi84H25E3poXZfCwDFEfKN4t2l1
mvb71Hcr/sa2rEaYchwWjDOrzcArrXIsTLh5+WdpUZHynLbRjnSciuPE0Gg/Nn08iNqQQz1bZHtm
7oRN68prJhBtgvCVFnwiGtPMRN5aj7DM12rm6OMYNm6igMowzSlQ2bTB0rmYqnpfZkayqZYundJi
6nQgri88UE+2TFNWLlpxQ4LgObbr6rd95rwsleQxtESSnC9oeC6qJMvDmC9nC9/eNoatStvaVYL2
uq7q3Qm4zot3Waa0TuHHVnVZUhqsGCKC1BZnJS3+0eUXUMlFsMRqoHI1l2PmWNFnDyh1zOVKdvZl
t7DfyxSfmfZTO8s6i6iWEgPTo5dhGMFcXlGfx0KeOIe/k6Q05UvSmlLzS7oSHpsbqe2a+jycmZ5Q
y9jVM9/mZp/kVF4kyAFIaMuGLPvivIbZ9vxPeyGTqxnoj/eBT1+AI2Jc8UKWhWe4a8dRMALYj786
i63fqh2E2vrKUunVC69AF/qED7HJWgDDTD/j/tqcBhrT1D6URXHhYjlAgEHVIpwd7GJhF2pKoTeb
05GfLzLQOPHrakbQilMhBo62UQxjmeqMHQEDYnBWY/ug7kFch8WXZNBc+yNvM4b8mH6Vu/bQbiMd
FIQRTWsEnacEd8tXqnjRGRdmKWKdliUUdwWHKhGaDMzlB7GLFQZ3nRwaAP087gbkV6PR+RlVhdPd
2pI2QMKpjxRjYyvyPetZ9Rml8kRXVzY7G5bXyO99D2QdhTIDMdjZr90fPtNmWvWE+qnuBvoTdCQ3
TN3l2uF2CrYFm13oeA2l9YcCkQLWwehr46DOL05DrRTSemfUM2HTfxPwOs1ZO6t4kKXo57n1z01N
Qq3DF0eAZ2IBJRPOEXHMdDnvvAcfB6MlPnuK0dhIGEK9B5dGVBmw0hKcEllROB5RODdlYrTCZxA+
wWvaGC/QWZQZKOdD6e/0D3fDx8gM4ChknKi9F90TvlMANdkLxA0zBpV9gAZN7xlggyimN1td2nJG
e74l571CtoTtEbNQ/HGSwBMCiVOsrCA7JD89Fc/EG3BDoVUWxxuc1MRPnDoAD02nQ04TKeqwQ3x/
MgW9pwW1hqPuZyS+tv9xhom2GI2lctYXZf0IyHQvW/3snaQSrgokhQmd+J78WR32m5jFP0z5jP8V
9wPj1m4M2E3vBPwhdatubfqv6P5kJvAXhhrOUryJOhEglTg5yLn+d2UXly85dndkwRyuaYy+KReI
Z0JTB1hdLq0M3cmqW2ixG4+lwE19rwdF8Tb3kC8Pi4wegnV3i0/SaxjOTWqNpozpMKxq/jg3dHEE
cMCKg9s44593v9zUJkVNkzZoozyi/FFEXKbCgY2wZdf/S+bwXzcuSurUYCeuLwUXBuvRvCNmPYlx
O9MwvikYcrJ0O2sbDuXpLsA/RhB2s2hbALwjtA7Ds8VDoguU85aqoauE5WaDzZWqtXZAi6wGoBpr
O3P3C0O/Rog9XvEiW4Zb8vwjx/gNvZTe1voxbf0lTWYyrXJ0HEl9eS6WOxO+A+F1V4ABaYP83vta
cZHJoqnoaMsqPYKq5USMxTlhgPzTqofl6aPTwz9IKqgGIkfp/g9AS1UfYEBVw+5EL7APzjuwy5OD
q4vfEUJRLDxpPiMikorslImzdMpwvmIdinpLQaYcRtw5LJQ98NBSkdCMcU2q3u/IjIFDeS5EESG3
XVTrNbo8rA+pPRBzPfpQdgQE51dLRiqDtBCfsN/Srbm4E+769hY71njHfoQW/cap4vQw7lzOjDtq
rWliWdYXlW8lRwn8Wueb2PmmswnXobWPBIWgDIIMB/F2ClODfkXzzN3RXWiy9Sc89ZTykNtQODJ8
7QqOSLja2luXqRIrDrqPmDKf9l4DjU2PJay3ZczyxR0es7faofZH25bp+YVE+pSGgnZAaswB7Pu7
JjmJ/GDPJrLKJO2Cmbf+DuCa0bqJmHOl5VPVunmSQ8M3fk6+75sQe1PE3s6wEdtnqET8qLnGvyi/
4ynkQL4q5JXXMw766s5yyf2P7Gm66Y/CS5WBTuOOm7jBv/+rO6EKObQjyq6+KJlQnEkQMATR0KPq
4IcR7zpntPDGlsW6Bon9CU6jeXaHfm8CWEqClBtoQQlxtYlqm3JcfAhBb61lqWmeaZvUaPT4MTVX
s79W9P6+zfHEZ1UDyRpMGMNAVHLWlvPpgVjUXjlwBfuJeaCJZgV+z/c7B51SLk7YVsC/WkUmw2XW
U8FR71ngTeaPC1iTpiNJB+sWU4e7onlroGsmlxgcz6hn95o2E2GpbyLA3hGrmilKeBx35mmS7xrA
TUZMixAt9TPhfAqBngVrktUUa0FvXHF47XAU9enExY/vHZidSRhZ2QD/JfERf6yZYv05AmaP9gji
VlfNmv4hr2/lXmk7HXONyKC8K5xnkAxqw4Vy+0lPpWgy2S3exnCM/1AkLKAtkLPjvY6qpi1kjZex
QiWwPxllRty+f7cSRehgbyAHsDZPCdo5E/i+6lLUKDrEVloMD20xD7JyCOUt3TNA6kM79xawNJlC
rlJPHPPdUrVtlP9CzvWPTXL1+4oAf3B82VC+7mIEz3+rYgz6e5t/nGyDZONRXKeJNgLktJ+zZBXQ
HB5dvys40X+D4b3shvWBc0lijT1Jpdqo/I7eBLXDCDcw5ole8t5xsyW/yMtJtcmED6+LUFr2+xiH
3uinLlJz4xow66R01Pm6uCSMApXqOYJ3YyjKeYfJA30rTzRjglxNaerFuIaaqif+5+VQdp82JAHh
48ceYTnRYU3/UYGG5b2PGynQzj/lEIfgmsoM2RNh9cw4AcPif2U8Xqo6Lbqt3/bb1Kf8FWBlQf6k
nbzKbAj5qpRJtiJXJ7nYLC0lNSesTu0UENlTJ0CUwoh3hD76BCYzVSPQnoKV4UZy7TqP/NXU/I9x
MiWznqn7ExZbpptKSX1X7jczVSl/DU38jVfJ8qNLEcb3M52tJRPe4sqSwSYJBTs3p57SWPB4moif
vttvMajrT4Hx/x8/Z0y3iQlsFGHq16zz+phv/8UV86OVR35vdUClhRvtUGK8e9Wnk0iG6djOu6ao
xztl6dekhIIt4ITlk8Hl6FcBK8jpAi3KYRDGBBCicb1wJJQtIhOKSGMKQuNV+fmQ8yNKzA0a9Ylu
D8PIQ60WxdAADaLqq2u1BU7WxKPQg6O42/XrRiHCVR0Ax6+bPy2ZLB8Z/Irm9WVnLs4vURSGduqK
DgrcO8HlsLPtULqwDDlW3Frk4MChc4Ifyztmtowr8GUa0+nam/ggAxXuU1USfzSfvazqjtYACfPy
CcAQM1fHEXY9ODoVd7pHmiKO41xD1Rumq9oSy5gQr3EcbmVd2ID4tXJRG5wqwHTKZWB+b5JKoLfu
sYDMDy1qinUvu/pRur7pI/8zxs2JsV9y5gaC/FIIEWTzsROv+p5Ub+qAVHk+H6mSkS/N3fjF+9KF
8NtL0tzKvDfrhPRTC8t5hTYHKnkPnqiXPfC23W7YOaeM5D3wVzXXV2d4dtG2+Mmj6UkHPa4DGReD
MM/YwKB+wZwEbqoH591aAZPNQgzc0FqXxPzS9O46uru1HzvRIVjYATx7ahySse/AD5ofAq9VpS5S
Er5XjdZEs9Pe7HUvFkwzbKd+A2sRLpzSADE0enfOiqrFWOYPt8O38aRFIa71aM4OiYduhRiaRK21
kpnHA79RUUTcGWdbvwMw2/wYvQu+dAUJsf1q4fgEV3WU52IvCaw4VBcCR3b0ES04G0yew+O9Wm97
zgBYf6yJQiBtn0kYL2qKcE7es8PfkxCG+nJUXrOZ5T//RjHfmgFaBDDzMtKGz+gJxl+vVTZk9h9N
P6UR8KjyomoWhxAO4ezFeuA/btzEEAfLWp65BiPBB4JmArEORggcA4WHbsp7JMVLHBdGt1t6d9GJ
P8Tg524bVhohupUAZPG1VmuidCbWNsqSHhxseBl+EOu8klFjclqa+pffJo5VuBvzaiLdW1APkDAq
tZpb8jY/QsslyTsBINk02E2bSH/1Z8YN1UW5+eqJCIKuZelAbuL79GswD9vJb9UtUSzNxE6HLnqW
OfNXDapfPXOD7QAOugw1ONYeNNNIBu6eWDu+rHgd32sYoqLA+tzOEQNLwgJHX0xzKAyrrFUc2Pua
HZNDGjwoSaykigmeaB+O4zZ5yFU/A1HtHr35Yk0ws/kO1rSW3CzMyNPiGDqsiNHr8aDVSSuXKc29
CMSujLKJjJJgtUXbHMYF2u1ZMXes78YlmaAaUAzA02u/AMEHeusBLKhmvOXie704KhetK+LK5jGN
+SyO5SzU0wkNERT7Q1vxhcZvdxqmP4IJRfi+mOOQ7X4Wso9yc4ACIjWUtol539VwG8idD+OuTns6
DImszogk72HiVflaN2X0U5IlS4Zxkhe8JUvs4aoaNlGZYRFrNnhlvHojp1kPbNF1fETbml3UPgRs
3vFz8OiAYb+qqajE1+Wp2qOx9Ar2W1wjC3s3d1Q8XLELdBn1Dikx/ihFvIB75TKbv0XfGXYyVPXD
pH9dRcaIwVIhOpmUFyl1YQ27HyHdyL6pyIddmsSyckOIk98u+a8OEFsxsAzKKEEIj+Isbd65RKvb
7twClJkAGY3YxkSSAnkKGF5asjdUHb2nXbacLtOTY2WtUmUKbs2IsTsNWNZQLe6GPkOzwu1legFq
GKZ3hVySefZ6ZrXpXcznXGFWM8nzX9ribGge5ORnMmxG8LYnXG+22GfnvdQkxMMV76QVPHy323TV
BODRA4OUCJrfLrJsAOpNSVHW1pDhh9RN9M8IHtjn4LOTCdzaqqcUxEa/zS5Unb1gGjYms1Es15FG
RcLnuMxC84NoqLvJrZEuCc4IffpyWj/37lE4cRQ4eXkoeAkEFsG7Mylxw1X5sBgxpS2bepOkoL6M
w7btns+cVl3xv9hwuoRZoPZCZBYvk2SuUGNw9f3eq87oF3k9qKDjsemxXydLBQsz9LrtVjo55YqA
eY1d4GJTzQ68c07EMkzSQlZB6wSPRQJL6aUamsupohVstMpNGzYtoxbuKPDfS/gq74BAMOUehHh5
ImeusW7uxn3llTrr2KwMlGdx4DAA/QkM+hbiauee5PjcbrUHMCD479jue6sEk3J9jKFGhy0lkP34
fhUechMFsOiDUecFS8y06DKsCsOTHMv1eDIhY2evKzXPm+5169NkcEv6s3SzJ1raUYnmyaWMOrJX
LcklCDi539cxRBHG3LzEIu9nIrbOnbARRwxz4louM5SNol9fN1h8tGtoUPla74+74wNLJqr+cz25
680rZTCF1GXBkGa2Mi5drZ3M4j6kXSqNjvgD5tCpFScb0yv16QCsi2GaOiXJhsUiba/IQXGEZwQ+
PkR+PLGlVDirfkBfw1Tm6BtzSJHkTOA1vEt9TB3rCsl0RJYcOXFnn7DSGsZXHS4qmiZeCVeIk48p
3k03BThkWsFr+qhWQVGhuo0MvlwN9g0+7bjXlwBciiPtm3RAhG3TTje7CNGvlkYBPWBQaZDfEL9q
LzLMvP5vcVD6R5L861oYHwGpxEiQx+NPk9IObZVPoFENgWl/9AKJgKAwUFnbuAXyHTvrqhKjbIko
AmBIfvGbQhtPqJwFZm9XLxjAPLGXKKSgz+aMXCHR0ltTOyiNpEIKnJxebKjjuKpAW0aIYuwLchuz
FcSaS5eoUebq7FZrWRmvB7EkHA/LCA9wgDAKoyDKRiwJjjyIreKIwuw3GY+EhnL+c5tyXAdVbuVN
bF1e6zIghxx6vuAysNh8mkuzAiqkZRp3hxNc3CtqpFlSIfeqCzsXGSlUji2Ap3oFhrjZkfHiyYz5
lOl0aGkW/kQxFhC9uuI0C22LQmOcSfFAAXaILmkE6JtSfjKRAUOI9ix4LioxNZI0UErABGyLyKLC
c9XrbUVZioLOTQyGHmtP2DBIqi+kkT/hGdgikBvXcA1rZOmz+MzW0Y9rxaHSHPkya402SVK5QJ09
YX/B1x7VT8lByHhOADphKN89HAsicDRYat3v9QztJTZ3hXoiAgnV7L4BJ5+YyUNZlW3SLaXQ6ne2
+G7ztZ32zffvX7OMfEygXjQHs7ivhwHyBeFhWK/BFyqZNy9Duc/W0kmbyhPMfHyjN93UN4t1cYLh
2m5JyN1Ph/zs6r4lWH1vHKfHvjySox337X7fCMEiv18P+3nw+31Z1fkHa5+6gFIrP55acvomO1aI
yzIQtkysmls6bvPMrqsqb3rsAxGXENd/0eOFAXiVUy71Y2sskLm8HO4oOWgrlRF52g32+pnkBfz+
9i+wbRmAH5ngqu3XJWyWgYeB7LLd1t45UIpkWH3W4+05K6S3lxuf0GB48iKlje13/YfW5MdqOH0z
Mt4vN+ON9tGhogq+G2dpW9kya+bKxp97qugGLdQEaYOFOU6H5XFkHD0QXtpUI/8B6BQBqclaRicI
1I8RLVx6Z68MErZQbCltnfa2X55nTwITVNk0EwTtS6e2Kfdn7Um9R5325yO5qZvY97kix6z7eNDa
PUidNhoVdEPHx2FtEkFU7rTyPtaYZcbme71V07zfE+G2SUztZ6L4cjmxV9XKa+Kcw49rlb7YTrWH
tBTbR2pTMQ4nB0q0hhAbyGx9el9PcQJ6zPR17f7Veam+Ic0gxzsE0CnMybiuf1b2iieJHyMRqs0G
NPEzBiq427knQVIp+go39Qn8kTa+WLHbRz39PKRpmJog2sThZfioBkok/ERMZvaIbN+Rv/rVDUW6
oKiK4L/Gz20O+pV2GQMZ224CNK2baCe+DD9Eg89PRlkUPyNtsbaEwC4eno07xlIUB30OAYpjtA9d
RViVeox5AdOv+jz89qGZGJjUfyN+8y4oendIEUPuW1jbasAA3yhzsLiN3fJXX03OrhLcHBxY32gG
pWAOnqZ1MYfErZlZm7XjYLBRh0wBPhqeOFR6wAgyVZUp65aRKbiQRfIj1t/MiH3oUGUlsyG02LCV
E511JtewuzT+M4bLk1reV1ju6zXhrC00OHx7gc3HpVgMPrR+H0J1KXXQAqmj/ESG83t/p28UlMLR
zX3cLdAPF5Z5pZarrjjXWAOjB8YypgLNAomXwVUWmqULfJomdkr/4Z2/e7pjkJgMQ3VRIvM1/75O
iClPpXXp3Dk2luaLnGWKHVckFA3I0gJrrW7+MX5HwPiNYkqcH/GF/5UmBOlFFEX3S/us3YKAxsq7
mswX8rE6TtTAE6QD7tZO33rmc4ofufkHcv8Wb1pTj5VwVzMlgyCValjA71G91chH+RtwndWvNy0M
7clEVIX8a6Z808W07h/faUV7fBEEFBr6QWOo+w1rvIcAV1gjz67x8b7GWlrMSw6UZBDqeQt2ljTj
hGNJ8qu5BNpMxZnB7Qo/q3zgZYsT403NWKA23aA1IGJYtpjTk/GI7/UZETaq8QJHK4pw+DWw53bj
gpdgDtqmdChw51ab89ABOslcVgCT6kbjOsvq0vlxarw+3mAL7eZENrTDm+uEqksjb04XkQHD28Vt
Bc2PKzg4ycj0mkowJ+Z3e4Yi/kEu3TG3qHQPGvqJGKjcP3hTDVuKH+wiWRQq7gfCZJ2jnVrmKp9T
gZMudolrwYu82hu44eZ5L9ICcDa1aPFXufXGFinH7+B32EOOR/qDiCQwo78DZYKuKGcWwXTybbyZ
Av+xWMuIz8vKbNH2riBPtYsXU58l4MN5UFXWNnrpTW/MSUWIXtJTMRA05HPXmv4JJ72wMYiQ6udy
zS5TLjfpi4LS87uIQ7K1FBY+0IMuzBOYTbFu3yOSK9k7GiPWLYhjOaM8GG3/jA+sO29iMy1rKpdH
MvZdaX79ZLPYZ14C01LtQt++pwFwvA1T6lUJv3a/I8luIoZWTaBCqRtkM0HxjGJcqNrLr+DjuxXp
c5HPd1a3Z+NPbi68ZR92WuMojqFGP34fJgq9V2YbSIrzkL0RPHahmtFZhANyuvREeYVvYStkfWsd
tzZhyaY17kqlKja5t9DSP3TroCPPc0McT7NRS87m70/YRZ/Xn+p+Dg21Xxs1M0kKstD13V+CjJuc
P2zAala19MMg0wx93ZRAPxzjKvOMASX61adOok29HPJEjWSerEcRQInpjZfjOX2OoTjYkzArY8ek
ub4VDlgF4izwrD/JTg2aV+IDbu50u0PViQtJ3p3CRhqg4ioW5HJLS9lvUXNuENm8y77HZOIyxAhg
vG9rUo1JXJl0rFI8VVIg7oLzD5cyLmxhiXBb68l+wJKHufcTi5MnzNr3jfxbUnk2dkqkuFQLvikS
y97T1pqRNxIue3CJ8XGN3M2U4PvPz1GNl9HyDnI1VNhlmSHM5xwQHLOVcTZO9O4RNwnYtONPVOkO
VvMJ9M0eMHvIDsIoGJgmPG3QFSPYuLHO7ah3wavauSqUlloSMkOtD43yzTphz8ElHNibHDR/tI0+
FrZyDADuc4RR9PrBPggz4mIH7ZaXQ4CCw8qBOxFg+qPnjknU9LihzmEw5HxMVmy/zhznXKoPk0bE
G53jHwN/k65BMQj1msTLSZpJv49MDUL6wprNtsBQxsTs15OlUYEihK6FA5McF96qk0rxg21O0Unq
cXef5iTFx6fxqZCKVYUA8vB2EDFOrp6cA3otUECvkg+fUXnHpgZlGg1f5DIswyNAHx6uswfhVSU6
BMeqHxLROGMsJH1IHoBVWq1Lm18ExFTzw7lNv+9nxdcw8Z4nC/pGVRCRIIvEsGLMUUsArR9auvnF
HHEo5XtOSxWFOEo5y6+GjIkItTur+RWj+G6VTlT2XfP8VwGY4XyAzhTEg5n4v9Mg2yof7MKDcIGS
QwRoUyPOqb5ubnE/m3aVMg9uuoxoqlUsQKubDlh+A6+rDpa4ihb46VOrcTOsajBRpk6GXoXU5zYx
NfRwtl/Qt6TacekCgOWQLkGTJc9+SHWjjFR6uDju5pQlUpN77vqhDrkIj3i0RIXsYmq1VBAWGWzQ
4l2ihEEoJKOBc0uSkEz8N41YNmfuzahsGhE9P4XRIwqNYByUtYqnTUgXuPZLsKCl/6TJNGFkspyB
blH6niSVqhD1NlG9Sv26JPhaJeuIiMO4ez7Rfc2XUOVI2ADzQb8W7jvi1s6XMaYErVQa7R1GlkrU
23NszqKlVZrDkwz2PGLASWC0fluOAYpdg0wzw2Hs0yAjq+0OtFTBo8uymiOwdPKUSq2hDlXCFbqJ
nElE8JC4kqqd8X6GYakN9dkbRKrh6y3+g1hcSuqEysdq418Jg1NvlARx5phwprQdo0cpxNwVJPfw
B0NfrcQZB3luFjGewhP8zNUFLlj78IixA6f+9pxw6Vcoj5olLN3nkVjCUYgQagWI/aooLeWY8EIl
wTyuygxwsBeuv8SPuOVwbFVhbP/Ke896kLSCEO4KT3XiNkfeCuW6yo2crmjAIXK2l5TWpeidqxh9
HjLEJUp0EcNBs2PlBdDPYmct8BVyvnasCd1a6nwc7VvmV6THOj+GAq624/HoLfxnXYfWgJlJdZ9U
NR45sZtnG7ZhWYs4YAwEooII+cNthaI/25RunXM1O58bsLKTtbxc2Ya8ydwK6vtlZkrMaG4gkVGk
TtuQyTb+KoJrcg2MXFD0pwvvF57YJPSR/tmJZYXgtYW558yWZn7gEeKkl7uZ2WfLWQDR7S+89JLu
gCe/tZZB6qkudR5wuFIGxH1mft44O0bbOP7pKAdFJgVwyKw29IJCHLA9KNbjS9ZqluXEFYkIHZWI
f2j696RDLMKqXQIxMEYv+e4/FllJ7Mq9gR4/rjEy3xfntQr97w6Tft5+5oOR3nB1jhpnu6f4/siI
6lcrVk9WX1jhly/5HNJ0Y7pojFImLxqgF93E+zIivnHZTLviAQv120Bp6ZlNfV74RIPXAsuNmjIF
Fr0uEA3h1ZlkmJZ2guyKb8yD+MIMjVjba3PZaImqpLAlu1heHqOIDxJ5nD9tmfTv9YcarPilYO2M
P5XslwaofbfF9wkAhNrPjPOKfsiVEfiY4tK496YvM5VdijD3pfFpHg0+P3t6Vpbeez1Iwnue2t5F
HW6iB3uoNAGlKUyy3XFRioBaRILOzOETnVYlyhR6KCelLOgxZbpk9giP5TK9kRCwLt8wPw9HGDQD
H5X+XYm5uIkVRDam2lLaHGx1nx+LrUSaV8JZoKd8+xAmRQem6kNF1//zRm0oLTH2Hrv5zKfH1nXY
oz75uVMq0+G2OjjOeNlogODXjEPInt7BDjCOxbvVpuNUEKI/83FEkZfszc8tMUUoZclbWonqPEYE
NhGMgIpKW7r1cV7+7chXUTNjBM/Uebn1DC+hJFbCVOsyHdzwMci9fnYrajavi2p25jiFbyGetuRp
S4mmcXpgovGzqeNNvszF4RRynQGR/BNIfRVs7dvdLCnUVnMlP4HPA2Vcdr9TXsCjQLQDQAxHxXO5
XwrBvW2/IXmva7z6TOp7K8CErLXmvqQzRkQEvmq6YfVddBZ+8k/ZyuJ4yDB6c/lahRXdgUJMzoEH
b+YkQdNaSDb+ERR21EGhahePidLw2rypg4mgPHs45ZsdUf9T51THOm+zzmljXkvb/gmfzruE+Htc
DlClquKKHbor/DaiqLwT1PB5DUEZwjSq+DLlBQT/DSqeqEMIKtH3Q/8akmALr+LGCpIaS2mDqbhy
a3Re3OWcFKOYLANRjI+QDik7+9UvQjrKv+nduTC8qa7HIPl0/EiiHA4hz4W1tYzcLWwY+4iFv1yL
7I6rtlnuNk2Iakkfh7rmJUfpXX9SPfP3d3ogw5WUujngVIDEexp0zZea1JPVtOW5It43WbMV14SS
4MexrfP1cNnCr+BT4jjZhOP088Vozej+Q7bVHOjtv30/ge3OWKJwG01n8/vkV7AL0njrooMsrnhg
TZITQiLUe5xrdXFax6k5P7StX4jPYi4Pm9UVFAACD0D3kckOi8c35CaQBhgvH5lxgchOI+JdEzus
f1X8UKrkD2zfB5IiMH+o4z9QUnXNKVeyUGYMHIfPzFwYypYpTayaXopOsuidfTVs+MOFeAHtlvqS
KtSBpa2h5tXrJC69t2U2Vl0OLkiTfrH+ju4d5JdZqk+xrcd702sSX24Ujt4PHZ7PRwUEGzwgbjBP
//A+ZKzmH2aIjtgFlDKfi9I6m6ohdvr0lCZg1yswXl6kOyk5CC+6izzgD6o0hngANmhzoq6qjxhv
CFT2HDb0ckTbhfyF5iwwiTrfQB1CQAeo26s8CrTEUHUQ19vU7bwWhGVk2PS0vc3eMi22G4JY5/t4
c77d4CieKBu9hGVO1IX3nQVa2tyx904b1AQvvZQgrBaqiGUURwC8HwNklnVLMXZo6thCIHlFuNCw
vMVpFE16x7UEXaRtzVWw79O6FK2Ul2KuRoGYVu4ro7ICXKN1THwYWJQ19Eq8K2tNdB+xwN0igTjL
G5cXP8SWzIR46rvVc/MeIX8kcLncxVBfp5sMx2JO3DtstAIVJq8i2bZdP4y6M03it7TL4NJpoQJK
5eRL3F+o4otNjaYNoazatLdr71tvVQ7DlhyTH6IPu3AD1FTuBLmEsrGWhsehdRnzaTHiRUxJ5QhG
yPMM1VmYD5stEOK8cxuUvWlDdQQc6CYl+xdD2toN1kgCxKVbepxguDzpLukdmsZQV1ypwfZquDAX
Qz6Q3XqO4Gg3Ko9XC4Y+DDpuvmAOPcKnvkQxMGFnRP3X8DX4uE4BpSoUDOqEG5U3k6ZPaxwAyOux
UUIlvXQqSHcaffDhdulu/cVG2HPQ3l0L8ZL30hLcZP/3SQGUXmWcwyCI4q6yt5CtQ4gVTYKvaFu2
cUxIqYPly3qsuHt2p0c5zgenkyvWTr/Yty9em1sdaiT+a23+lHzGOyUPOjosZ0KsJTi3KYWTXRgA
+6NuSmq0HRr653X9Dv4XYS2Z7wf4D8SuKcg3x8QWEuptfkQFwZztF+3z5rQQfqlVQSrKIXMhT9oH
VHMKT0AR46yynuPcYnXBgmePgQR9yPOstrkVZct8tGjPFCxp6nAPJAxLxFITt67F/L9xtm0SUbYp
WTcgP9b+Ku2+2YwdgauCqCfZ7kAqLDU1cjrq1jbIJhY39oHmN9zMI7RnFUKAyb2fgABoD6vMIqNO
02rY6wplHos4NScP91Af1aPYJTvIkWSg5RLh484GQ6xjvtHM/hwNPyi/Om6Adbn6+Cr4D0bxlSs2
tYGf4UtWoD6v3yOdLJCaiqXVueYx6NCBEqBclJR9cONk7Faob4GiOLYLRzIDT7uz60RIlQPjkOre
lG/1UKfZBEA6sOO24qy94oAIjD8H1rPvGzmf0O9NDE1+dFt9BKWZ+2a5iOof+LQVxN5BaavKH963
2QA5cqM0xzyYaZ1tc/5ObpaSK/uQOpzF4374hU96DSBqmW11N2YaDS5K5KmtH2kLbI60phN0GsPy
kZToPLEvkCn7SK7WULc7BugldVMUEMAvrCnaH6uqn737QyWOgvmW8VhAYSsM3ce1o3QuYWNXcX2R
h+gTlip3YJ37MhrB5DUuVKtvMipbqzMDV2/M3v5K8+PZxkiSEI3b4TTyoCjnCRmXNJQHuChQTqVs
08v6n1x7a6bJ3LRcBFrYGO2vSXomCDVbvWFEaaU+evLdmiTp3tOo8KGepcUMrILiZsmU9ymXdIGD
UcNAstLcnwkerSIeBacBhaUPrFOKqsGTnzp+z4N+nAYWftC+xsI54ZYkyMU7Kv26R7yqqlpWfYTf
evHmhBJBxGIb7H8vnrnLALpC1nz50YSmat3rj37815s5ij4e4iha+dObXJiaiVxHo+f9I2G4/KAs
1fY2r23WIWLKBgLmQik5qnm/VliLQXliz0K/bE5MkimsKJXcykay6araaRhCtXGYFNPF/gs4OQGO
dOhDbmGjwSbWF/NOlUExDu6JNCg5K4K9xvUOvMGooWv/tmidqxzBYtoRkSbRBW/EGJTLLqMnEq9c
WKVb3oAYIGeQ7JZndZfgLYUgGPj2S86dyZeA0YThwd5Gc4XMWCAeBlGCafAcUPUx60OxcouKntX/
EyLLk45onIrk7+Hji0QDwHqCmqVlmp5CWpLufFf9CtnoCV9HwbpfSGPafo+caN9Jd7DphjpvM34P
SUCeOSARUEvJmXMuZZIXiMYuJAMKsKOzWQ99V5jJ4Q9x6XDKM1BY+oRS1NvLOoB/pFTeCJ/Ng0Uv
U+gbfTpad79yY9mEjuJ2gEQnLSWCi3/HQn7MGu2bl6p7jS/gTetvzZ3mdgFXdhMQXY/oPrvuliQW
w/NAf15QtKYhm4o6I1n2incups42EulyG5M5Muw2wuQ/cRZ7+N9+RB56bIE6a6a/VdusSZ9npLBY
EVs2eYWhD863Xj2G+0SSNXZuBTQ8QEL/W16aI6vxlEgj6gusVM72eDa0u28tqt9t+MaE/wSGyTLK
QR9zfVULAZA/HrQ38BLQ5PPfktK9p1bawE1iEkF66JqIlrOx0Cj2vNYcL7K6A2g64HQREGgS/aRC
ugr1za/URaf3EHxLvEW3M/wfJMftM7z1pGASOfaa6VJTwYSSvTJimeUvHjPd6p6kgVoa4Wzjf6c0
uInPz+sNXGD3O/UcGmpTBmmd0WJagGzsg7VXsE6ETQfQKHB42qxQOlVgmL+37i/bPPpachRAkzJS
reAZ+a4fx9E/QxZWV2lqdoGNvKr8krZ5z22kuMAy66ZKMaXtPSJyyUucgrJbpFjUQyOyzekwSz0c
M4RmjqM7Esced7Yp3GcUgLR4HYEpLc/FGuRDYyyifkdS9sYmgIZDfxinDiRRjKcMZTzuqq1KnP5Q
sJlCWbGXUW23ILxqrwdZQ7fpypT/JN1VsuuUsl2uw8zRXLZn9HkBl7LIkO9mZ7qotehE+HOP1l8/
4rMJJ0itNInO3ngDRXzltqVc9MEwSS3leBvaX2mmJ9KItpiL7sr3izbJ4Nr/4vHURKY4RIP84pAf
4bDTqv5eMzte2AknIbYgahpT0woxcAOnFimkwzIWRgXooAxNpG6+kPoPqQLItFSKIueYvmJUQZjj
/3/S+bSJLme61BKBG1y/gJDFrdNXELhxGicl5HIMLZbWYVGalaN5RAeblrV7LZzoz0K5fcIyzAgX
n2GuppgdDlXxpZRuXBwFgitLpJL9C8dJFUa2SbRMMb+GEP1/85eGp8OtlreSJbjzAPV/QiMuN4Nh
7X87VEgvzx4gdaM8A9W1+vBt+4oAERDlVav2/220kelGhZ+GcmLutAxV0GFFDgAciy8bLfZWJY8H
DU3XGSGDOG47DdbfH4tJbqbNe2sxY3JULTdStmZ4OY8cpk06COlD2Tzu3rwXCQeOsBfybkpl37I3
HD7xvhy1Oc200ax8CInKf074uTp1C6uPWadzW2GaEdqEnn/1qdWM5m6pRMSvv5pPtNleEwp+EpKX
voX6Uze5LIOUtNazoBYucKEAdDmGfLKITJpS68CPbKNZ/+//VmhFZKv9Zl3QSfoS4O5cpPeovVCx
m7LahHULEbSXWSqIKwaMOqBfwKREfONW08WRfPjB+8ozxyRQ2gqNnV8pD6Lz2QIuFy/h41qdUnFN
Lt2GFSuZZOXqvP71O0QFjegURQitEDe61+q+8a1T82L/grIlRDqeAvbv1xWj2Op0Bv13BKYeykdO
8cWJJE4VDuCb5MK5O33cn/mjMlsveUE5reVAZGO8AKA/e8Gnt5UJWhHgiBQK7v/WVBbmKv988zfh
MZC/Hme8+zm9EQtLNlSOwY1DMn7nNQLISX6V0VBZEp84w0NuhSqrqaq4po3qAC1lqe+LWjEI/rxB
wwdIISqfs9sMpve82fYBlyOzazbRaKu3ouDav9soNznskistgyoQ6g2q/VU+rJR+TrHUxtyjaxfI
D0Zy8uzUH4dQn/ifsgR7SlENqHR8qRDfKs0mkUD+0hs7+wT9swyqHngksjowlw7VL5HfcEmTNrdO
AR3SD60792cSyMYeCnkdRmZQykVw4UXkA/UrvshwEtQAZ0M9m7kYtpIE8S/F3wYd80ade/EFC+8A
uS8zhL9Z+aLska+Tq92lZn5VjZSF3TpR+kbFBCmhhtolr6DEq6wl1SXA1yhykrCH3ImzBVV/lyrc
HuSoxFKe9/dGM8vO1r0Ctre8sehySppX6YBiz0kBPultrzcCxoqXP3w8HGSRcbPA22K/LLAH5zYb
p9iLdrH3GMz0wlN4HKcAEOapK55PQRMfYGiu/zg5yT+NzyAZe+8VBHOYnCsg0jr/EIWajAr9H2/0
rOiL3S4d44t3v7PTrcy2LBspevwphsnGgaeiK+mhhkQ8a09Dl/Kp8X6cHhsHSOVYqriIhzm2VQ8C
NUpRV7ll7dq1DiOAokHZJlnU8lGi49LlcWX+8lUR0+YH/NcrR2Ki7pCN7jkUSrfHedM+sbdkqmEv
MBst/1alzBm8wWgYbpgYHA0grh+eoSJVHi5zEaTcK0eTZdvwJ79JzS0yKseDk2x9/VUCdxILEzF6
DRbzX9ZQSM+jMfK2HX0dafytyvk55cQjz2qtoR1CLZV/iF3irmEvg0KH5YfMJX3NPq4EtccR7K03
5e9Q5vwEdzVOEEETbo5bZN54pNHu90YbaLUVbTCjbGvZSIjdHf83lw18zBgozKXyJfG/dXrLuliz
as+LWTlGnWaVLSfded4nRdRQ6RqT0RDsrMmfoFz/ObI6eUJg4aAt++kemh5WWknj1y+DhFZ5wrbo
hOAG8j+QE0QWwu5b+TV3Odzm1H6BQbQTXRjN/Ma2yEvIeJmIpM3drHNEfhHhDGiQcEmAETkWzUDJ
ZQK70ksOA/cyUAxzBJXRIU+bxK7Opl6jcnRVi4g7vmqVbh8FbCuTr2+i2wyo4ynN1Z2fQjcQkU24
naw9AzEYNPw3e2czRZUvh/OOp+3ABhl7e+6net9YA3FwjgcotXg+0rwoDCQAnmP4eAxzMFpJ6jph
gxMn0ntu1jYcUUJxNUSrtZuiJP38sJmLz7d4jHEx2fUIV3rMTYKAyMI7klbGyzjhR2aGinEl9+xY
XYdD6nF/fzdlnyz2BpiFC/WLwWUFuzNTcJPj+q6LSYTeH3lDzECSoIN0jbhRzlJft16Uxz/5MXpX
boDSTatmEFG5dVYgldPVirR+B9XLlPprljLNACze4pTM2DGxkxqRbrD3ncCcF1P8hvm++NYAP9fl
JpW21A6Hrhc1T9UirC3zx3pyWNisYmvKWcCwpDIbA/JvHNApa5H7LpUZWO//Y3Tg8Cyasg/auHYA
xpwMlrvzAXLtdTElfNDsxCnHZ0eQS7fTgVWJpYoEQl3FguMko4RJcl0X5k2yEizRcWtqysezUrI2
hEUncBVLmzt6/GQIPd/rhL9MS6xMqL9MkZml4MwbJMuL1YXuFXaTLdmV/NWyPgnhbXVYXWKXFgSF
VQyxz5Xk2WxA34onyV8LGRLApTfyGYRzeYyoj2iIm78tx9RNIxorlIOeeq623q/CzKbYoxgykKPm
6w5lsq5fTM1tJbZMZhr3rShZGEQsVcoI4kEZc3yRkIPocP8WJ1ODFqI/WMOfPgYgdLMndd/16IKf
bR4Snvovc5K83n2iGu08du1BhccUCs78vHwL1kC1h66qzjK6mkH2oHXFtR7ZushybPVoAn8g0STL
ElMKOChdLjxjbwS8zg2z1tsG22LsVCDPps3rdv6jx8nnEddIqHywtpYCPh/sZ2Sg3gqJgSmwmaCz
ZHXiLTn/JdcY0YAC5AxCJ0VNRw5Kto/pJ3G+C/zXNxTF8QM4J7Rcm3gm1L1xabhyzylanrvm97+4
RE0MJ/vdit9BebncDf9dAgClTRVxqzZRpxNEXGmU4/3C1OYMUyYJQjYgUHEGFTu4qGw0ar6PMgnt
tr6efRRt3jCiPreZevrKg42Ks/cp1LjnlYdbFmhHZoQRQlN3sqQaseFLzeanG2t1Jc0i5L8q9s16
uFh7o+FBIBG5ASPqKUdh+eWFbqBFFEMIlOn6O0ImpiX6G0iPdcN+4cTkoUUPhZlaqFnsvUcT69j0
t1gDzyEVBVwYE5CbKgX6yiWzpBmXrfvXRRrnL2j0uDTuMXJU5NgKNx8c8U9oCCmmzLSJU5qaRUlj
whhDN+uIgPXJaI6KgQ0MrUSoWp9509/lqFbhOYnBh6nUDN/JGiwqrrq6yvkHtwa+AU5LH6PBha+1
PQK7UKWF4Slf6GmogqGXrl++FOQbTv4n7SwcgCJhQUxhMUc9gNsMXjiS5xgAYL1YhwaHpvzhoF2i
WrL/rXLDgP3OiwHw3sMJC2T/DqcfT4Dmu12sVnZOtr/WFWW+m9R0+hV7zB8aM3kEaZpvjDl6i8Th
HyejG8q0cmwMqgywr0sap3k0VnKMMpCsx2QvYOdLvpezf4LvGY0oXKfE7lukQrPixkU0D+JPxVqT
b2hF9pcvnK0i9QHahnhhKA0iE/xzTy+ss/JeyypcoR5Kjh+M3bAYX5UYFSomktOch1KEei44ObPf
fe5MVSK64xEh9pbGLTE2ajd7Suxuj8Nc2oEBV+xWfzhW4g3E1RRject0OtQ4eNu/aucs+ZW9QUVI
2jjwRo3NAg89g5ZdS+Vp1l2kOZBZ1ppikHn06+SA3Cs8IhlYBxLB+laHN2zNU43vtqlnKaUCK77A
Daw6etlaw1neV5wKh9XrRup750XtKRaz4jHa8MwWOv4LEVIUIsHjYwJzH+omfcY+/gIyQMQjmQ42
KOwLIoWNon112OaW3cg/SWS6WwtzFvZrN3TP4pCLmAkEGbRfogYGaGFB3Obc7luQOu3ua/QsRJPm
W/YCzRmSh+6Z1erSzb3CZnHhp2WHaCpFkmU8KwrcuPtib1Mtk3U3I4Wn5XVSu/Mdq/4Cuz+VOMx+
7iPOFsP96xrnL+GaySIH/S6B8xwBO4NH4t0l7JohcFf2C1wlkSWZrntO/6bJMUZ4C/Pr1z+cTQTA
xJC1cYRdzEM52/4A+ImLrD7eGumsGJ2OeWlCip+sslbJY7Dm3xBZYCBK/cc6Dpf26QSieQ3akdqp
gqarkf24FIjTemycvOqhzHBvaXb9GOcm9cER0ZRSjz6pbCbxGq9kKVV5fQgRnUZACbxyPzcgHAGi
obZueE5lhlb/K03eepf/aE6Va6Jzj2tqbhdqDCxHYVcu9zy0d3SRAqlPeHXhOV6xJPyuaaA9R6FX
wj8LZg4+LeYxP9FsaX5CRQbPDL8/Lv8eFlGKU4B45bqcvEo09WnZpk5T08vzbppkd9WgUVaHRfxt
5i05DY2OzUAtODICgGEEfVssM8A35b8beWqvF3m87/eMPlz2XIe6lhtXlgaWTbamdyA1xGQovHSL
qaOsFfhRRz2OSh8qL8Y0xYeRpjNpLBI3FOsLcg0QjiRvW+LL1rIAlIIDVWJCWAx3QTPDfN9h6LuC
bVUvG2ME0Fc2hvQ4XAS7C0EqW7meDH76GcXMW9cTmLDKwOqGHFaDhxJ9cHgd/Y7koAC0xe7+F0fO
ohgezWxcdZp9Er1pLtwxsI7aDOBnojlqbETAzIhFWy0YOYHKpYOMqbvZ8GLBUZFzUQ/ltI+6lENJ
q7Da4cd6M6pDxhnrmzFrOz1LX7MtipsBgehDkDJhoQGXOR0I5YnvBe80iWIx9jdFUREnQ4ZuaOpw
FO1QW/z3zm1W4vpTNZGroMIl2xyvZOMvdSCJOEig/ZBj+Zrv1dwwiapkvFrfY7HW1HKtlpTYaiAS
24hFdooXf3XdQYU2Rgh8CAqKvemO6z8irdQOVJPA2RGFvx32PhDuFsUXWgsgyEIk1hpsTvaGbaxW
Ox3vNyD9Y1owFyS27sZWS87qT2VPZZ/CIwIiLgPpiixhgjxZRFPIARB7k/flxUpWfuiTXIC8cb7k
mgXfu2idbvyRqSx/tPbfjHCRsY9n5r9qDtUdKhruWf4gqMCayx+gB9R/ggsvc6+Dyj0XgKfCKt3o
N7chrtQRQoF8tO04tiDseW5Ai+u4l6+0Rd7SPrq5V4mK/Yon9p6jCx1tUjSwAwIiU87PL5IIvZOm
8V5DLOxWqXa3acXUb8Wr8s6Wmr3CViYwfIqZWng0Cr5GfLYWMS+YPU0g6wcbxOQkQuRz2F1MVgF2
3N4rDN7JTuofuF/LcugZ3t8boFm/3jQKRTRzufglNnH5aLpenPA0DX8OD+VwuUDCUUDDBju1RdG+
WUw8Wo+QuaiirBjgVfTpICCzBZy7E6Al/4Juo0DX5cgqN0/4HCFtt2i1G3R1bloS1dYKabFN7irk
rmCWwjd2e5dQ9Xr2AwGA+GeXKwdmG0iBiTnSypDAZwiNb/me1sPm8mZDlVFcG6DDUF0zG9Zq9gUE
rBO7op8yKZS4pCitBkW68nkAwttTatd4DkMBZJNcxMb4Tx9pY7jIzyleg1FzKkZ839W0dpK4v3A3
1U7rhm2JHVXInGcuuGBzugcMPm7dOnFy7/7EPf9MeiNr361Bj1DK+oRB3K0S4x8Jg0Un9QzytOO5
pcUQvOISjk2pHupane5YIY+jTdVL0+2kh5ODDVSAScCKRREXDOWRUybAw6y0izjUKnyCmUktbkNE
CrvS/NUPIRuIFyASbfr+VNowCBiOYcfarbiDORejJqGqQW6+Pwr+6d5m9zu8xgmMtBwpKTmtCV0T
iPAl+tjfg8Ecld7ef19EiBy2X3WniBbF7H6yC0I4zX4XXO0jmCA04i2n9Dpjkoxx+xF+APKIrjEJ
+ESuumTZw3JxvTmJOR+RTc3/eRmNvzquNfpeO+9N9ZxhZVIfjPBtrmzX4OQ2rKpHkyZmNP4ylKYB
obttLt2U0gb17VVFnTvPZj0OrPgZbSCQt2Y+5wbtC4YDHfVZRIg9ZujFtEz7HhZ+lxUODfxwjNUB
NzQbM6K565fPw2xVyXzpPbS7WcQJ59ZHHQUNuqG7sWCaJqY3N2IbpWpBxnesqycY6oa19+CQxT+H
LrhLdEiAauOt6xSaOBWhfuYZrVAi4U3KQfHYFiD581UuGZawzSLbdbCuYs4yDAIYKiElt8t9Xxjm
4aXh787/SJGyJUkk5UO8aAQ8/6rS0+UfvcXxlcPIWZ4C4XGqcRcG7kYzyy8zuMkwDvbn05vg9Zw4
sK5q/EY8+boHCGFlrQ7eVRkitJ+AFDdp8LxBxvz9i3DfRTTialn0ng8BxkXBU7auHHRv41JYeD53
3bwR3vRwjrB/+hQOX8b4Dvi8oYmU6xsQchb+Rj9SO7unQ6P6n6PXZ5saoequzGULKBuCrWZ5dgbX
EE1IILGeFhh6wCf7nkcQfCubvEIcw0KPGQHNVaU2XqcGlSjppTCAfrHNTYRR6wYP+oVeJCunEQqb
nHdIA9YGtBo3MHxA70d7Qydum7+lk+wca/9jKcfIaDsh4Z9nfzTvjLtBViIonx6cmA5Ka3roJkiC
EW2AHHZ6Hoy/EQRj2FDZ08GyRsPwLSJHICtOzcUzznZOtvcz3gLMf5hlHD39ohCaO39w/Omi54TI
4xc7ZRzWPRShiPWxt9yPlnmRe4cwVqBfhYrlHS+IcZJrW1hXz7eCVKjK0wSasaf2NGlpI/fOa84t
b0aPUbiUr04Y3G5Xyj5GB/GHw7R4lf/M2rYnJXBAKWKZ6sXM4eLrsRR+x44/upObiaINV/tOqN7v
81SOmMPddlQWmc22bS3l8nbENka5NIWLfzJWEbBP4xPhOQwUHpSBGdAMWL63F5kBGsir1nGSAh19
hzaPsXGMOfRYhllj+EUIP6KCtrTqndlsAYPcFpkEwS0A15NZBzbWYtvkkhddsaRau9qKZSGzVd5p
G+m/gdSuHnKyaIOTJFJgUJ/v/ZVEQ0YWgAAudVZvhxn8Bj8pVa8SbAW6U6monBhHrd0ALeDbiDO6
1+jQZASkSthpSYYJvk4gg3roBFOOFGTYpUR5luCkHOALGdB8hKCIg9j9g5ipXN46KLCZTXz4U64R
XRsjobLVvmp62rlymFRCzyZxwB+JUCJLJFAriIWLAg9wQrO1YLLyoaN1pM9yLosz/Sar0q6YiNn5
GgH3HCXEwvMzZBmZQ1/apZheQPSPF1bNdn1WNTVG3ixQoQxHgG4XvPY02tPi3dtzMgYP6fWMl2Im
BpXiNNYJ2R5+nzUv9lExieaIilZD98/gpWRKRFzsglvGJQaXuf29p+aNix19Y458OQHXI5V23LuH
kfy+n1Y6HqulPaYBp+OU9aTLmLknDtbpFvPrK6YmlEzU04bQTx+iNJ5UFDQVXzf1CUPiP5CN5YGM
JjVmezQAmY/ytmoTjYUBamWqgWGnNjKGzj80s4hKNnN3RVZzao6N6qYPn/7zvWaDlwsax7/c6sy1
HwEaD8Wa9G0VeiArcMh2JjyO9Bm5OLr5KnKL430lNdosG3Ug+lyJWTvV4ivXXJ2XkiPvWQUWB4rf
9t9k8oVbPCimaqFab62rnKth+vdM5F0t1ifa7Te7vtPq4Kseux0FRNap4KMGLf2sCjy2S/MQLRKA
0+JAs3umrJlnDVxuOA13xXbSKeRQFWnI3TZPl/BT9MJ9BFrHyVsUUYrYBg509WCYgRHhRlY7V/Wy
6059x6TYXzR6UgiGYIRsehfOFC7radBnopB4xw1zvaPtC47SWHpnTrTLGqwNMiUS7aychCMeFyZ0
EHpzaYoQ0xNYkqIrNgVNOxHjC+sLg8eiNwEA6oSYr3+RQKXHzN0w7WUV1DX6jNLMlDMI3/p0Cefr
77q7/9+12LrG1/b0uZX0dpvXuyrz3UcIKfB5qBX5Dtak5fHb+z3u3pI6JRwc3xYfNIv+CYySXBKX
AZG52pv+pphFY034V9IlJNLe8xCIDb+swsx6EmDCMi+P0mn+ngre7WyHR8hXX1eOPvglZ73FaAy+
XTRP4YgpZ1jZD5areeATWMWIk0ZmjmbLc1Wmzb2tQxMWj7EwmB7Cmz4jeYR7nGbO1CLgs4PniRAt
1EoC+V9YqHBB6m5ljeYzs6ACjGRLo+VnDDwpY7sDAcMXauOKizbg19uVK1u8XlshXD/4iMcNavZT
O0yIkAl3WVRNkpX0s+d+Rn949jUxI7IahNJovcYCu/d3VfLO2ElM14zbu3WOpPayKrqp+bhivvDW
w/4Vv+dvST2m+oKzL3U4tarBnuJe1avKb9pJClwkMRDkP0dApusPgdu7FHE7RnCJo7M/XYM9r4on
TTlfBWyyxutZnrmrPW1gqM+Jtvwh5fqihlbiSZKgEjqKE4WDeo/y5XyzXBdCQiHWbrQK+ON0rX+7
BwS3bw/jFdBdt7NJAlpkZf5FLB2WMt7UPaTvkI0M2bb174LqMMiJh28i6PE+bBnQt6jxIalT5NkY
0bgclPPENriNqbAe5MaZBgqM4/FmR+pa4qni0oe89346X9NFmKq4hTmeoCjrx1wpI9pYLLEZYIKS
AdqwKwJMGME8rg4GcoGckx07gdno1DhtkusLFgaUcWH/YKhSgeqzeyqFcZ9MCNsMAozA5u0Xoefy
qkAm0ZCdHtwJapobe961JL1Y+yq/t0owiILKEf5FwicMhn5gAObwnERToTs/LlSK0CdPExqC20CF
ncdGKpQCJcVYBWnFpKLb8xdbjf+tARgg7DlVqSBHKPAPDgpad3QYX9odenMGI8IjLMoGv+/2mZco
GsvOnQAFWEorCMK4WpBk01G1SdkyQK7tzXSVHvNo68KO8rj+1b9p39lVO/piKyN8Gf6U5xhpX9l4
RAhzPqP1h673kXhjGCuV2b7ks+kTePjpZ6TgjG46QmKm0S1Xt0KQ62ZIJAHPpHQu6r/e8iHXzEEb
74CLWkZEGR9eTdh6qNfIUfQceTn878TfVynY1v5br1fy3V3Df/r2xQlYraq8wTWtZRRpDmFE99MS
6K4oIV6TXRVNDh1R21dHKqM5HS0gf6a4/t1bNZYRiU1kLHQ/LvBvfABN3kTEhaabLcDWcSDzKKw/
xHtPR1zqWP5gQKLdhesHuNTBZq5iH5mNP4JyoeE0j0wgjKqJP91uoN+2N2HFL/IhNCr5mYh/ZzcX
IU2f4vdJ00+uynJJYBeMuxtsYZMzuIrgaysMDiS8LtdFpF5jlc+YACWjcenRV17vZSNDOE31peMC
GYKNCdyyFFmuI0OKIiof3H8t/fdmQsBFxMkzUPPx/dLUvfKKUhsDdRu4ZHMzH/V44jCxEgGYTNvu
rSNSZDjVyC6V6onThmJDO1Bt1oeRDyn72J/k06sIwHlyK9xqCX+LWMkG7xrERAa4g1yOmzBisRwr
AIkL5buTwnq14yS2Fw1M1Kx6Wyyie0CLEcwFSsiYgx3BsTg0rWGhSv2sZnpJBPuB5wri7wAE6Wky
djeCfpx6dYwvC8J+tIhVvScCKafrQ9DERvcWRJBLgxsxacvwvOtQlmNdLZxtP8KzCRnxsqCKTO3U
eZZX0jsWzS7aVu/pzO8L/2U218drHiGBSe1o5rQa7FQR3QY1ZF5KrPs+mNuGCmOMefYmcG2YRbJI
Z3Xp2xW8N60peon44tMKUezfvPAQ8YQ70qYOntah7mi7pVsuu0LB8EKLdmY/s6EH26riCTThU6z9
pPrwGXDT/qQ3N9TGNYYmJ1+BZTXb706pp1feoL3yuoYlIRoA+U3Eil2z1aBYfFEBqFrP7fAvSfk7
OBhvlPcO1mjnNpZOSWq17J0mzXzEiZicMhOadNR7svsYZlNNo/SF89sH+xoL4qnI6CupEVWRAQA0
EnE8cHUJwnfXorSE5m2apn/sngfS7HzOk/wsPMfWBqpcO/y1iusmovznUAf4TPtpGaEH+LTZi5Of
DvyFJhFD1G+zAnjkphXPzeiLB1Vm3Eq3fKES/ItFFnUje3/k1DCIbtwPuuS0GFaFFj7Tqe/Y8XP0
MJx12LgY11CuU3jT3wKiApJKa7SxSMJD9DomATxFJMO1Y75sDzrpEoeISR0ljtE9K78wCP+EIRLc
bLMApm4Pe7zetWC1ArMafIeNHTNnzFKJRRV4wKCK3DOe6RHdqfjjK+E19YuH0cngbF+qiJ5IFn2g
3LLtE8y8D4W41SzNH8edBGeogCDB+0lY+nPpggQvlZMJ+B+da4b3aDHhnPiqapkjBxk+hU0wotqs
ZQW0w3+07uQJtj1a9q+3iSB5hauf5igeZ1mUAO0s2Cs63iGOHYVScZ+Dz85kksSSMMJJfi8p+hdB
u20+L1S/Z/WU1D1SW0CJL3SB+J2H0zAaMFpM+75HyHdc3sGQcFGB7qnNQOp934S6W8V0LM5ZCJ8I
vKjLOEH3b+6EGP+eWbRIaHNUefd8o5j6655v5l6oexicvWMy1ZFvRl0nLMp5gTUfkYPqKyOIpLpU
nT2TzJNQi1v9yKZ5S4n1KfAFVQ5OnSKX34gcyjPzv8xpzf39yytZX61qKnlijeoWwM4OBF+zxUAF
tuCi1qu0PaJyQ/tFr6GXIXnxCu5EQgU9mojv+fX0BUsrQJp1FKVz62zDOMLNEpAN6oWbuJMkZ5/n
DNty531jEdfT9NTOdMUIZ64DqH2iTIWo4b89gWcOLplfswKuhuW0AlAkTyxu6HkUzJ5y6g4gi3oe
2YidIonAp+BF8MsRs7Wrg+MTqy83C+64shqKN1/n34Xe56a7uhYn4GuDy6c3GowWfvGH0dRP2iL0
0Pbx93hrPkcrhCs1Yli1HtQky8SgmyxnRKiDBcjWkwmxqCOBd1CwHE4SgHqimA9T3VJqjbaZKbok
9sbgP2/kRL+ONz690IQRr1JxwjAD82Y2AXkymSjFLApbxK2b6D+utMnsyKL8ue4ggmZ7MN/UFRC7
T7WS6s9tXXkNtfF1fzXnHSSOmVf9L7bKxK+vkMbD5oipR3YoPGBJ2tF0moUPXmkFMxc2YilM8rLU
O2OlrDqHWqcuV3f+CV3kRGrtxjv/NIG84CC7/aMaxgyxmJJgXOD/kmaAtBJ/lQkIfS8RGyJ3k7wE
iEcHXjYuYi3tGbVflBiiz6rdaOgAHKkhHEP2umC7xW18opA+1Hfw2nIKhaXh+FoBKSRe2igkVhdd
kGpmCikfqgKWr7Xm2tp45qUH/szCi1PUdKF8OxIPPQEq4FnmkA66u+ZVTmanBrWBNBMhLXJ8PVsp
dV/UzamQBIPC9L2b2iGlskK1XVGfvslQAT05p29YQy50rxDAKEmoLhpsXUaA/RIRXIOZNHkQasXX
6wztQcYvdW+/bq77f5otsFmNkQYFq0PK9BuJfkxEkdG1Jz1iisbR9fcW+ngNjrwGyY7TIwXELBZY
sIHdvGVOh22Qc/U7qUoQ152aERM4QxVlt/esTeQpIJ6qXvy6ZhkwZ48ChDl7Oc+8lZCbUPohTYtu
AsSM0p6/G23MSKpHc2v3EPZSsKnEkJXT1EgWP2ZtD5aZgJ6BzfPenvm31y+3CtOb7z7aOV7TOpQX
Wdekv4CEcjMGhgUavkHlYxFuMtTYPR0wlhi4dadZNJbvnX7JC53PU6CGItlhcjuaE/9ZpbOFKA3Z
7mHtYEcypNbuKa9gqL/uIBtvrN/NHcJi74GowU+X56pAoPcwtj+6FsG0lKIxd4HF7Go4ghe4dxH/
1hPd8GsIHQ9sqSKBzIL5Tw3ze7hhfvTD2pN7SiHpmPsrjKLM8YgSRD89hgrB1xcD7kAJq4dYSM/B
asZSsLvOaQXAE5iep//AbM1KFk7d9GZrvMScBKDiE9Jia/ymouLgR3hsKXYX7VJPh+VxFwnL2kqf
dBG7+b9SJcO9wHZWRLg1ef0eTNRWMqOECqqpqx1QvtDrkUA4Xmlfi5SkSeiplFOdITTSxxqFop0T
ZhcynCizrnnmzCU30Z5xCTPE3NMaow0VVmMwY1o/ht11IsAdnO6Sao5RXFEoiyfNGaDYJW4v9N3o
EKiOz3ualpg02ispUsfn6m+n2rknxYLd9fvsQk5Uqauj2IBB89TVtuxqB4VkL5Tu05jvAyrfI+DZ
aHBBqiLo+wa0Naa/ZVaZQVBo1A29IMMapa+dUZhtqVQi/TlubtXXs4XPYvHAyFhNwe4lV55Xih+J
M1A7resZGW8M9vTbCQWszwfc7A8D3KXTv3z7U5ON2kGLHK1xJoZN9M3HfSTSYgjY7/+OZmgtTqTb
3CrrVcB5ZhoV5ANP3poVwPXFXGbLyiEtZtWwq2katCSiMEj4+dx0FJxDp0wgX0tFNlbskMVspohK
e1sBkUczna9bBHeKVF7b2rvqG6WCKkoBfyzZXd4YrS7ew9i8T56olciE0pZOY6xb8AL0/xhyv2an
ooGiyCI7lHjK540TzsEq671vEUgnY5rB2yzrOnj9hRUcRZxF8mgmEMW2S92MoJMYPQzaX9X+q5Ct
D3u3kLpQ4cyOR25FZAynudTg8fxS1DcV7V8ilcROfALUO2lyk6wqUbnBDUYOA860+kEl0Olezcfs
NBGUryl4gg/Ik/iGEVnojcyqucUu7Tt1O5YsxUXP4Pbuwx+r9Q8z1dJdRsBmRpix3EDM2UZdLftH
56DZvjgcsTPKazRsf86F4nuju/2hBjPt90fV7CbBkJJNtPW219sZv6/7hoifcZ1d/uUqtT2+qrz2
0ptQQFCII+mQ2lLlMAi/ZhfUF4pOTXh9cbA8KD3zfkGhyI3NXkIeQuT+xTw7OV4nCPuKwph4M9qo
Wx5N73k6emSQ5pzi6Z6+cp0W4GQcqQhAX8Knv5XqsSvkboXj/XJ4ZrGb6yFjTAhzNnVymYPr5VuP
k6vl1GmSWgZok/htKyFIyNvqVi95yzM9wqURRAmJxQzNygULb9vZfa4qUPOkPowkHuKDdIgK0VI/
KLOAx4q9A+3PS1f6x4N5acDIh4MvE20DPoe87fTPK29nz0Es2wYuKnPS2hfqXr6LNRnjzbxcCLOo
AdtYwwi3fvdYibEXL3F6YAbapwxKXepwhK7JQsQXd0G3xUC3nN9+lv0lGqupHsirmd8aamyXK7S2
pBDvjbl2gwnT7yG2FqXuxbPn0uVABy1HGT7G7IxI6NuTacWKUthUwWa1apgquCsR/6552PvMnken
9gqGv8Cj9z3ESQ1qKWP0joaGsMsH2jcYxq+dxt1lYS16mAxQU9FFnVj3lhxEWKIc1n6ux8ZdHukx
A02APTmrxCG05D+d+lx7rC14fWNqmt+4uoZ0lcnuqPgKXCm/SdV5HOHbC0edlnYGTd0wzmYD9OAa
CE/e8tVk3tiP+NUU17G3jR/ujYV9n8cgElIuvsbqM0oYcHy/J7IHBlsuWXsoVrn0aUhty8oTxHgh
kOHzpuCizb17IJKWLxbsudPqox63RhF0G5OusfNw7HclPd1YXNlNbhpEwwQaD+2xi6uPvttehdoq
OSdJwQPmkwb8Z5BeJjm/DTvBCoUYeZLtObxLnHwfBLMLXcmfmvb4UYErMnieClafH+TmTP6trQYk
0/ZEiE1M0S/kgr1iXiP9AonBDHGsYjFCOzxkBrUY2z/2dKgSW18vvPgWPwvkBQnJMGbp7UFzF2//
hKwrSuA633HuIn7BmrCoBdaFm/8zsBJ88X3R4adNeJXaFle6zxZRNjD/FSxalnZfn0CovKBGwMJc
N9nEkWak1XlIWxHct6S7cjBEwgsyNpDZlJUu1mXmMppbUCC622BMdPEEzOa2YscBr0/YNdUKDTXa
CYBN7ccpzyGqcRYA2AXLGuNa96s3wxpLrBo4OSrNZh6t9rLIK9SiM7hSaTAFPXBHg/fDtwCrv9nU
J76G+FUiWgRPGK6FcCX5kLRZuTBpndGij/0MzHLJqZTkvNp/vFI+xMUpvE9cqktcLk+A0Fyszlcl
GVS5fdWyxmithUYk1PDwM8OHrADnZWqjswUHiawpkOJkHVS0GlFQ3j/tv7o2rQZCDw9ySEc1KjMG
ORD7hnBZX0VGpwHaxd7IMlKkciUJVXFRfW0h/6ceMDKjezEvraBujFOrd2yLds+m2W8usNfuz+0B
1elgqwiFXApsyF/xjIV4PUTlwt6nzxP82mcoqnoB0di1R6C8J67uC3+Te8WGkrKz4V3QQDH3AaxB
gkRgoIyl+6+o+81tw5LOSUAyX2vOHch5qnBzMNWmDVU0FwkRQSjXD4ByCLPIvBbhQqXmTEIN7aoL
K/nbFpZxBLvM88+3XUY1qLKwVpv0FkbgVdQSUSJnkg0iWfWjdC4fPjwmWjWvxC0jLnKuxIwzE2Gb
7sUqw47/nNcZqknkpbTdD1HzvkIALabY7coxA9u+wnWb3OFk/Urm3525bZ5dbV79z3ixwqOB8+qE
laM8f2G+dWbnMA+3EwfNc0AkGyg26fyMo1a+P4dCY/wSETVKYPK3tyf70POjhnjfDA5AbQVv/oEy
nqLW6arQQUV1KETE1Jn4GLE9rZsWByGLXIaiBsV1mJO45M17v5s7WfdJRJnVVuIX/Wlob222b228
MWD9DTufgRsLtrJFKNEOPDrol4mLYXOLIMQs9fP+yvrMadl1aFccjyIJIsru7MOVVcuq1wTmhT1U
QjYYCDl3MbZsbLXB5sOUvJdD/4ItGx3zC6FViDaayIKJ6A93BPpiwVNN89SJCoR5V16lsQ9GdGNG
kMMozU/UR3VWmGKGP60YygYo0h9J+x1u/ieyH+CuL88LWyhwYdatAbfqLHHJTydpaUAfTR9mSAuE
hYDI/dzh/Gf3mNrGXCCijkR4OEXYvB6C/v6/6C8OcUO2kdQ77z45hOFlG9iCDYno6ozAqWxXxuL5
RCVS5rdyFcyDkfi1Y1makvmr9jqylPFwjTIYVajhLKuWTZZqu1HwplKTdkf3/rTv8ZZEUoNcWoHt
PskKMzmBmHpfLMoGaddF3sfL44hhPUrYZ1Bd1ZCnRnnLXSkvffwUJ/nKTrpLi6P38r8CgL4rDx78
UJPHNq+WrhHJakbve4clGYGnQMPXPnLzDL2VsZ8MXrEUwz/TqdSpjSTda/vDzWAjh8gZNZL3FMTq
7t6jpzuWPnyuAW9AaOYW3AdSP49iprzfSTbKpA675JJYgNlG3QaoxDzwjK0chRtMP6ImIH1g2FjS
kaaay4t7LlCmodLmj7q+RDFReUkU18iSn/es+k5O4tWvsLNmlrygu9HW6w6fUOKVwb1uBz/AfNRo
5L8o+M7DMig5zNLvTJx5+kT2Iaam23PGTzrZWDowx9VKFKfuMgjXW4tPw/zGuRXmVF/Mg/K95px6
TiFUO/5pqnBgXi4pBU298ZZx11963WoL4x1/YQBFziLK8NhvWRsv29WHDgJU+CYKli2bgaccBFye
HwHwz76zszuOJFrgyxb8DsywH4wJDQm5obZr4tEpsKNBIZrEWR05PZ3bqZ+W1/78ZHu3N0raJFNy
PxN9ICo5Zti9zIQVXNcwy+Oy2EUMIwQ0HXHjUef6tVgpuLXTUmnDzCY5ctfKGqdee6X3F7hl5VM1
cyJ9khAOOfvz2VpO2UvZUz4efOEsJIsFP+x6MVRtFV/432oRAbtwfaXPBO//RAaaSmxFr84CCjbp
Xes+sEtpJmASihsVjn/x4Ct+o5GoiihSjMiAK/w3PEW3pCOF++6k+rUACV78SOddsYsTz/NUJzzR
mSyXi5pD0KkUJ4IFaQ/Y0mCe/ZFEYNBY5jh0a2Ez3RsDPYuN0RPBqp4BdvXUJmilkErJLMuIR9C/
tpJ0p/Rl7gOB5MFp8OBr/TkguMMf/4IQWQIx9MbAYSUIfV8MQp1yXe6H4pMA7E8ePrbNqUIDUE55
BknRY9Og1sI8DVQqfKl9cw0Qbw9lPcTj03T29FKyMWZn9pAfAdJxtGNPVbNo6XCTHJ1jQRClNZ/V
vu2OvXwABZg0BzNdCbELkIU+D6sl5aI4+BJkpkjoP/ABM5h7Qn55teR1wy9VWVdgdO5zG5Ggv/5q
91di1udKrry2HDuRWCYVWv+h9gwlN2CoAQr+abFVT/EN3SlPpzyk4oD6w9sYI270ltDzUrhRb3qX
Mj4YOt403M2CCdLUjJT4p8dJc5nhTXd0EhfxkkgMiYrWAzLEX8N3N1coL8D7diIESp/6wscU5eVY
uspQ0EkbTG8K5qdIf+U5v9Z0aXpwwhfjgCsGVEtj1q7/taNioE6sKEWyh0UIi21B1Npr9B09pCBf
cqVaOEX3YH+oYhaYamP9kJRAdDHUDNMR3PuLPk+w72aME4kE7nA783CTPJB5C7tUMIL2JaAyFv1V
CBwI54QyBdhx7DDjk/mFCNp+XbfpJXY6pPwsnTGaOdOfQ8GhYfcqyx4AdSDvW+2qBe86Stdq+WUS
PTq7XwiNDEetj+9dwsCYjoWtjkEdqcPg2si4wQnIApoelL6xTisYM0wx/B+0Wxink1f+XgN+DsYv
pIt2FEWkZiTC2CQ7xaSVjsAq15JnoW1TG1JGuMeq1AGCWSIVBj+Bvp4xsWEcTMoP+VUqH2efkjrj
U9r6NZSoD2H+SmoHeZB2BS+BmwqenDrdyVzCX1LAFUUNV4mtE5buVUM7kljIeL+5fzljVso7BhrH
AR/S/QCEb35KczrY4iZVuWx/xvSgfqaOVwT3kse2+9VObtWNBLdfTSKkikBwmVY/wG/VvNiUP57w
fghHB3Kkets3wOFVa2ma1TD4583u+SKZwbo9/VUJNJVZAFI/mLslbLus9ur1Yo62O2GxR2Mr13hw
AnDyZgVUEAvKNLfw1tGyg09bbSR7Q0jYmqJWSK14gwwHfRRPTu2uapmzEyLI7tdv+Fg+0SgrYdLf
gWTsH4O1VLJW+9YGCd/ZDUef3ipzf1VcUW7dN+DFI5av2ynlSFbj0piTRqBEhFPcfXn50Pnnj3cJ
THRw+ah4wmk4w+8tVh7VtdQmKSR1wP0rL8TurpfDye6Xro2d/5ZoKDWD+EKswpMyPL58f01PCpA9
J/THmno0netBHEnzHinFRrP6BVLuIMWhX4d7cQGapTIZKlMwM2rxSOffAQfZ3oCom24h+Btllqr4
9m+lm7BIWNVvrIdPjw6kB2K34fzunKZ1RFw792WJF4duK78rXc/xEmG9UTw1F8nlaZAtRqL5eFS/
5eApe8ADzOmhE7kkYq13KOx8SCC95NL5/5GP8K3mMwZm2izh8tnB1KgE/8MlNjMMrBDcxUtb2d58
MuBsCfBjkAQ2VpRxm1CFezegoJQZBC+ZrbVl1zfKnugeC1sZBg6O8o42h6KMR8ur4eKhyHbUfjrK
UMhnKPPkLIaxKvcfV+dR7p14xfNwsXopkFnHUpEz1JeXyLwzIMcixxWYAXCccHHX/EVEpOB54UH7
V4fMsLeyfmDF8b5O8/zwmdu5zZzb5NoTy5LAfS/0YJMC+up+M7u/ZjhZHI5ktApm+Ua+DNd4n/Vx
ea9FhBM6pvz23F1AlRPx6pimRRdFRvFBZVuoHc8haD3p8ZV6is7aHQ29zr/tf2ZQcaPEjMo0S6/k
cy3jdYCrSvxm0p/blHBvglSVwE7Jc1rFaCNnM+LRhPRsz6WRvQ/cscvqJ3JUqxUmWbZsZl5cbpO+
I7GeLiYq059UEy3HSO0908zp/qYTKHAM3a1wvEA6FqmI8f0DfWuC7TDLSHkgvbdmgC8azOK707Fs
vYBgnKGu2nVeUdECIqGTnkMoV+90sYHTrULY67CjrJcx7f8rzK7hkTHop2xLH50z8vuZTnyXqbdz
2+vZaapdJV/zn+PwQfREXVCittKESe4ROjsMDamgHa19rI5PKb2k0ivjQW0+E0JuSuOQhI1uV9hW
WaVtqJ+g/+q6IVeWU2jNV/dzMLzuqQZIss9Mmhf8d3qkn00JDDRIo3pzxDZQG22MBTlDUyji1bBn
/2EaDBEWou8QypIZZwnJAoaiHmN29OORMmZnLJipZ2HiItUhF0AYY5/YHA1s6WMIwwdscPhosbIV
c2+hXG8cSBs5LHMQXuLLGHPouzb+uqQGPcJ4u3hIHM9wiLAaviTLYda9YEcaCBoTNH1UhJAtQaDv
7/gqOnWsl4kS3ybZUTp4s2SWny3GFk64xc+IqRUH9yZgBMSXqkKh6X+VXy5cLjSgF2yCJW00yJ99
KewdNqkqdwVJ+p3xTQmxMwYgrS80vv1ebz3ck3ljtj89gaElLX7Ue4MT71QlqsJUTWJ59MndTKfR
GHuUDgqF4QEBuahzJB0Av/LcZsjhRMseNZ5r2S0/0SYc+x3qjRHMeHN4qtztTvZF3c3uJjhjWu8O
RCEXEvFUn/qbjpu/tjvUW3aYhgz6xwOpNyTyCCdRBNyWlIUakNJkkmr15OhGBBkHz/zFITt5zes7
48kZgzrxr5VJC0eNFCbIR75j44MrVDqi8h8L05UpBpC0xbb2vKBD+XlMseivc86tbp67N/iy9eiO
Vy741v/DDlxV2WiA67gXTTjghDZL5qnEJaMHifDz27vbnPr0RQxPjpI09jgv4gaotUUBjRNzX4r8
3Vk4i5lMYuksK/ijwsG0ledwTSPjjbjgj9mPHxI9EryjnLS2qtZbIPRWUkFlUBEdr1ixweFdjumx
drODi+q5jd9xRDPSHHo1AceabtiMJU5Fur5hrZEP1S29mX79ecDOKXtLMGlasR22pFrDdqmyPLMu
e0rMfSiquS5l1LxCZCsJBfU7Y8jo3yYSXNV0l9rLcO0/50oZWgk910J/rnww22s/JdRWd2oXpRqj
ZdQK+jgl2tnq/zpsF3OcCLrHSwcAVCYa8nM/sbc89qiEpQqxy9w+DZ9wzRyDJnzsMoEoA/XGqrhU
PHbXhT2yPJ0+9DgL7K0rXlHDbAZ9B/zxLZe7DPxed/nYyZQbyjKKvtPdty/FVIwudSjN1Mjs0bvY
y0CIrwtTv0Hj+klrz2muX1I8YFFQR/eQaUMKu4O/Bb2gDXp15O3ToZQpYybge5N0YjNzXlbWZbKj
ZSsGpGOghB8vHDih6R7LJmiBQn0x9R5cL35JbEw2StNLwjEkqYHdmWvuTnqQUIO1xFxgRX87hAn0
USDNalZ7b68om4Zi8SDsbo0fzgvabYeIduzfz64jsbckZAJ/HzPCtsEQM3qsUpq4rYTXXQZinrAR
mdfNhUcBfdgcrqsd+N0et10y9CW+8MpZBPJE4Zx6EhGiqfg96oJ/3Pkd08FHmL6h1ulyO8HivOV/
rMByHbL5qOS3murbKi8x1sUpnSKG0GpwG52Whm+ycZCiHSnjSxNwGt6r/Oc90o3Uf4oiUYtPn/Su
THLoMoMg71BOu5+XdS2Qs+FyKwJor1M+dEkAxOrUuMxkKxXAMViNs1MrNW9zLEZ3lEDC88Rv+gWk
kMRgrhconN+5GrRFh5DpLkdkCcgNdn/3Uti3swHVkJzzQ9woQeSgj0q9oSVP5evj4wH7aYk5MvTQ
ErT9ZTYd0oaxPAkY3BX86fi/cWFTx9jvp9PKWPQcE0g/4JO6CGUxzl4IoR3umQo1ONPChG2j02IC
CRr04ZnaCVmoNE8lgWUM3eIWrzszE/3TW5M/6Vj73tzIYd5jDLtrneoM3WoSJFkulIiqMKQisjjU
IWwH90KR1N12bXY91+Xok9JO35RsLij6FdhR0BY/0isrjBx48fMGA35V1aHNRCWWxQw+q6mxOK1C
O8YpaPr+fOv57dgX9evXUinJXN7WuISxnPa0Tnm1ZV4Qo+wVY8hTkosH7Q1NcwQcTRPKyD+wTsn1
uOCm2/Ly6sOr0x9JV92Gg6liz4gMHLj2tyX9V5AkYTpx1O18orCwd2/r2bX+nZR4eJHdOUsV403e
fytrkMDa3WsMMajMXZ/Y631AmDwPWTRyHdN68jPoJLfsR4OYDs3g/dSExTaXC/PxTbXImz/X0hMc
fYiSDeCFnGpsupmemcLRZyjuSDMGligc7o0jPNvlUDuGPNXpYKruQHiKsrFSM9vGkR9aGi8mm/vK
Mcga9FWxficVJ9eQtINN2Ow4uLB6vphezw3YO/O+yp65viikqpaEoydQ7O9nfEr7dJNLCpY3mHxv
Syi1E+RxC7eqprbGtNs6FgYq0OiiV1kkQUKrtfUl6QvtcaNA7Gt9g1PfhqeHXpY6aQcfTCbthpBX
4KxAwVUYV7gXA2IFxRU2HN4QkN4p9TBn1eZ5QlSBywLj4dy9Z6WG+w2GrQN07Xg+myhpZRaGq5bG
1BDRObC6YGMosX+2IRYaFVQmS/WUTOCbdwnR1eCZQff08Y4olUIuia3Lr2rY3kCJcqdrS6GKtGfu
R8g39znM4A1JJ8nOh5SijzWk9RRTqEuFeB4a2XiQOoDMUkuBIuuB4xFLKbDRxTTAeD4hVebJMF+x
aai4hQdaZpt1Hx+5LAQuqqF6HBnM+H1bzt6kZ6nWsohU6+gOgtHzmL4BgYb+3xL3h3xmouU+It6W
WpavsnXwOlfLmLFKpBeWhutD5bcTVms7P0yfMWe1EK5klw5ipPccoqZ+BQ15Ja1UEG3SPHoMj2Ke
XX8D01ClfHh8jRAPVKGi67jt337BujvZHoWyKCKF9qP5vgg5PmqWx6LcaKsX6uYCtd47IlIdqc/U
nw9QzAn0/GVrHglyCCEBTfFekr+kjNk8hA9pMTcgBLxW7Qb1eXDDHTnecSn+9synGH9NnvnkyBkt
8KhcwJZJ8OgFmsBevjT4aMNNUMfqml2asxPYfUiP4rZnzhMqnglt49gcwh2TjaQzOTme3cv9ctIt
RNT5dOcdItLOx4R8C5sZoiffaq11KO1oCCC/wUHLB86QnTNiiHvS4clskHQqN1QfWfib7q+DAOtX
mx/GZ6metPWL0TvsqZ2f3KhU/RLFGfdlo/ur8uEFMWl9ijMMHyoYcunGlg4P/u2oMiek2JmRbYMD
cps7G3jBMmXgpHOPalIv5AMD0+eb1IDEgzmq1pmcnRxaezWAhYQf7nHNvb6czsDaz9A/9jBPTgMf
VzZRaLfRXVjc+pijY+/TXUkRZmdOhviZHkhhSIatxprjIzYSEadbY0pJZZ+VYhYMX3FRzMO50Xv7
JFlGJ+mDpLwYJEY7QhqYJIJCFmBlkt6EdwHhhUX75yShq/aXD92PR7ekvPRK5uUBx2Mwe5cX8D5Q
P6PgSXTf2Y6WBVvMLohbuXiL/FIB3RfgdWxV2k5s06mHW0w25i9VxK6VsaaZPy0vc5GgC1CwNQhq
QkMB2MNdXb3tzTh+7Oht9zCHwva7IIrgj9fmFUImytYqS4YiiXggDxPL/m5sq93gDAvI1W18Q8hr
/5rp8fIUredtGQSGv9fdN5ipWzgGXNkdK1UGWecOKnTY3T0tUEiJjRrUlT7oHJW67Pxt1ZMwE6b6
vZGelArMdKTMDimRhyL4/k68JwMHQBcXv6SdaH7Gybs/h6OBHU0AudyC1tp2He9r+TaNsd8IQA0j
TPcsRcxXSOwFQPp2XyMMO8GzLHbGiVMoHfOpsEOTmTHWR2OaOUEsIoXnh6I5NLE5PGJmcl6Hcww7
lvNo+Hw4qaFbFzerpDiLIyLqp2J9qVv8SqSO1WuxiR0AW9ne8fbArT9BEKzzG5Swu1X16qNzPXpX
gyGGopufQUzp2BGaOowD2/KJHpVJtI0zP3bUnVma9Qd/+HmuSXyqisVJL+KryJlxpxGB1VRimsZw
IxZB6BP3Aimgetr78WkHaSbBo7YpdEkx1pcHQqxAxBjOzLwz7BfVenEcUdngXZTuDmnHijd4E3Fd
ay07FQsdOkSbG/minU0PHMkVy5p78K3n2P5fEsqXtsaAJDqOYlOF1yhFIDNwapgF/TGxTHUr0EBr
A0mxuAYgCFWpj/zHs9MT7zuZbNamv8X9+wGof4ycUU/uIwCq95FC6Zbo3GtlaSfUmtNSSW4cBbVX
RS7eVzZT01915RjemDa2HucrYv37PtWo67YR02+JFMovh6A6QBaeFkSMsjlS6pYbsANIhWHxozK8
gzGv2iEvZqEsCzXFv/tUvdYGEfrjoZfNuDUuYYX21eI/WN15XNYo85op9HOPR4Ce23hIYN73UlIW
CmiQ4iaeV5e0GuZuBqdviNsKS2Vic8SorPVzR2nCS7fnDfUeEwwklLbqoe+734Kn7s99PwMHLvsk
VnkuZmuRb4rfMS3p8ZEAu8M1vw/mWThYgMNeeS8j45y8uZTemUIwJTkSIk4noWgDkQx5pIW28UgS
vCFTXP2cKTY7lMVR2XKMXus/ziiASUTz5dLsBNeR9cYAeUppwSQ+niD8eoQ3MA+0pd6FJxahWUd5
NLLEISgsA1sA+EzyCS/WbISGyNQMwHXZ7NYzEg8dZX2RimBdNu3fDU+tGzsl60Tsrgt3vwuGAZbK
LT1XgAZ5G2PaUusiLx4AA1aie7m8FgG8Yc9+XhUdepin5cSd5aeFw6+1kaBw+Lp5mBAZKJ8thmm7
sXLfnrEeyHrNkdckwpaaY0LKxUdwfIAM2TRIMImwcDgxXPFOQKzdPivFl6S5r9X3QP4Yx0O0F+pd
ZJu0UDfIlql8K32i3Kl4i7TX1IRrVCIGN1aStzsyt8jKlw52EmRnOV5+EaZjcWeGnTKCYU8kLOoS
JdOwgh7RNRb/EEJZ1Cgu5i2lOxvdzIP4svJ8tP3pxU0fM9eBuH7+anFFGn9PrnLYzBA969O4u6Go
84m59Crm7TWs9vLnIaka+PTvOr7qdw16bprDHbXVKAZi9tsMyxOXqzGBN53Z8yl/ayk6wQopmJrF
4aVClYojWDjqSeKtFlZFkv7IW0m6BPJVI4fSlyHQLi7EfB5zTU3MnvQHPbwejALDsExDqW78/+Aq
6x16jb6du33mYM50a0wXoc21E+2BbMRopuVhG0cgapdL3KiZuDZnIN7LchXx18YtrBfHJnoaaFV4
9gyq5vHPTwLpeFetxIbsnrrgPG8P5P38A+maYgrFWs+BYPUrq0X7eQNrhygi8J+e+FBiy6RlwTpV
aJLPGj1BnsmPykq48IZ5LxDE4VruPKyey0kbz+mn1IwwV/Z0xOqS25cBOA1WChzm/CHkZaBisqSd
mluUf9O1zrbBJXQGkp/ufQQe72OZYVkesI6AsAr4hJMcuqQ5WU+TtqtDYxEZVcDbjJ+Efpf+Tgpc
3S7DXAM5F26+iWKF/PbaXWRxtGlh8OqUvIA0V6j7dvSYgKTC6uMIg+bAqUNNJc5k5GPw9QHVt4IF
wO/VhpulMr4KVCdi1IgoCkTxOdNz9aLZpAAcvLg9cLju2onNj0A9bsTP0gXgA7D7PbRlyUbdzerB
jbPdwzSEAMWlPHUE6NknOV6o4mcfreSBYBws37e1kWFu6bckKKmdILC1Eu3DeuSf/DREy+BVQC45
RYe1u9jh711GGBOQgwoH9wQoISMGjbq9VrB8fbyE358ONcggO5mQMngM/a4s3KiitidzIrliGJWe
KW93dxrJ9xQjH8zmNJ/PS6tGIRkC1tnN5j4+wjEHkRMzoEgCcsNx595IZvlvtSFyNTzvNqRHzcz0
G4wm+cjPAAtatR7DqTY6VYwQK8k3ZrsZqIC03XMTpW2HOhYbN/f8o3CN0mWPknjeDWSsFgB32Z68
X5IBWXdwjhntctclDKgKuasyUlpuQYubXPDwkytM9MDROrmavo/DOZYertOV2rRNYxHzhazzuVyC
5PNEGt9RIdhKoOLo8soOetRdu35jEuD5Aj3rjYkoZxuWxFjt4qyZdpzS5HfXg3ibx2lwGDnaR4HO
ffVwG1m22H798tJqOSqejd458lWcEy4dVPEt22tUo5RUO/PE0kIaq3mPy3WobQJ0DopJAezI8fxd
BdFrhUHTqFRXyP6X2uICuNIqdWDR+SCFd360/VInO+yjbecbH6BBv5oX3B7DYBJ3XnYmHpzPfqxf
3RxFFg82hkNRHO72GsLAW6WVaXRAG3J2Dbiy8BHWky1wXpUKddZ0x88nL/2LPDuuFDM9PsMBCknh
83uPNuBdpAxsPhsu7DNOSE/WwSYNRA6VPiPETzDnNpnhVLNxHZRZuG2asfoozyhM3bTPPTVmGO2G
OXp9a/9sN2PIEkmpOMGDu9VGLutYHdhBH/a8i27aJYZvHNbRagUgp0wLYV6PyIUJ7i0oDGLSsixH
IpP641hOxmWBusXjjn5Ov26zk+N8R+l68xOU+8WY3X0Iup5k3274FjSFLyZ/SWOljGHPZCgQJhbs
h0EUDcl3sBk5qLzlyJzMLSf44FZZpkG/WzNDF6GJRRaPUEaIzZI6garl7TCGd5EDRzSACzaMUzls
PQ21ILoRCPoXAPyaerw6a/emBBXAaLlWTnfWSarBmk7zWF8qdl+KwAJnXEhpLYsZVuVL7QGoiwIm
470P+aF6AN6+IBwVFHR6MFq3syDi1Tebf24sMallosq4M8Gq45AIq7x6HLxrx+O8+4J570r+e2pm
AUoOYoX2NlqTH+yGxz/qrcBWtocjMb6F4Wo1uSjYdstt1joA1WYUXrB/F0KHJfWUaMWUGPKhkN+6
053+YilRHxye337LVY71kwumT8SzK2/8rOXnf1bj2vIy2cHdPsMZWz4mfqiueweoJ1c71JiSpnYW
Qax7nkg2zJ11ZoRcML0i8kOCtD63U3Tt/9oqqFyfnmosSp0/bBbrbQel1Lg8VeSycNGK7NlSLlQ+
trRgfuYk9MtPcMUnmR+zHBGqVr615Jx19MaSv0b/JAlq3UgDlC9Slpaxu9hvyRJU2QpF/bfdN2Y8
MJYzT4qdlvTMcLhnGsst1E9e7A+oNSOp1k+IBV8RMQQO3JIKjNLiniG2VDWWQGcMa0gFtN8XPIcC
ohnfVHKqZJ2axbKUTl50Id1daFQ7IFuVwpsjOuLTcDQEs4UsopAlSuDJTYGJhyU/R9V9tQqXsYqu
E65wlTVh7P9GE+mwUDKpV34z9ExJ7W8zdafs7wj/fT4nNm8P/PCnIJD6he87tlhIx447y6c4y1pi
EqTDksTVEowKzzeelB7EW8xIMUkdxJBVq2cD0hSComrf2mmgh5TVnoRAf1PemeN4LjNHD6d6Grho
xN2frVpIhLTYJrhSMPciDDMcOMve4uFUWzFrtvg379C4XgLPpNtXKI7OsAlSUHdwXEN0jM/qdkSJ
sXV3r+KPZ5CVsKEwtojhRcie3mueZPfF15KH1TK8oITtIdHngLf9KINyUVoZek6WZ72rSzRYy+8Z
a9rRrmcmesugREEgN0HYM7CpKSSwXO9qIUJZ9RDh2jRLFQ/m8LC8M6iLElL4b1En0K61C30uDCm8
LJKBc4A85yjkVuVe7f2VISCzVeVpvqHoEVu4XmJwoegcWlPr7kadET+Bxk4VMsTYGT4QNhfD/crP
RT2ZRLDzcQd3yVhU5NE7Wx1zQTu1dxvhSIY1Dl+o7rIIiDnatCySFL/U4gS0w80fsKR8/B1Yb6Xn
04XkG3mXmGnH5kMyKvVILtZoNAdbJ97TQmeuR7EwnLxKq/M1QfuomCZ8EDo1aHjwdEODZgBC/yur
HSQxauzKWj0Yi4qNeFauYjML44+3IZBgsgtYm7v90WKQ7cuUJ5b9DrM/KJ44YoDPBUuOLV8PB4j0
06WwXnydFesFRcPTcF9oUet5Fb1akDzweiobXSrfVS3NZzwIyWCrCP2TKPHYp1NGefC+MUWMF4Tg
PCZzmnY0+CTEPSwCZMVyQUud67Pae/Qj6xG/RVV5JPWfq64GjDO8Ti+tDxYBo+Zoe+eWdEMstFoQ
OqOe8lrM/NKJ3K+WkginGDnfLpTgCOp+EYqYIcJsT2iT50j/2ol16QgQ+KKZ3TBhR06JeeOIL1pJ
QIHBXCSAXgm6a7VVU1CKm1vTuuYpyo/lKKPSVeCwEwKBkHlQThNIxxDFwnFepSW3iRLO68G5Iy92
hkJhXd8eqjnC5xHA3EarNYeffae3Ia4L/SKZFjbWvETaxjTJCRvFyXBULrEQ75xWKJhB9aXiwTIa
GyWAVVYBCRGZOs+fBb9J0kvn8R6AD0DpfvOhHaA+5/CBBzS997Z8RDPaO/EqcN5iUBF5Mb3u5yRz
19La1ZZFHDZuRXYB57SGp6mbysJet3G4V8xVEjaoMoOAKtuIdJB8cBG2uptZKTNqbVsDnXRkhmc2
R0wgIuP+xIXa7FSWDRI4jKM5V5esi3EmKo9f/0Huq/LUCcCpJB+oH4vBo9/+26BmS2iX4ddAnLZ+
ESfpvkva0FtqiyKJLiI86zedYcWvNB6l/lfBsuX4OC1oOYiYuBgsQve6GNnPASpmj7NXfoC0WIXl
TdjNYyd39jGZ+UC2VFHUeurps9EcvScuFkAaeh7ubWWaV+Hqen5SyTbK4UO62pXV/Oc2yD2QdeW0
XvwCNEs+jidvqtxa8Pkag3kosbfYRMe5ESbTbVsWGVPnvXl1Fm0YDRXZOLHHQdSAxRCRibTTaKSt
i3iJ5ZFMiuLRoTusYZngCjKbEVbf2k97KQ4LhYZFL2nRGFzm74A051wvIn9vJOHfOpMXl5DRI7A5
O4xCUAYUCo3dCX7EGZ+tTEj+Xef+NtvQpk6Qow7Rm1kTGQoS7hVjaENc7W1aOmNPOwh7xlap1v3i
BQsQxWPRyU2UfVFr0gbFe9yVpVEkDjG5WbGUBizk+EY2yGX+VMmzbMJ9srsX5MXKuiZ8DFm7fGR2
pH5ZHL24neTcvN2FYqXMaVAHFs+r2+BVbaGDJmGGyHstOpFcC/hmPQE6KnSfR72pXEg1axIZNC82
oG42BrRlacBjSlfSrywdo4XCEKY70Dmbv3xwu/tZZyngfRI8Q//Ag95veY5AV05FgLWMXH9VyA8T
LIBCEFoSfzeOqh51vT5+7Cwzur6TF+3rNhokbJDaejNurp6Ef+7nS3hdf2+JYcR26aqjeedqLrfO
bRZHTrCU38yj/lCzT1EZkBS2GgjMfjUDoFNdtmkFOeI688U5pY1jgcBjtdOvVDA5FDqHiIxZ+Vz4
EV9S8rNlWvIHDXXzjISxAUhWj9F/Um0kngXx/WJXrVKAgiBUZMNSbz5l2HM9+5C6FDvjI+2WNIcm
hZvgAs2Nf5cU9ZXM+Rg73hQccTnRUAhMgZ8kxBz8DHu3bU0GNi9Wws2I9GvLr6lS9pnpvg1V6vdX
ZIpCFvO1OhkB8Lc6ZORyGjoMTDcDmR4VVvJ+PegsaoNV10/1MJXvTnbdN2dGR7c08D3ToTrfUmWf
noJYXWv1HOicC/0z2aXDDMo1OFVbu38FEqdAhcSGg3tPsqBoXHjxI83zb9gTG5VhHVQDg/nSYim1
iQnOXZLRgrMfpr5zzOv0UB4ZQnkPCNwluyqJW1ezhQoOlmPUY9u4okcEHvJbFhZ2iHuQNMaIqQX/
9izE9NCGwYBaia39/TZNJexHXHwO3nfXCGaq88KzACZCrO8nn6F5F4ASe+aJjoVgaHkgkiiFAZJS
vBpbJ5f/gwJS60d7qJO5hcCQAXg53dsBSmOhNF0pcznM+pBHv7tDKZjilIZn/7ssZ22ODMfB4RmV
gJUubTs/prPOEsTALfVUh64m9LaS6ByFHO6WahignOs2bxC6gTSs3o3yDnEFOrKhJvH9XLpswmIZ
AuKDBoofNGHcm+8nCvW4RFIFyD3u4HObEKru8ZwNHa+5W6RJAYGDRQuKAJ9df73YaFVWpPFOQwvq
pWn7L4aV6WluG47fgYk9IE9gCfE50MNSaGYlQNU87SEJIzze/Kmqr3dqjk5C4JLZYwBTQJ/qHl5J
wEkSUgoxWMRNDbVHZ/gAIN0a45C/xvm0cWbqxu8/K40URHBtLfEPbJCgApddbPcrI3aPuPWTFBb6
pGWY8ajMwRNliE1jrVCsUGWQ+sv6+QN6lhi/hfLmLlqLFI9/dAqx7abzF+v0lmeMQkEs4I5A3ep4
VYfOwvne4LxziUBtpMr8adIx/3TKgCSJ/MSrA7Q/2/HwMoabUCPZO5yyeP3JjSuLgMsLT8okDcT5
S5uH619LrcKLld9NEU8mttx3AoGhA7OVC4t//gO3ERfQuPtb2VoK7Pax/QhA1pnvvtaIIEe0pSIm
FmP5fQznViOlYq27bniy6e5ytoMNCcsOZnGRSciGA8Lm85zmudznW/o4j53xzljn7Gq8cUt6OE7c
ViZkoJW/cWGp4s+FxlasK/Z9BTUFswzjbroULItMHgaq8W2VhHEjnoqAYfOFgm9oQIk5lf4tOmE2
uejuOaC9JT+pyFcCD+T7kx68cTD7fGSYh9dB3s/THIzghfDdfXUk0LkzlC/g0sRKV7FWOs9L1byC
IN4dVKknxbDVFnVxed6TwaQ9p6oNClL4xubej11MXn1T6htYXpjATj3tRpgkKDeKECLlct0g1jDA
TDTTAJiuGxc6YZ516wcpv0U+L+ssKD9+w8xVrHL3P3KbNgOu0b6ibc8gj/V74YgN6gY05XwhsA+f
nGmDFiCb7YaCoq8kAU5BLSpY8c6AOf8Gq2mJ51z3N01f2yFLts74TqdA/Tl7HS1hoPoY4GoGtPqi
x9OSjEKFv/O0RG2GaIyef9PZkuiDpUX3UgyrIhBc517uQm0txTJOaSIzJXHGjDKuVuAr6LP1X+M3
7q/z1J2X/jXi6wbgswmTHdTkowlCXoZxRzgACVM7KaNkc73+zGmF47efoIL71a3kcQvtuOckvC+q
PkSeGtRSN6A0Vj/HSWfKP4n4OKb1jajeQZw5IALk1LW/EeBKezsRpxKceMriWTkDCfvGCB5hZ2El
a4rri7F35vKAu/a1cxiNELsebEpxsnnORQySkMi1tsH6mLuY1ek5bocWHeX8IOgFvlUX9vevcVND
gSaSLfEx6xPRKmEcxvC38Duz2LYpWH1OM4FBHs2lHA+hR6ZS2ogOosaaX4RWDNENbbJruZydO/eD
GFMLuN3ewCNhlmvPRG3oSusxBdLMdCi+FIuWWJqVt+urImSL7zmFJDKWRqyYJZK/qrRG27b+esJ7
6Cqx+uYGRPSSQHf8nd4b+6vweAm5/VaII8p5KEqgzzAENlE8Pq4VPyhmZ/RqrpBHcjRCLNG502xM
GgvNplJp8CAZYQCYxCqWLW7tb6g1Kd4+lugNl7uBPp5McIXJMYOvArD8KXVYZvYAhbsLm+vOlygu
PSzJJkwqJqSwST/KixFpUpdCx+/XioYyaHcBeomzM9FrDiobl3hX//S9uB4Giv3tzrho9BEphTP7
XcueI/0bRgtkdEHUxeP7mG+Xcgxy9D93Vpo7+Y9SZIQRal6ZjX9Eei9ra7X6yBXW5qH0h5d5yFyy
yHHlnomfTq9ulDAf7INVwfATMrE9gbRJLahkNWmukcIIdt27GstNcUPSEDLO4TeqEdQFbRuZu/lG
sDUN4HUUbrGKscirHAmIJTcZ+6sAgf3s4ei3YgIhZbEXF4RAYLQf69LwzsHPijfpDAOtkCwMQ/fV
58NwD/jMeMhbZn2pi3Wx1udYoBnhZa+GFzDKYjbffq4ZGBGU8lAEp910PsDzuQ4R+AyoL5CY4d3I
mENwyzk0rcP2VhwW9iMCaRpEkeWoBPwFpakVpIY0C5SGrIOWSN3X5+gai73tq/yyzzB2Nxl0aUZy
WEBWqxJABF58c3hINY5HqMutrRwChMwVB2BzT3I3TKlXZQcEvyREZwA9tmg5/eE/U/PDxHM6q6sq
2omHx++0FQiPpWW2wH8Ze24JqFh8ij6GPKUgZdFzVAvPk6csYpqmkDn6lhPpWbR0AKM7qB4gP2rO
V0cD1PnRh8DOwmAdPV3pph9k/nBCupRAmWRONoATw136RkSIEnoVieTx/Xy/k5IXHqnlkbdyH7wd
hTcedQSRc2NwIV+IIZZPfQbbkL7dNGs+Lp/IJ6Toc0hf0TxPghcpfpJ3UbMfOsQdwsgJVYAyDc1v
Hmdu9YeQD3XS1C+VXD3WZGfDdp6FwBkEltkFlxPALztGdf4x2h7pG0pkNpvikrZ3mRSp3V+yuqWk
IaM9KTjmgZnXZQtiCZD7uTuH2xAaKhSeYlrII1u9qQ709rgwvWw2aQS1tQdyIUrMhfb5BeX5EbIm
CXd9OuWKfbccSUxt3pz0tFr/dLKh/FrCdNDGfaFsDxQJyt0iOcFgZuFdIa5vb7LK/sIy8F3GzkOy
RPPiJFnI2Eq6JG3kPk9qwMLvU8duZu200zJpUkSV5ai2W2j1mCEfJ2t3syuP2wM1RzTqVT668HpI
dsXI9tDwkecM2/6O96oPvjPDBlGGyq2BkuCh3trm3FIqqg2QUkM2/hIUPt+lGRMYIExUtp1fgBB+
WCWCwfcRZRmUuJ+B/AHmDsXW52yRzFJMa0f2tVzwf1ZXJgt5LIOXh8oen2Lhg6dqwnd1pNhBln+M
3662yWGSMj/uKwaeBoYsNKQDcOQXpXPO+vJ3FvRDZwTbPcSd5mpIvTSKBYAOMj50F5OJf1dcCTGj
f9PPDcVYm76oQQQ/7X2A71PuZRGOyNJv/pYdJbsA0acxlR3UfwZSqCZkGtX/iKhhaUDS3t96pTES
KjxjgEF8JBdAf5U90SVaV8yyQsdpUli2P5/ov5rBCIKW+xb/rOylIcCL4X9JbpIGYjIDCvDGu3xb
ghMHegfRGhpXzJ4Acb3VTGY+k/C/4IpnQnVg/IgUxPxxPYPrAE2yhFxWEHubL5n1au5ITdJ6nBHW
g//YZ2l8lnqwV3i3SIRkSMrLzqRexWARydPnS8c6mScDpxK5vBawgXevE7PUhiLXpf2WLiDJ4umL
4oKMjL3vZvWOxeBi5ew7o6XqFwK9gEQH4i+PpO9ZnCp2HB9PwWRS15xqEsrYfl9zYikMAZ9HKDKr
CeaHNilly24TA8TzJzKxjKsA+LVx06dJreERODW2YS2Anl90CUooWRKt6g85LsLgJn1WaJVcpFOm
yV5AE4H4fTTTX1jyfcG0EvsZOR37KjqFNwYJGnxtSh33xHN4rn3PoS2qoXKA6vFLwbWAK3CncvP6
bETRMNvQ7qO4H4g8EE+qgIKkh6tmGr9b72WOCS4b9VL0mIRcknmSzb18DMJW5cRtq63Q02867VQS
Re7byIwkcXblMoVaVerYHMriVZiJWzhfsmbT3359fIYnmxsMlJOHBz0ODNqPuWXRl4QGZJ3kO7FN
Bk/qCPFc9Zovw9VrqJIe7O3tdnhBW81S8HBg2rxEXQ7nrZkFxHwspwODO7dzwUvHWxVPZBaJ6Hl7
YhV3DKD942oU2dPwcGPJt5UxVKlGDmf7oBS5yPBHMPDM6jQNkVmLSfj0VzSZqKvUjSx/2RjJ5Da8
Ex0zJqPUPYjSyLsHwUm94gIO7FVARxbKeniSBFZ+fEV+mpK9oH0Sr0jx+soI7L4Jfy7MbzJlNFx8
QPABawapa1+h3EVR3AWp63NaE9Zqr8aSbFToK140R6ppPZmwTnaQWqD3WtC2+m5MZwe6WC9VrRzM
g60FxHQDEcxuShyPqLamSK+499+c9xaZxgidyR6BZ4vtQPe2xB/IUqQAcyR0WoMadAjAfOavT3Lp
od873mCr2Vsko75III+ZNoxxQ8hrRCTkaKVYte4/jXEIW8v0Ao7391rJSMJ7SFKiBDyZSneWJWee
9l4E/P43bE+KSMMUi/d0MlfZGU/ZcVxaVbdMsu9QF4TbFqDAS1OxHsPHRBkQP8hcCmXk4LwZoGTw
LnBZ0aWAQh7qx5fBlWBjlK/mZZ0WTV+iPrTqF+0yEes/KvRg/YpaAn0CLTuFOItJ+jWOvGUBo7Ml
x8nH96xrpSZITQK9KILYzcnvh0gCW6SHvp8Q7V9/PREBrmuF9fQ1TEFNQ/IyvijeHQJFDqgyaQT5
Ba1VpmxaMI+F0KmqmnWNXnxj9GB0mMDRizgG2X8Sl69W8YYUQSGwEscmFiYQDjcn7RDkcpoytRzz
tBNXcffCXHZiwtnYOBnL7vtuvln16v6y1Tedq3hLsZEjihXdTHNQ4dyvD3m1Cjh0oCBe/3Y3qE8D
N+TfE8wdxounOMUlsb7pJmEkcELd8KPaL3M8MvMf9lXguz8D6gvHqAGMdMZH8V0OqdOnlfL73Fbb
enRkeZkRt18I6XL+4DYcfP6/kmUmJ3G7mJWhOS5qh4I4WNyetMgPH8WoNsGRFf/8OfRTP39B933e
+CnMcxhopX5b4MyuDRURD5jf3QdNscYjLT2qCmdXKOzRDfnyNjJMCRM+mXHocdTXhmvrasd5rplN
jYDnfiGPJWvucHqxsFAynd0D6ygMbDobewYgDzdtYrAX3mPssWCRYH0vUnmkUETE/qeMYMKX+uxd
Jt+ry7qao5aD+yPACIsrz0V9ckhHlJhIYNA2+195q9K4MFZ1Xv1fb0WjkRg/YR1wRVKFAcd+Q8wG
zzvwWOkHOvsbEmYFkNjNPR3yiP20WAVF5/wYUNmqsfju6ztr7Vlwhco3W747/t35rFMDTp24vlGv
aTMF9uo6nqzDu4vVsMIME+bwEwRlhxuspAgtuUKkebxqLmqUlL6yfSMcZqx12Ee/Jw983QrZ/Oky
KYYew/rP6hUwJrA5jdkhPLLEtn+0YKWbgP7ImEAHIXFq09b1fosLe3RRovlPx5mHnXLSsR51/S+3
VjHBVNIalKARIpnHImuaw/N4Eb17Xd+fKhgPj7FniD3N5IXOfsfo9F4fYuR5yqLu3Ph05YjZzAcc
P1Q3VvX7lCp9qpt3xjd1WM6sBJGTDEkBdhvkB8WOGt3Bd4OjORA8K8YyTC7B1TgJRv/5J5xSMIhg
iNj6k6TlLlokAkLxlQxhUK/T1F3FY9pNQl4C+k+dgPcfV/XeNaUAiGJY8n4FRCVQWIV56yxHFXiD
n/nweUe3PNqYohIWGNhqAF1uDMh0dil+pZDZ3EvH7zBGpGUlZ8NszrzClkNpdbZGxW0lkzXOaoml
ogaNIrmMudy6sfHTCvxyzbshvUjAfGdEC5BTuioWgj2oEXYSWwcC8UCNNl8nME/yxrHSPMuWvYYd
JpZn5iQDyfBF3hbCUuWgk+0RYmM9GwpVbKwYXF/FAseueDEF0c8s4E0XHjSURc2fwm4ZFVsWJJBU
Dk4OXp7mqH5/B44zeGE2CtMkMLM/hYJOOOdKPTGgaV2A8ki6xIlid4UMXFp3mPkGXchhnnc1ruT5
WgSw4eLD92AtK/Hl21rDUMG1mt6i1xglw31QOWy49/ZAh4kOHf2FccIs6mxpXoQSlDDl8mErMy11
dtqfIJKdkLpmV7PCYad2qVMNrdX2p+FvhkAvkZh8c2VCFuYRimyKCW/wY+2CaYW7IiroK+kyVviH
NFjWGrkGxVfte4DCZ0r0XhTXEPdhUGqjVhBWc5LZKo9IYhqKmnVwS988hGIb0y+XlGBlS0cd+Vlk
XVhh/a032WcUuLHJvwR29xuIAQKh5PhpBqkAB6xikR6LGroOg/GYy6/8pi6aLAxK16mBiPrvMj1b
E3hoLS5/cQ+UnePFoi3v/7Yzwc4Ga3wFOLuhhOtPiU+DjvK+bcMYLvpWTuwXBCC1MRRkMKeJC3t0
3C4y5N+DeZReYDVR4epk6aC5ZzOb7klqrYMRaYkE8XpbrHXgJOlUDNhrYvmqyJ5zPswRb0f5pxoZ
G6OD3pZo7u2TW/DruVn3tDzh9uiSigVjQzDnKaagZFkrb56RJwKTHntADwhfNkBuqg0hTuS2HI5+
EexydcecYOS5hTZoj+eQ/QDWeM/CrkMhayypyThNByodBUXWUWKjZzFruBZvsybp1w8CilWNBfek
/aYUJyT8w7lgni89WVLgFRWQYu4bXedDJLD4LW8M8fYnqe06xdT/mIn4M0ae/WATpIt62ChsRIuy
owfhLRJW7aYe7INLe+ppsa/x0ZwRRmmYQ4DAbYmLhTo9QWhzpcjIwSxKMcE886NhHjeB5+uFVTDb
3Q3PiDSIX8oubJ8KDuuaZm9/X1gV1s/Q/7a93kmeFzxMp5hX8LTYopJ1V5fjxGw0g3nbEhXSo23r
6jkBfQDENn1h6Mi16kLICQbz6xOQV7yGHUNTh3HUPX3ocgt2bwd6fjxr+PCPoHQaMYP95ClinRdb
Yus5/vc69Pk9t/hrRum62qlLPSY+zk9Q+wMFXMdqAnnjBrk2h/yYJVblDH59rbDApsLlDZGwCR7l
QfHgqVtKS74dgdfZKIbnaRyqaU0WQrmX6Kz4Cx3Nc6ueIBBzMO9ArEfnJOxXLtljq352g0zo9MAN
WvdAnvVTZpQ42B3yowalxKcunzQlvsgf5wQeIh9vc4hXTuXKaisZzi8PixDmAvX/CO76OSaN4IGB
yxONOHzcjRakBeyrUGNaYuKGQxIWSslEp91gXqBqbUmIUdEcgbKuY2sbOtEnHErZY4qo6jaYKK6w
t3YpfPLPJGbEWil1xXk6Ppw+GWmCmjosPe9eb++z0lO26C0vOnVdsqHsVOb3xHSxzqvBMv4JhE0L
RZ5GiMYp2Jg9Yb49pLzVXm0m+9Ss1nxSGUkLuli9uO+MPsllNmoS0KS8LOLtQf6cSQ1g/iD7UcK6
68Kvosemf3dj7+ClOpx9ZfRgY7+/G8U04FYHqPRPKgS/93y5WtD76kHH050iQY3NnW2SzVaWsGC0
n5ydIV46w0Y7y2y5iA7VqTyW3Scc4ZyhiftT9WU7egKAUjaW3ja5JhnWDHEepTP7JMnlFpL/Efb2
OZOA1G2Qpy1xIX6ZDzo7ZiXJDjg6sFMu5VU0d6jibcSfKQ1gU2PM8uAnpEVw5Hr2E4LdSu3KKxs3
Wu3SvUC49+kRfgD4UhYT3eiRHYWvfdHcMWRWDLkOXlhJPMK9ddIW/MJ+TWkDf9OLU9Xy35XvGYEe
hthBURVi92G897Jcx/eLYNYQoOgg1HGqu6BzdCOKuI2Ad4c8XCv0U0+x6MERxRRu3tMcqsQbl5Tw
jn2KdmPuzzHi+dYJH4WcAwv8B6yzfGp46sEuJlb5r/pRid0kIvX4Zxw3Ehh5SrArjfqnRPJHZdf2
E2OENCyF+4NbeUAVGk5H7FeX0ySH8jc8y/1VkWRT8wu4MrVaflszPk9GLkmobDDYH2M5mnRc0aaY
y+PXpW6RrkaCAdV+NtefOlX5X442SXqfIZCFDjvvy8XPVDfC4Ce4bYhzVj2Ibqd045s5XgcfSwSQ
WfAzkP1HySnVOyAoE642vmbjkliLbxSUXdokiGfEvxNHk5tFDXA1vFbEZYh7VwJNPHx6MNWH7cNS
cg+D3E6FLO++tKjaUQmgfx/Mu05BWhi7YQjUzcWj76uk+ZylgtdsoIQ1HoBwL4hPzkGvje2eHTGW
L4DVlnFASX0Y96LYuvGOlgo2Qpo9yn6+6uPmlXZuTwl4J0nO8S5BUUq1DuzNMDgoLEcFSlrq3Ejj
p5xIv4z8NcZq8qARd4yDfuIB6BzTDfS6jssYgP4+nsMOh7dOa9QtYYne0iO6jL9hvphI3TLnUi7P
2FWF/YuWWhDYbyr+Ng0sHQrRh8G8USm4LsWoh8c7jNqInmSj+FxMhQXIZIiZhky+X9aPZWfun6Nt
ZopY63cZGctN9sUjXVb1ELz2+Fu9Ap5df3m3NS5+C8/a9hcQCO6RY+4UavQgtrCJcuImsD9vuenV
kejkEFCKfTQ/lEArxMpBqhTfnQ+fWtKFkCU1oVDbWBEpCCL3RJRirFClBgKBg0vYffPfFm/g+q05
gFALO4AllanTSlehKqoU74AsUGidGxpBsPl/xlT8FSUl4Um/idEz/A2yxX92QcqxSuggTK14EYFC
CiSEE0QAHibPE5nrl6Vq0rPKxyaOa9DoxsA9K6hZMZcFy2TXY3FkXFCXGk/Yc6jKeRlLxNye0h4b
wNfoYW74Kowv3Zp37nex2JPqDLTcHHdWRgRwmDsSOyl1UikJG/5+hlGFBJpj29HiLGCvMhmrqP5O
vME9y1m3pnnf2fFaP4M4Xupdy7ygYtJHOYcQjx4KKoK9tpHHn1L34O07/sZAwBPL++kXfk/DK8/M
CnE3xJsSLuk4LL1/zxPKwcnwP7d0k6R7MYuCFjDRsV6oSU8HAS63rN/6cbg576Swi3IxGSXiNSpS
WuvoBrafT+mMudbnGWfHKuIk27bNNHzLmz/mlmaE9+PtQ3oD0ZNpasE8D81aAGvmwbTT2k/Dy3sF
xU/4gZl3H1pylYLhF4jyzw8rYkr4nHcEMvg/RrkESXQhhV520jm6zJhaHafvStdTwtocTlp2tqWB
Y94MnRidBkUMM2msKtajAZPsqyn9irfx0fBvFQfnDTJCrwggJJuPKl2Ln+krU6GrZNN9C/QD/HZ3
z5OlI/sHzpO4cUzmNsDM0S0S7oZgwvkLBTQ7TNVj1LSQAybtRmyBOnCaYHvO2pA+EPC970oQ+KzX
dJ1tuydNkI6mHxzbCre4D2lpuFSA23f32WmFxFXfpIgzB4amdrpBYnEMF5awS/9EiP2X29CG4o2M
SV+YdTwmm67m3Rn5yF1u+NKP/GFJGhAfPlWk7gi4nn9RQ6m4lVXPc1Aa6HjLQSOzj6USTna0ZfzP
5inWCUxnrXKEAKoppEGwpiRlJ2JfwqjH/YdQwhkZM/uVlRANQjnDNXmW9qH8PRX8FPXNnFKxo8hc
sagx/DtLgmfX6TTR3PSOZ0Q5HqwKDrCYuEE5kJmKi/YMqYqKi0DgKdkqsDHxx6/SES4BL6vR/w9W
A1BEUmei/28+nT4ewuYKwND6RmLrYbv8ru1anZRmb2He+yMwa8bN1OcXkXmRyRLwshIJ8He7uOjo
EFWXl6BW1zkGuaqeguHE3yEI98AxlCgdgT3K5chhzcwBLz71svxTXcE5AuZja0uf5lJcaUGECKeU
AM5/t6aBp5rAJVAdv5Qb+AwatQlxSAzA6Fc4gAq1kh/Km7oikEsTUUVqMQtqUhglTNDn/W05yeyY
QHueKecMtOi1PBcx/9tEE8Hsx0iboZBkC1wRlOBZ9YamUojTWkpee7AUYC0fK+ejx9JblBlwIUss
z8lNdN9d1A7N9Z5qyO1uUAhTRzIzowrOjOEs9BeOfEaz6oWJegRd9b86FtzQxZlqgS0B1ey+qgT6
v82qqMru+u6saJAJueFBI55HkD2141sqo7k1dCx9AZxPTObGp5zbb4XyAGohA8+GAzauxWhIZygd
rudPaFCN2eunrCzd7Fe6ObKB9+Pold5Ev2x18mIRbqOh2mmMuxsIdHncfhtOkvULtQeWIKAOpkHN
9ltMWSSOmhUaX1jid0jw07OSmut2p0OE2BKHZZfGypsuhGpZZfcgF6Taq/MvLn79ZfxCblfTu17y
sTP0hyEWfwwop2Qvjb656dMDqlusXtnabwfguGroVKShjCdMwGuFifLq0rhTZ+RJRMdCGfXIqj9Y
aZqsE0QjG0nqLEejHuGZdzrLh5gH5VDPIuVgnUfsFaNnkd/MWssI6Aw4bHX0VB91/bNR61/0mNa7
LFPRXAeujh8owQM0fAHSsGXXu0na1AOSQmP0G4r7JMTlBsOTbz78afQuonliMWNfnWqybeealP7J
oIqY33ebs9pSP43YsSz6UZ2PRlGMpQWv1QkpPhieZgy0UrjLU/QxIBJOzfvTKjfQ/1NjtA1iLMwn
ahbGs/t3QRZWVSwsYDgJvXFny+pokDTTGLHxDe/583uPaw1+/YyZwsLfO5dTVMlt3jHUbAcNjVBB
r/5CdDDfyvNRIsHuZNOzW63P+LsP7UJU7Qm7q+isdqCXxkfbY8W0YSTNEq155kZoVha0vyrDUyz/
MCH2f5UJpySp5xYSNYLPTj5riSn/Zza5YqVd3B9xqZ1sjacR/znjN4/uthS9/NnC/ezYOmO80N8e
fvpIySp783iJrTmVlNzw//6uS76pOr8U+DLuVY1oEnD+rlB/ghiO5YbLwZZvd9TkfzBgF16xhpfT
jEO1TunFGNFKIaFagWbL
`protect end_protected
