`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Gy1bKdwfkOwrVNhaKcvvIZKO8+/R0WH+p3vmFRvIRouJ1kQRL880RpRJb51DWTVNc572RH7w22lt
FmubnQsytQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cptZRwSfSWv86xbTzDYloxfYzXCdBXxVS4R/01WRRdPalvsctpvFhC3ERManlqltFltRfQbB//G4
59WtafJd+4zlPfC0u/u6HRPjhBx/mZLONcXUNh0C5NBojEcMtyv9tcyRkelL1MrqnfXeljULLH2a
4RQiVKyQbkoCA97tTv0=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AE9QJBEg4nBxW0EA0pwMPZkiB77pjy40C6Crkmqgps6AWs4VWZYRFULx/teWb3qlvGDHFb5Vs3Sm
4ixXz8GiurwD+glOgoqsIijQbe+Q6L86c+1lnTMdHV5IbCaWoV2Bo6E7fvo9lcnLWOJw9CxMvqiF
zSCxd6jSW/rL/uEHrG6Z+mV+sj+5mkcmUq7UKieeyp0jI/FAox7UL0K3xdMsJYCgyVDoAJafMbDh
8uHhopEkCZGL/PdKgO1s2TjYM9R1mLnL8VLGZmnHMsyRsp2A4bSz+71pvqNai6eR4PaoNFjvkW0G
EsT9eDDxUtklKP3fTvepmgqDRrLkeprGPm8J5w==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
s5ELqUDgjsFXRaTB9d/oSqrOdqcWSVf3VcaUbdiYVmSnqXhuyUoCm60RPjS6vs/aHeV0TyAFWT0j
grgRXZ7rhqdq6QLul1o7rivd1EaYwx9YZmvEzviMGG3uyLwFvdbQYYz77UZxCpilldIBKiMHe6LA
ZjO7vyqfhv2RaBhMfis=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ph3p2XHeSe5TNcoNotnxhk0Q/EYwzAjW/AjlME9a/HUzhfJVd4MV6v4aBy2hV7gPnq0halfvmEyt
qJxomFlaivJ/3YcQnIDLOM/S6JFjvnEPbClDF6mj8B3M6AxGuPmSkAs67+/8d5DGY0mdyirfMp3i
7TXL9Sh0ZzuYXpatpkIHVsLoeQ2QruckK++/1To8be1EbrEnwqsZqt3cxXe00DO8MSJwrz/vxFN+
Jla+PE2/PjUhrm+Y8HHZuAWE0qV2DaZfsjwu0TGZNZ6lXQj/758koobmltDgaEHGyOjFjd4r7xO4
Z4sVwCOZLdOUskIfVy6xPO/fSjOXLfuRsW3aNw==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g6xnTpZsELkh+D+mLYUAIF40MPA4fUYcUmvrMcvS1wwKcNi0KjNbFftbBNl1Hwgc+GD2wMBnTw2W
nBLKI7rpP33fTMmvraIMGRUWBECo5VflbCcfcdiyzUxxQFIhAXHG48syQQZ7uHHE7uC3zBiE+Aw1
mrDf+cgBdPtLQe46XAcuNefQ1v140ADOVPXi/O70IurIVrZ7rPu03usmzY1n549gKpzEf4xbBM5+
9MmEEOt0wn43d/hEPlkq2Px2Lla2mEkNm0L5sPXI7cudTDkJ0AfyliAxF7Qg2wEWRzwLZXaKzkwc
yteDcvGmZgib7V19AXbxEQi7Ooj2DkixCmBceA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18016)
`protect data_block
aHPGuA1lf5zO1yrhLrujBZ+HrURwblXM0wc/NOKNMG4HSihqs9zGYtz/VMvZNADliUaqFVsrrtzC
DS835lVtQy/vsJZgzAwb9zGyY3tICpVPFKqvK+dcLUmTfmKWa7K/tBoc9b208SPpuUEJZLgiOa5h
5OFelLptLEvWIKdc/9wr5BEOrkDUxHEVHmFbMea/bJVjcIuEGZAhZiOMjCWUVSksItvdCI0gk6lQ
SARZx/KpNIi2kl4SZYdxNTVHfMQ03zOPqfIDzGHsI+uV4g3JqlUYMMwuiGe4UFkxFTWcz2qrAzLU
ryrg+6Ipb6cmF3I2rbEPyg1J+kumyn8akYRUIufdDBZgFgwPMU6V8suEMC280m0xoVfwbTstm9Ef
z+MF8RuMLP10+kc+2iCbw9x+NdV6t50gRDjMClwg9D01y9D6qlKCX+W4yqNXOtW25T/z57yDA5mA
zOwb+1tWYbPjMN6Ljht7Ivv1/bbisE2fOcUBBf7YBqFNAE6lYVuTE19lChfP890L07qBnBHJX6/x
RiwrzNvNZa6M7xrc2nU0GLpQebRfT8SkLlidHv9Gy62SyMfpRdsxpXLlOHSkSxEpfPxCt0shLDf6
lScan/u3ppppkwu6IWgr5S8JwO2GbwffSjB2cDUmCFUrKYrkLgW85g673gAfS6hDjBcNJ6mxYvYr
5ZVahEL8d1FfQ7NyTNt7+LfH16fzsG0jkbjdA0Ni+w26VuiBHEo6xj2p4J+V9LsZgZ4P78bH00nA
QmAi7+BC83MHpmYxr56ZTR2OUjBl6cp8Keyt497xfsB8O/zlIQIWIRqDC599ATV3yBavvBO4FKYO
f2/qrbvHYrkhmkaF6SO3knUUv4wUt5pMxr/gBCwMr3yAQbsFjd5JQNrogG4vgw/lkoaDVPofyYgh
OiGtWkYsudaWND7MpbpSix7xCh8coYnF/71LY0EuafQo3MnWxvb9u+2orlHPwY5XFGON+vEL2omU
guNfaiuWpxOjTHulhIqC0hCMGqApVDKGLjoD054QIY+uDhUVh5mCiCP2n2yJPKTsBoyv1mYs1Slj
Ua40ThclKKSYVgGi/gZgo/uzFRjRSSv+8UeBzNf11FItH9bJnvKDcHtrR4cNrd/pweKMOdY3bj2a
nuIBo5TZ6ykHzb7Imex92e71u49sXCuK0VDHytXI3tXMk2ZatO9vRroMIriNeOcwHI/gW3vKyG54
2wHP1H1BmvrGedFMEXIZ/e30MQk8qxyyZwKL1LSbACF3VAbGm6REd5aecNbYRtlaxHFwrxt4Kb9v
7EfUBe5i+d06F+Wf2efh2+2M4kbY/GvY46XwUu6NkpaoP8ukZWHgoi+fLbCaBitQGzWu4C5L+ky2
qn7b2c9uf+vCv8M/R3KEzAX6Igea2ZaYAWrFVWfTG4Z8eSxvrh1smwS/mcxzkvRcEbSnYqG8/3CK
H/OTaHnA8Mm/Ckm4SaTOh6ql2wKND8ITdN3eOpLuZRima6vXHHZZBaJP/epbiF4v/0oSfz69R7fJ
myNKyeqZDC0cCHcvSv3hZFH6o7NZYyKx0q4sVNS6Vkd/hLoDFXFY1D4l1jfZhSNd53AbpAifflHG
PkLypS/z7KvwuJ/E6/a1o+lYMeLjiN1WyBhgv5V39uEhz0apenmBSKmJ2uYICYzlCNRPnxDeDDWv
6M6C+NexaJnYfGSC/VErNLNCpnG0Eavt+KhlUKn2KLReN1Dxt/AimnpCHBjhFEXmLaDizXqbDxRw
77y8M0MBKt9kp9se6mm6h4iMr351/A4tsTi+q0774Jyb37w/U4e4McyqQY7pQDTzF47MK3b0yt48
yXR1Nw8Ro2h+TksiAuNZLRFHuVKRKJITtxDGKtEC0kO8+SFUv5CZM5GZE5L3GXY81RkPlNQL52A+
EVKgZIdq/vwYkirZRn0X/tNuzOcfT2RFUwWDza5+Hpab5Y3yxPQr94Ciwyj8ureNWJzJ1VadwSM9
6YJk92gjeIHlBDz7SSOLOkEnp2C/t1pF80Lkb/prVMMXCX93VWnlrqIBPPtga+XqpD6NT6t0+uGk
QXQ1EmDDPCjVZGe5Hoxisrp1HpvgT9+f/8YWCgFiQJprsBjaXV78mS3zkFv/wLpSgQCdyth9Al91
cT02TgLVY+7f+/vOKM5lWX25E9iN3to0fAOY2yi4H/oQf18AUBc9D4zZjkyQbrI8oPs9p4o2p/3N
wiMa13JO7Km3EPLW/5HxPDlYTT6aqsoJUhQBW+NNxv5t+bIe9PVCVktsvssKGET9FjiYW/eoHRYh
CgjQQ59YdPGKa9RbtaVqZ70OtfWUjXl9Z1sJWaLmjpiniCVA1zPiNpeo12kRFzdsAYH6NvVWyROU
9HwsKYbVnx9J4NWHNQnl+BUR/uYvbEZbA7ofQeJnjHLm1RTsmzLm5lY98qmI1M4lHb+yito8fdA9
tjT+RaOwGHlE4gLtHkmW1ErTJ5isDdswMFAGSwJmch8VEegR2Vbt0UcX9UvqKW0nRr6uX1TmDZEV
hVsTgf3ROJmKkFKAlZQJsces94IMiocqwsfX5h1L4piD71ZcdYTNvBkNUMzcldKvcLbWpe6j2iAJ
3Y/Hw+F3rzN3CmhC/77cE6Gxb9RNCdcNf8khOjsmRNvWfT4DoGAtDacXELOxW3HR4OX7fgiSSDsp
Fyy8tsasIeOEuLOdExW0HNmK7c1Tneu3ho2gBb/PP9PWLjvEiYhKSiwtMw+udU68cjL7iO1hmtbw
ILvwSZEQUpNtl2Q2jZm2MkikuT/1yDcflSF2bz8aakwYKkayL+N6A+WVzOB/uUqjW8Ao2UXLbGVW
UptF/AB/WSNeScoe30Ly+sjahkO57kAhhfgTg3l+zR/XZ6DjiA3GuhamB2FdJtKgydk+8lcSgqzg
aFGM9c1U8y+0JKP9vifVxuHalZ+8hpQMmRlX1xHfoofc9/W36ZTrI/8eDLrUIVExF1s3yCBqZy0u
17o8rnvbTRG3UPCq2bIl6PMYlcCapUy5b6SfhNykJeMCf3BkH4mIUXI8lqWQQu/HdxSbFKI5FmWY
4o/2SR679jhGn2kWqnYf08vwy6cMzXGwzZBzjB6653QC79/rwugPPNfi6ZsVViT+ggvoYRFEXz51
M/pilLjTjbDf/R374JtLAS2vHyUvR8BfhCuDIbfJFozsdmBiToLvHFLjpFTeGhTSKkSn58NLv2GY
6evgTEz0upJoqdAeh1kGqbnfJBJ0x6+8TXRSZsQMeFLb8jS0IEdn5f9tBG0xDz9N+BJaeLP9EiZz
/eyR6931zlKxSYVUWr6Di6HjidILw+ZgBNt+Jfyz1OXZZYQoDqTHPc1mNBY98h8GMw9vcQI20Qyu
Q5haG2ENzVfA/gIe2tgMIF3E1SFczSBQk7K/ZmS7p0BLylBmMM6/7HuU3vvT7vqE2B8lO84z99wC
vTiLKZGceWSyeGDw0MOO+76JVqk13KS7QIWUUF7CcR0t26BfwDIMYNIGaXVOW+7VoDCTbGiYfz7L
uRKFtR27cFEdKNXJLrdVKQKSctkSiIhqL+FUMRxxHYpc9fec2HB3MbNVzAQ42svi50882KIyPi0L
y2WqUEV7Lsj6y8qO84hLGiiuB6gd7mFcpUSJmQrOnQU+D2ca2yvC27kL2XgaE7LSeFyAEtilb78E
PRizMSmzkJ3Cu8U+70uXsa4dfor+aoCHLxZxiYZ/sqDZfrOeQxMInrsJsOiSQ/hoJ1WWVDLb6kQ/
jyoPsahI5TV5+hPaHxu6Pi9eWK5jCEXCV3oOjE6/4eO6QDEgP9LVOgusOpHdFYdnYwIf42kbgf85
XOtLQBjB5aelKqOMMQoDnzAKpVBX1FzFovRMbs5YGnV3ebiwqVMFrUgJJz7asymCvbzVUWqRSNYW
aG2FGr+8SkSZmyzH3Kl8yCk4TA+o3QAofbymVXvFtyBUpz7atj62N5U+6RCw7MaaxP2wpoNC8jEx
lL/R3Rg4ZLYhPzFuin85mVLZ8d3tnrSpHOgpHfExgKapLfgIbacNU/73zRTgjIdj4+Vk9kM5S5uA
HsDyRkvA5KyJQt4e6uGFiexU8HuMU9He1/Y3OqBAeIMzpmPTgfukcmHZT1k6lRvv3tChh5HOnOL9
Jv0BKTNWOTTgnNsJIMp3m8Opn7fcPt8vjUYTsboISssUqzte6MMF5SdV8QlTgjhg67xGXQbuFA7L
lxZSmfBk2wXcOaJQGD6UagUK68hbqSXA1mCmNLLltsfE1eLNypjy1SrhHcrWwiWmzYf0GKZ+Amxp
iXR335G9POztohITGpNZp8wVs1JQIpNEqZK/RufD7B1UdH6EKIXXnjxz1SxMk0rWOxbMhMasCKC6
yVwjsYqBeQ1cDue6ISloOXEnimTOL+vGmSSw0Mk5A4keU23BC0G4HkUSJsm3kCfg6r0IfqYvXXRQ
Ma/7YAp9p/FwUXBHisIkGOaceQIbVErulsavue19vRHCspBBOMY6d+VlGi98q40y8Hxki0YkKYES
FxDElWYKGOqfcrKKvJgd/NzjfiwCVZOEhVrU5/N3Hnx8RKJbD2hTXe41+y00/y2fublD+qgTRlAl
FRdZaP/4fnnkuWzatUV3hWaXTY4ur8qYEnmRvclL+MjvEjSiscYsJVaIaYHsu8qyHshbfbSmMOtT
UfcCJYAHGC7F95NQtnHCH3QhyslisrVrn+OqAmZ1AjPYka2nvj7NyGzGagTrZG4R0DLPgThxXlEV
Dp2YezisLhrCNoNXzAClW07cFf29L0Exb3jtNTEfS4OlWdZ3qoiz8Q23nQXQfFcqRvEyN9LZ3rWM
zs8xtIZTZacZBT58VnyGETCZvarQhk3ihmCwcYzCexJPDWsP02cVmpFVrf03nSt3ZKffYJWPJ6ON
Do80nHzAAYNadHRjbBqzmwc3+5CAM9CZTM/rx5qTvWeLm2sJsjpbpkgmMDxj8E4Ydust5gJqpept
c8EQKGaoQXhlgVNReimAQAQKaATmCQg42mxYLR4k1zbQw0iCxvPAR27b5shzBcbH/kvUbsS2IDff
zFg17lkw9YhFG0ZWWArlUAIKnoSQl+x/2inftOV6NdZFcW/zrDuaezWRAFkQZHRgWMSgD+3mqlgD
3xO9yZlf38OXgoB0YIOAvXOlthRIuyeioe/Vz6n7O5qO8AT7JzOsJZvM7AMw23Pfl1RsMckLN7er
K/YLqlFH5aG0o+sAvhJKLY8P7TJJm6i1QjTMX7TwPy4kDUpGPJgL9RwmRKCV5lqUco78EgESo7rA
MojUhHMOae3poK5MjCO+FapLGJtYTgJMmjf0Xr9gaBqf011tbX2YR2ZumG6JKYuqirPpQcGvVKVW
Rgtc3/HLdRgQphSgZzY57dkxgXkBDUSxr7/t/cYAaRsBYKLBuFhD+x6zepN+sVR67ziYamxa7tMW
DwGprjtSWjI9bc/KTa1cuGjPgdMpk6+UUbzCD1122QgdQ5Y591qlJ2gor0U3p64FLWorP6C7jqaR
qOI4btOu/810x5vBQ0SyuaZhgr6ceTBbeZTUeVe6xAd8tRWDhUyJLfgsjMKyCjbMnks60hxcs/0M
l93c1p3t/NIJEtzxaGlUOkdIW4p8iEvzsRSo2f6tLZH/MY6ERnX+E+8YvFzwUyGMIUm31bZD78Fi
OyqZ8LNPYjVJwxYRApRbHiJkPzMKmuV8lQw9h/XDszmMvRjXubVjX5wZeQmXjgDYNt5dTC5dtRIQ
LED69VGFBZBio1jGK8huAuOYIcYD8PNeDm36cK0xOEqYcod/dxL99reoKAGHSpM3FFgPoIq3SQmj
4ldyjNV2pkLoEu+G/dH5UTaAY0Rb/1yjkGtOvMojk4qQOP8x3SLh1Ow0YZuVHcCIeaJqTBPLL+WW
66R51f2eNLMY+/yQCWDOcTbU9x8CRTSkMFy1CnMPHH9hUec33UG6vnA1JCkuDTapUcslmAoeFD3b
MOI4UwlHwFUS0ZKgxzuVxP187sEbe2Pd6Z7DuudfKZfqTJ7/FpG9096CjkysBNXLOFCmJxoE4ew8
tpkBin+TiD/iZNp7SrowmYy2xBIbD0DZ0dXZuHr6NlsADHFOMm0oxoqxk+k6iSLRK4G4NfOJBdeX
wBdrMB37XI/1RbnUYu0m8TzyzL3a4/gh0Kx/K/d3PIOI/kfikYzzVtoBc+J853aBFJS9miF9VywB
jYuDzrBcV1vvKGHOazyLoEhPljeSbpPvy7jaL/fxtsN6sdWsTrP6t8akxtimaWgjw53JQQlDI6Fb
25UuEoWIb9HdRmU9jOJMR4XEQKgU2yPEC/4Vv65jhKG2ej76o4xcdpDrMJo3e7Nf0i4+CU4S+vn0
1A1vBi/CR977gMD/NIaHMh7Had08E0EAUY4OQtPVmOoeSPl2jm7ITEt89P5UZHjxMRSM1c+deRgu
G/M7ZSm+P4t9kmNbgPhxkxJftiMVXGkF+fs2UHvH6DM6cvEUMc9fF14YE7WTzulN5tA21na5ahTB
/JBVQ4jggsjO10JFu+MxEWe/Lt+d5ue5SI/T+4Xb3/rz9BwIQxMF5E4ZoWmsC/fO7JhvtVWcSIud
bFZ2qxz+7yn3Zgr59B3jkUxyB0yBdkrZg4hnR98KUX/rchFmWH+f4JCFrnmlTSklSLD7b6EBOi+P
O1b4Pc740C8Ia3tYe4tuvs4EB1J2YturLtpv9HeUWRIBAI7fBW9p7vOwtafig3lYi76aaNKc5JNi
bQ5GT0/dJBuUz4U3W22tfuK1P/s4eqXGgbUX6CrQFDWOsyEEOQHu1wQ6n2/Y3pTeCG3aC+sp4QoB
2doCxLJ7leck/hr6JBp1AMozdzm+bzCsao5a9QDNWRD7UpolHCmu+dElTKJqhpaEGesktAXzqP9F
bSoPRSuSmZTedt8j52Nm+v1IlPIM4kDImjhyIk758ABZHSWj7eDF1LFCKFzQ4LVo7f+05c5v7T/C
AIn0x96XizECjLaxPlnAOJXs4JKtLsgl31K7I9/rmnwyne80W94CjvIymylsYgbmPcdWXxXexVUI
B5OWI5s+ktSSHSqbD+E9DT+jWZ3puwVPoNy8J1dl2SmAf+3xQSPMUh4eCPz5YTpqUoJ2ZuUyhnWB
XWd5r7tnNEWOF9dBT4xCZk0g3nxSoxlKhRuj5O0buKO4HxNNcWkZ7hKBByC4pXpRWV4e3dLZ4iW7
EzERq18lpbrEqayh3JBqvX1ZD+sYOkFdHr9Ve+OQ86ySwhaZV6Bz3fV24QCku+NuY4DldJ42n0D6
db1FPpU+nopDvG3elQAyTTsL4Kodi4Xc4Syb9F+2T/CiHVabrkR+UsAHCkwx8fxJoXkCqRdhl/4m
WqbC7n5r87OVhzt87nCjoGkLhdoQp+gkZvHwOYbXZDjMfeDgYl6dwj6N/aIlc+b2YWe0fUPaSB+0
1F10QYPQDZGHdSthiDXA/ijoFXTKMFvR/RwSmlGZ4vHTQGde9rUn/+Ys2uEQF5PA5DPyomn7bG3S
sEBDN8iXdCCQ0VByBmqFlhtLiaE7KD2ci12dP+ekeNztczWLODls7REDD8H5xm68sYNXfE1Yu0AC
uomUTp/Xqi7ACWGKbY9QdOdcrlzmG6uJ/2OUH5EQGmdTiRQw0itIB+ROzf02A73uzYYv+79quocd
pfuoelr6N7lENYzQyVk5Zklgu5AmcUNFE7DXRam6USOHVOOmEe9P8chGmbPQn1A29WL8OoukvQMR
jT/CMgvp6PaXd8hrq38HynBYMBctLnTW6VPju6L8UB6JSrpPWEvyVImcIfkQJH7R3BnaeD5uXk0K
eskdlxQwk4sarAlq6THccZaXCSZiZagF5ncQr0k7bg8eJQnopS3Ni4K1nM6vJOdgM1zFfoH1mSkj
hq35xF0ij6g9KhDnleMzPirKpHmYEfiV4zIEpGDUEDAUwqh2sv0+/NGDSbD9cOalMppljtleLdN7
0rAgrJ2Qt4oTsqBBBmzwRkCDQo4AXN3br6/fY+2hNQbIToCK7rNvMLRkIKJPEsqzQg7MLRyuzrgH
bFk2Xp93hTRuTkluKAF4AYya+lwEUUcqQwAmgD521PxInVhP/ruR1WxFQ15LaaThVRmVSW8RQ7bK
I/igU+5+2facuKdOcF3UnTEJpOOzLpVAaJwmTjsL5HPHVIVZ3qrHW2nqTmpwCxdgF4oP/oEoAJn4
qD/Ij1enVFcBU0njVk7Ov0tQGHRWCSuvFEV3eYNk07i+EJELj9nwDH2AITZByhJwl7ZcUGJnS/qD
3eu5j8o0lLXdiF2d88DeZpKA67lSCmf7QyYvHS/a625McFVV3vsge9oCyK8RTEPIKogYholGyQnR
aGA8pUfF8UQH43sXXLOnnT0lAnt9xR5yJENTUxQsRiJSXQ78aRnz+nDr5TLCx5OW9MBAJTlUkPsI
PvC1nF0d+exD8O3BH0oGfAYF7y1BQnoj0x6a8Eiv0Yk8KjezlU09Hqwn96VNgOhsveMUk1BxS2PK
Cljzs5I95E6T+fIaV9d0wFuEUy+Pl2atolG3+lW5Tt6sCjTAOdIB4+GlH12fvR9uUVhB+xWkErHA
hmyCI1psVPGnhgtwo6gsUjtgzUciKxIH36TAWv+fhzKhdvFgy4QwBxR0f5KRgLp3iegiIPal8zyj
9F/K7affVaTy30xJWVdgneDFn7GekKrk8kur13iSWGQjflZm9h1aohUx2mZ+4ugcWPMQPLbHeDeY
XOkjupBNO1sFdK8P20g0mMtbr+eG9YNehqjlTHSnZkM9PZCV2iSiCr7rLk0uddfTXCpMAtSOSIgK
XTXdGEfj0/sN7xHVWgPxqRMNg8rH9Z8NuXwjf8X4h+hN+XCGRHfgX/QBb5GK8n6ICRsZLezBVfD0
qyBcy3NjFQ1WUYKDLIvrh7jc7yZEM6Cj4BAeCQKxT5rGVX4dQv9UB9zT/kmaEWru3yMujkchZd4I
13CAc2qaZIy+dsrgPr1OdXMEHf7SzHn+d88UP09cRf2KDT1bMWVbVOvKkL0ZVOk6ucB+03Zxts4z
igXYm516MO0Gm73VjAOsVsoFKYqlRnHzSYoC3nGpjsX+E3dlv+Ckl54TRredVaJwMVvGyHkishyy
DVTwNk+FLjDqZrVOk/Jq7YfEE5/myIVZLrC8roHwLKHAzB0NCDDLNB0eHKpckYGVI6842zQ+KrEY
PtWEVYY6LW6wl+Z7yEwkPs8HrTvpRPktdxCtp6WNYvG3LItnH+oxCFg8CVOSjOo4JFK+56eE54vZ
Up5nIKdqzTFROT2WfJWkeBywvEbve0T6yR07+zmP3u/oNMj52NzFuyYWBmbbPTx8jpjKvy7Z1c3d
faJ59Za5WTYnd7JGkyhZ7h0bwRkwxmq4qMR4a3Vfkfuau4bZoi57khyL2o3Ms2BxeWUZj1bF+hIE
pFYK2wN7PgsNQa0Yyj5OMtymy+m3t03CqWh6mgZU4L8XhGzBnA0FoOUDgiZH2WkqYSLJWdcmDeYi
T+6371x1pi4Az232um5KPydz4LZHr+3oE1GX3+Wa1BcbRM7lt+UDDnk15466BBprTu0uUv+iWAKC
o5e+uLBwqZxNf3ZJgdqGA9S3lxlC72aL/tkJzG62d4NJBjscGrZIco4Rs/ZEQpuyfdFMU+QBpOey
P56AXT0ZDAYT3z63MGag+UfXI/q8PAMHyZrmZ3GERR3OQNMEBYpR0rX71AzGxam++LSpI/2BRBhI
priWZQ9y6QopqqafQLQMgvm081iE4fggEqGy5x7bO7IqZ5JwSGIR0I6WLmrVTrLQSySob5r7ztaI
sZQSgsMQjFSdt1guB1a20mDyltbM/BlPgnN6akEaN9SsQF/3nzvoONQic3zfElq/w0DTc4UiO2P7
N0bHP/Kf+FLe4SO0RaM9sVv6nXRRQ+I5QuAWm7XiKARQ9tgBUKRSpcvYHVUxi2gn0PtFT01C+0X6
E8N2FrX0m1xige4DHQfRKfgaAUXn88FQAgDjP+nycFjRzZGKK2RZi7a3U4gfBT9xo2NmIlrMGM59
wqK25Oy/ufjXj2tGyYFzESTY/254qYimu1XCQB9B5MIw3YM2BOFuePBFb0uKhee2N+XrTEYhPTt1
RZBP60LtDBG+nYNILoTzdTFn1AYAg7p1QkPAjFizFMe4GDZvlZ0FOuNgkQIo17WEzTOgR/94hTLa
e9krW/vWrp3RQiMlqG0GusjMZvaMEWfTz1nJXTr0mrDxGocclvNi0g+mnFhqVY5B1gpLkU9QF/Sb
+K66kbhfR12LK8awfoHeJYY7XYQpbd3p+xjjxhLw6P4V0QDkaFmRQZ28Gq5crwsE8o1QH8rmSl1S
750UnVn8K7Hc56uhp68Ezr6dml6U3bhp8oQ/tyB1Z03IQp0Pvq5cv7A4IMfrPdpSZOwAgyuRg1Vd
YZVNlTfAA3E2HKnxyMk4o/Z6uEogsejEsJBXgPtFanLjq8C+gGjUEkLnM91pbKlV4E6RJxsZO0Sp
Q0ZGAfK9jFJSepXa0gFNcgU5wWLE8t95iXg/bwQPuL41cjNmI0TT4e416yrX6xBYzR0oTjbhShdG
iqhA2YD8GALF6MWWRxvltO5kG1CMPCNg7uFPQY5UDt61/nNGoIB2F7w91biUSm2c6ZibMoMPmtfD
bOcPDsWLTaYTF55QjDtI2CS5xevIQd6dHvUcEPZIFZrwRBR4W7t62SblQ77y+Pv/tiW1qGRUBXZk
iKN/r9H+17xXB3qVJp0TPPbgiQNeZo71bOqVkPOgOjyh+XETfDi9Swqw07mDuauHaPNK6kYSvdNR
VphJeusyBTg+MW6tiPnHo4AauuBuj1UzPzo9pcWOySVJ9hM/3/w19DfxPQSczHUUV3erR7XSTf2F
UhAR3I0/SWJ//aW74pUbPcPVffmnktLAQbEaiYCZjFZlxe4/xuIB4Gi9sg5hFHAf7kHaAMrYn5GI
idTuGyqqOZ+Q0TaGSo982LllBn4uQrXiIbDmqDHQEic2TnNvxJZ9t3AJn1xwWrv2I384IqgReyL+
qnCZQePYRxq0L+rA3HgPBsGBE7LkvMaiRyrQq6XVaoLuEsvp3LvIQoIF1VkfofnijktjTu1SLn46
8qRmYz3SMfOVVwf3zrVs4C7v0r8/EgoTwWC5rPazYvMocg2oA7M10QJzXAGwiPGvHQmn5XoNv0nW
eiXdZw8mhIBQJiyMa7LAod6ClbrEoznlhg9/6s+tFRYw4Nr+XwewkPKScfgrFpSTIc5EwypOtMEl
WVQnWu6i27a8hB/Tbl8aimLpy5PTlxZoD9oymfKLoWCYyV1YQUxtY/FPNclf4tl4ZzZjgaB/LRoU
sHMmQsHNWlvJBvN5mbvbYuib1W8i5SWzoxuJ0gUFMpbfim7vdfwj/enE39um7bJkSdBsEvi8GbwV
HkhGnxPDQ0LULz3GdndXIJFstdaWy73ztLkV62G6GUKOZs1dMkhSLCOo34VPk9yHA/iAAOg8RZCC
0PDmwF8isL70cjRdlhaPhWBPIWEB1SN+VHiUX3vGq7F732FrIbToCsb9yN5SiePutfQlAASfvX5q
lXtuOfz00FaeO46NAeRVXcvotOy6IsvgXso0A4DtmYNohtoGJNzzP1AL2PUrTNn/jeOLwn+0p8je
SOBOcXiyB8+Ey18cFC1ahNDWlXg2Yudao6p2ThOeFp44bOrJOYBjEJEvFlQlfwCahzIhhiEjEa90
uvcycbo+RYA7Xqgp/z4HAlUg2yR04yyN+Qgt6irpYLvUueqoy7oP0vRtlCr0y9f6eLdbk3+om4R/
t1qz24cooSJzFOX6oLnY6AOAYQaRIUHf6shOKflTc5O3bqKcOyUigPSwOw3oWDoVSp/he6xN1j6F
I3XPuWNPiWIZXk1BAC8DeTffR4xbLFR7ogWJm2iH1A2SRDPP56AOIRUMAyIYG+lYp3yyjuWuALB9
S+Xk2Ob9i2+DgkhkWOd6cY8irBqdqxw123Fcw8paOoZe1okJ3XH6Adv2tOlnb3TNlc19QsPTOY0N
I1xPLkipHFweL5xy929wkQoYCiMp3SOGVLchbdcDp6ZLOdrN+HM9QBjYEEzLeVuq8/XFFr6yVITf
KQ0Tzqnc2znkXhjGV4MebUI0gMXHDPGON4iHouDrhRA8+ZW+SIvhys8V3sse2CGh99vyuXNW+log
YZL9wZkb9nKWJmhMNLdpVDh1cMNuatn4Cw5r/MGA79uCvTCLb9DmZZgN309u0I7oqIBRcXNdUnkI
zie33vHuBGqqR2RbQKVf5aXJUlgTL8EmhcIaVzEpbs91qTZRVxgxjuT74aMzrIYvAj79olJvSdq8
eHh0Wsnb1OUGzVUd2xiFBGvelBw91eYfsR7mHM9IOGVJ/SwXTzFkjEb+ly1Y5NgD/KJOkEfq12zP
AmKgvfrdS8Ue9NJTm5+Z9EM0r9OvXGdqRgsYI4uEEW14mK7R4MC26AoiXiiNJ6K45IjJELJs+vSW
yUGruFBIbpkjkk2oWZwlhSY4j1XbkqfBRYIqxW7/MG0+BzaxDwPN8lVo5xt1dtZxzU0ikNi+nYyv
8GM1DMpX+UOkvWl42Q565mFZOWnNsSF4IS7k72WUVg/dCEv8SaIp52Z6j6q08sFZZEwWfuKybR6I
szGnrW/HyiZ59vlgj/pWnmVf8KbH/0P0D6vpXt2KxLUaiR9E1g1iTnDdWRhoEgbbJHI1JCt2LqgJ
BUr9nO+s8cEytt7doU2F3scNxsgW99j2QotX7xxRJ0vGkzDLjFA1YmY3FQe6DtkIIMNKMHQ1e4VM
LUcytF7RXjFfLEDB26KLYrMA41BQNZRrW2b0ZnJfxiDH3NVEoMDK/3jvS9sblX399TNNAr6liUO0
n3ZxKKGnlHvJiQ5rr+2IFohYUavFqzLyfJ+qvOqqKpIT7Eag8Yu+Rr2DLO677lvFFYB80O5yp9L7
oOLc7yI2EIpNnSaR8dypirA1cI3/cQ1uyxBjgb1lqgGl3isXFPZ/ZaPAviiz/BelMmVqdOkuEhek
XoFmz0OaA3rmwmnJF6czd6wkdRzOGllQuQWs5fZBTI/rc50OGtHMWCRm2ayKAfqPcN8WBHtouwEo
YIfgMCyefmpPtyQxO9qUnffsPpk1Lb4P3WlJDEZ9u/v0XBvo+HalAZ4P1HQ3TSMjT/wD8ljdo+mE
WCK6a9aqXHj4ZQTVdGOVnKhRJOFBCreZ5oDn6Z2EJ+/5fSWgS3LY3wbgA3HFmlQPh2Inrdi+Ie30
bOpvTWyIvqIbg5LP2ZfbM2oUKYN8qcX8hnDq+mFBnZq7z1pYIFAxVLanpd4ZgVau2S7DY16v9g1a
sfkJSPxExsuNtKQf2CtRYRnPpXQGhSMTEpAQrfaQDw53AipRsiIc5OOMrDt+Zu4ReEU8HsKwKab1
MZbB2NFzD5hqmJ7tNX3uZ9b2Ywc2vb6TSQDx5RQTj36lewh3wAqhElLjJS/CypAYQqDCsxPa2mvW
WrLlmVhgEvVBIR99V+jFHhkLNXorOLJBZyVhMvom6FQEUdFW5sdqyWMJflEDD/M4qZVjcVKQpRi6
6vsTF5Up+chteDeQa/Js8AHP7jHOVJWp3T/WesVHqJzR2aNSuXyA0Pky2vGkjKWH6WDHmbsFVTJa
IiLmQdcy/J5HlAV9jYSxEOSrL8ZtB7PaECmqx+pcAnsLhGFB8f8u1H8LwsBDwXzqYqgpXo3sFZ9x
5/cXjZEHJMqIOBObCiT3YX0tLLl1V3elUX+YKliN39BE9eYb4q5FPdi48wCCT7em7wAHZ4WtdPXK
Ay7zMPbyeQXNXTZ/HdPqSa1XA0DJ9qGWGupYR+x8vpnplw4CnKxgKiIuo3YNbMqSrP5yCEtBnuw8
21ynenytzhaAsDzBha/ARCsI03/DksyRnFrqUmchD71Lb5wgux8oXAlqPSKkGdI2wHUWdM0aRj4l
q7A9HApuKvG5jxvodC/wflVU2fYDqHvM1qzXfCC0UizuMicNmqH4L35FQO8r+mSzKcV7otlS9bmD
g1xDPXo/eExw4V7DS5lDu/iTSW2GSj6rPacnKZHBQGQ9Tl2NtQWyWWSreicm0KWDiMSDdvd3K/hV
cpU1hp3P2HLikFx0dLawqls0YOnZrDWBVqbAXwsoFvweRAfvCXY7f9JGAUBOCE4JiOU5YQYtk7vO
Bl87eI/GxHSgXDcvE8a82UAfLAPdvQiwIXFt2uis39ysDGzxVT6EG8g1rKs9grwpn432k/Kj59bh
+ribzEXbWXp5BJnVlUxdB6Gl7pabeoEAJAIDQm4VeUjhSL4eLp8M7w/g9box2woFkf2R6JD7xyds
0FWeVJ1WlBwJf42mu41ZkmwBU+X+9qwXGoIMkSxuXhc39g9ZSDJq0pIffxrLKv1lrs8u4TggrHmT
yasNoBX9ERNgoWolR7ttp+MHeyEnu9VwsmHlxN5u/777f+iMZQV97XQnQzWfIlgDbhEKtJVAne7f
DuJqe3L6qxdY2tZ4XHt0sNeUYu0T89IDyLScYyZ1jm6MPmjp2wILB7mDiSq3ahlxZYO2AveWiHWy
pbLJY+Vk7DMfKLoLZYnM0fQNsi1XGPr0VxKuMQT1Q9Id5f3hX2xv+cYDFHFeHmLKaNdhpFdxCuhb
7Bz8G38tKobN1262OfoF/3d4jtnc2LCxTF4Of5Oy5as/+om7UfAfFv6Am9XMqR4kMQkVqMDxiku0
lLvuxO/4+0i+TorFCJh4sn3dqpC578uqXDgiV5NFM6yxvc4TpmGFh69LOS+X/+U0zUVbfaZu+JNm
VdjG2piBno4oxEScvFjVfGGC9UCP+xi73BDkbCRnLh0/49giXEToDiR8+7J1EN07PE9b57wjxv9G
2Egwr9Dh47HkNFqs1bfugaCBlURDuMvC0xB5EeEN9V6us6xMB2igLg7tJRobH/DLMOslinZ9ljpJ
53LMQFEI+CasonWX6+eELpfFGeQnF70j04Oy5bN1YTZvLAm1or58MSsRc/c2TzMyvAj2JoUiy3qi
z79yQ2bTIVvRYvxUGUIJi4nQhf8v6JmN4Z0NXmV7qZRp2RcCmNlIendpE7G7EcTdeGnqAFlIi5hO
LKb7hg6oVcz0gDVgOgoofsFQIUKwKsjVnvMbtyoYV2jsWElj2lR8Q8yMoo8DxJ87oNgNqOp1C5fH
owi/ZP9z+SRz7TlFrptbCXWSDYCVEkrgeUrkhqPaO0E4zZYOHTGP6hZMmi7gvfq2NziPyzEm/wLC
+OKtoyFR4WrU5Q0NbhT8+jjQDfCTifO4JTY9d0TZbARMOUIm6H92SuBjl9R3D7PffZqjfldjpt0H
dOJsDNGQPfGIHJwPgkMmCsyrEvM9JDkUyIxQqIraMvyh/cXnDjQjbaTHVPvF6rjHmNFAHzxYV2hg
v6Vv1kA9exSzHTTiZvx0CYfXXB7XoffeCjQRHSwdnXWcnv+eW2Bo3JHzqePxDdzMVdsXHBOHSnWV
1ouIRNq2EUWkzX2P0m0ilWkuEkem3AydMgUi8Qqir0GOwG6SK4fZwkgMvzITkyIIIxkAMrItp3dJ
EP+KT8hf9GX7SnemKZEaBNGtcfrkqgNYr9kJxGC6p2RMFqPeEKQ9iHHovjmtRtXAF999CjnfTIh2
Z8dbLivDLAZziVrBRq+UGonOSF7FyCWgmWPv4D9/YKqAuKYq0s6mtgUD77wV7rn46fZ9sRSyJGsA
M59TXCplQYWv6HZ1cvyym6yb6W/+LnnVFH8WJTLOO6XhqRSre82LcoDJQsfn0PDRq6uNG4e5OBig
VNokjTdPUwYICjUcBTNlzo3WSTxkXhcsCf4Ob/eEcBvkmUTs4rDPW7xWd1kFd47yurMzr+zUHR4E
Pj86JerwtbgJ3zaqNSpwVDPSVqPustd9qvZWWceMidpdfHQaJSZhOux6S5SHnlt2oe7se6o4TR4k
me85VX/azi3CktJBwJP8xa5tyGrXasv6bpRLQmyThjxFideNFWsKd0NKRAxTgLa/9jCGkIFB36eP
E7qhxl6bX8VHwmfTPuf+UrAEZvpMWmgPZ7335G5koD5tA2nvP9rmdawkEErPGBWoiA5O5a4F2fzY
Wg4Rt5b/PufTAgALj2CL/t7/MIXQtKw/eZNgS3T161lykyptyUZRub6ro0UepiyyTbPe01mRVg9P
2FIuqCVqbUhUSXnljsjl2b7IP9WCLcpGyAEViBK+xlxaJSIid2bTUol42DhxkzJRrWszrqvcMRCv
O5qdDLkUR5mLUqwcMiu8p51LiqmqQbuuxtuZEHqwFfMaO1/ZTXPCKe43G4d6/Oa8AdwiXjhNCPhB
jfLbYKrw+XE4jhbhVRRO7xTyZ1snBVcKPZn4PRCrKNDF0SnkgF1iK6R/br39uRmThmjbKRRgLVPw
a6mUKodUCmyeXu63SjgcNRICuIy9caljdWsYz6CO4NDoyHZxnH3Q5jKWt/OJVIYHKK7UVlIH6OjO
Qp73lK3oHRAFe2/zWMy1YC0agkZNAnpEyESgjfh0kjYedhWm6DWS8m2/5UosjxPdTl/R+0/Fe9NX
A+LOKINe+kOwX1edK/f0DFDG6XZs/d1HPgNVLrmCDfjulblQppGLWCItReEeb/4lvX4VhQeA92sm
jYxhom3PtjrymZmcL/TgTMRYujoG/x4AUxt8aTMDSq/sdXIvGiPJ6iB6UDgH3aVopAOy312WgrML
Pm0e2Zcnp2RV/jwgTxjIBc/RlYcdANz0YbUnksn0zZeq4Fyos6Mwc5I5UJMur8Xa8MPjqdkzcCJQ
uXQSWC8h1zjr/Qld9QUZfzapqZse+RIT/affe6XHb8UFAI/CpILUZ5U/phxe2WmMabWne0WvwTUa
hZm2Aj3PUE5d2lyjGBxVArShq3MsoU2gbIzTIJQgSkg7Qzs5bN0Hsio0JlWSaJQcxyiduk5rcnzr
vdrnayBLal1v8eo36jeF3wXRZyls/sf3hSEsJMvXxLVvRnlVEM0U/HWhujZeOIVv9ImPj2IOdx6W
LBheIeCyXYmqfNQep8zmu9dGKB64JUHs6868h69T5+WueNYTLuojxxuY4r6Z/s9WwYzUNDq2zmCD
I6ikdss41vddGaPhCi6Wwt5MRJ3E3eCxmBAIryHcKwAgssi5tE3aQIB6SJLv3ezz7r+ArwE/DhF4
nBFidEx1x1Nmw/c+mLri4JxYJRIFVURN6J1pP1HgBgZtFM3YgZgLgG3vMH5DfeNnUQurmf0eNkJD
pXgl3CM67pioG5Yidqaa6rfugQ/p4EbZzNjfUyecH5S3KahfeKresBOUD0LKp11wIptaBtpyDcv2
/1M1tPYjeLshZ+3Me6r73sXJuKwrdbrpfmqQ8tF6lXGxlV98GolxD9vtO7FIt8RyHWibrB2vqUc9
RPaeMNJRrYbh/eyYMVla6IQCPhjui6MFUH3lMSDmwXTUnmhQsfmObmzJBwk0icnXwWRnETWTdrYE
lB9/TTYSorNXRXESKLDk9qhjAJ3bOZAWcAE2kFRksiVS42yJp5R1O6HT3F4C1+rhsOaJEG3wGNni
QRbQlVCL7Oo+3flIwK+VwrwyQfcBuPK9zrvuctK2ra9wgvGT74Eq4VQDZ1ty36xUO7QnEmAze7Q/
9UWAmpXzCXcp/S/KZz614GrKmpRndbxDtVgl6AuWudqJRAQb2V9KkQVoDnsFgSvXEZRiucOA/1Iz
xCRHev/oYhCAJVL0l9T53H+0IRyUmU7ZX7rqEaPiOsEJnIizDJTZhKjAZH1sBfkGvQfkLafbvcIR
hXcaOENBZjjPYHa9VGTYPCDSmQdjRQ8R7puNsVTHFpDaxFVdRHqv8rPO7Qhawt92pU8i1Jwhxt2V
8BL8k1fHK7RLvvAnCMcac8nLJW0HRk5Hrv3KmLI42p0onH02T0zwsKopenn0z1DKWKfArRnKokXj
A+vmbGcVCPHwpLJEaDxtyilv5HX/HwAg4MTG6gvq5wTISqOMnOUl560AlYnLqwC3snI01cZ/9adQ
/SHQIW8OY6esBJC0MFpobK73KTyCeeGvT2KSrI8cbGknxBncAIjfnN3hXPXMuRtWzgOAHAGfCdpc
CzHvYmzAccv7T2XS+ZjRBmyMrcL2jzd4SYWlTVI35f3GoRxWewYTOLDqGcgLds77VuHhp2gpmUP5
ylxxf8C9bmJbqn/Mjxoeoge9hBVdeIduScZnB/XY1gia576IHEa1ezrtoqhdWxLdyTnLG4nwWTzd
GjfZ7ll6FjxBfeL1gO9hDHMxXutyAOiPBNElLLaRuIt/CjmkoqwLaXhlSJlOlrLs20TiVDCrXzBj
mjiB+iRFTaVDryHwwCLHsFc45ukmVxsEcnrXvYkAg4Ok7sEnbcuhh4fbPntX3RWemmDGO2rT4Avq
TlwUXv57+uWozQywDML4Z1MlnRHlCbJ5P3pK7G4sfiQ1rl21ihKNLOP0+676dn6K4u/fRgzxFii7
o5hz11gK3+JT6pXXBYPeYmxYI+6LLXTFYKkMnTPIKioQ6AbaViYg0TCdR2x3pHy3Ig7tzkcKkgqt
myruUIoQ1ouKiv1mbyAOtPhCviG6iyoXh7Aj+XAhXYwcgq5uaf2YvnSkB8YA0YlwbyKX2M4Z+9Yy
CNwoAXhDpR1beGAr3Ewhq5KyROyiSa4R9LR8dlbYTHWRxe7OJskKryyuRAENLyVdoghPaXn+Hiwf
wLZzEmwjdGTgtIHq9VrbOFfuuSgjcGZeYETqjtvYEyBLApTbT4P2kJ7vDO5RMD+pYz0WxZuFfy7K
M5rzPtO3BWXpP93qZd/HHf1YZzj+kEZ4C3Co+CvhYsadbTNo3Aq2x0ZMRAlT+8UJaMDPpO+4HpLw
VHtnyYPwc6BsotqH6q0fe2WJvLceZUSVmIPNesfEG1ttlXSsGxNM/M8SFT70ihdKGyF4jLmxkSDn
dHtaGvC90m/kwuqzlW/aTg4UrAGD0U2OzDe9cuVMjeXuxZV1aqLfPha2PsJgvLlBbQU38cKC3tvA
Xexee10bBgj+IN8Og5nm5hnd9KlVvmVZPULFviBzVgSaEmxrMbHOZSXciPe5eWpIk5vqD4+ws23F
O0EHJYXVqq7O6l6uS+LYORod/ab4BH8nhqynNj4QRrgxCeYUNPygPcL6r1eVN0Cfri/+TGH5tv+c
xgYyZRkajroRUedUESsqE1BQF2Hgjbbgzw+sDxrMwNMbhuQbfNW10VzknVB5OoytoDI0DrElHfo2
KC9NJQGuh9qs+RQPhvrybPLnssRi4yngoyWTea99H3sq8s5gYnTAkqutzj5VUZTLBC3FqTQMFjTv
/CpoU6DdB74dJvXjiFahOUUtuQW8I7xA3RqNVZfQ7x1PPh9Hj4eJqYtUj+OP9NfwtfdtXeb8sdLv
RL4etehKxMcwpbanNtUdQigGoxojb4dfltcuFfqIVWQZUaJSqr5Zm+FGR6Z5QKxSOUjEuoW5Tz5i
CADAUazJ7qSjM7wof0a3BjfMYDYE2M6vHVV4V5KP6STLjz8OBmxoU9DqVx4dKr1YE5qNHKCOLOM5
KqSVetMKbbp//kbaBHGfifzHEaumWNNiVTO59jNarkQMt61ZGhYTYGFVR9NU27nJ6rBhH/3yDeeE
deQh0yzv9+xlA8X3c3Xavm37IoDd1DqCTjmsLvOIkgHKxOr/0szlv6Zcj2lkasNBtWRx3JxPDuQZ
j2jpTnPrsUVwST1zI/rhvHetUkuy5ggzh8dhInJo+uASYBjb5htXawS1G1NA5XjYSM8aSXclfKtF
Xdqc41MFQHH7CQb+nn6jEStsGmwvJStWE3P7yWgUM3VwaLR8TjoCTme3SfbZxZIYaScZq0ftwM3C
o4ZeMeVY1Zy4PUYUZgZVclIv7sMU4kNJ8PbDpxGvTZ/OJ8xChAH6gB/W9qzyRXbxCuvQuVMBYL90
1E+ZAQTtOXlpxbZigJYQmD9AjEvfL52p63tECW4FdyElcmsyp6/ArDvA0HHTxLGL2BfgmhxboUhr
bd+uLtlKBumyx+/mH2bey/BsHJ3ZYpW0jZJMRLly1j5UX7J3XanOFdLRZUkFM0dVqYyEbnUUw0uc
7AIQvJAWSpS+DmMwxWGiD4Hecj4ZvhxTjznMEEzZDnei4FbTnJQYYFe9nXmJ3vxCQdijJU2YxEBn
TLuu61mItgg2QuUnoGwhSUBlZ/rpypkNVf6pPxvpJwcljuQhuG9tD1mzdrevkqxXaXCvX2wGA0Fk
YR/F+k6hqtwJI5zgmar408eYpo8LFW2nD4E7cP2hHB4bM8gXCsETSAKf4bJVlCKY6bbGNkfgBRGJ
VZOarX5ryRgwu6P0389cL+rw3395vK7zya+QcqZlGmvHI5Lo8bX1b6+5KwfEc7Ket4I2Kdb/4CCp
785xKZiCeoILqXzq59qazkgMoRFnN1b4zamNIVbaTox2UbWU17z3Z1YRyOI4aipaYqKjOgZrjg3/
FfXPixvrGBJpyjDiOVmV4TMw/UblH1z23Zibec4oPcc0fTUyqzsZSkZlk9X3pTW21TYepntsx7Fa
zUeCnNuHevWErMVpwm8lCq66fj9khbCFsM/zuwJURjJI7zz9ZXKzviTASRzmWqIe+iOY2b8MaTdt
KaHgypE5PJIM3yb0FAtlFpxOvCeTgfILJvz036RU/wBz8u8byswKo61qVBTkw1HShhrfZdUVaIIh
eCkOH1l2Bam9NTrQanm9jNutWvGTL9JbEOUZJ6Oz2S5oCUrvSupQPVV9Hv8Rb4Li0/sSUmLodHCx
BxZsZ20rBAyZYPrlQV/FrPzSQ1EFy1BYQpVE91W/ZwtCQtUD0tEFg/zzoOxKuEOihW2HEb8w8yJz
0Se9FpOQNByWjqysV3/b0zQwLkUuH+X+q/Cgzbl1xZHNEtgPNWwCQcOQOifXG4NM2TreEILoi3+5
voE9lIcP01fR4dgmWaD9sprk3OBW4TWbkNUT7D22jUQcgtbNgA1d4zDWgXBzIvNZTwqCuuRZ1P2G
bp4oHOZTLeZSgest0yKlRF1jHIL2MauWelJ8TfHreUrdYD/YF+g+3jJ3EwiNb/6qdKc7K0k7do1z
Xnw7NmTqIhYcfd5eV0BMiNaQI4eWyb7FCrcIkwNe5xWs6ay8SMbNkQHrMXF6qx8sXd6XmahsoMMv
adU1ITYiJ4tJsugiSMHL8pJQRGNV9xJGqmcoaCh9p06NjBoiVL5rrwfAYjMcUSGxam+zHgUp92FO
vK1Q/oVcTkhauRGoAa6YyA0+QLb/G2zshkqvYq6q/u16FwYKgM5feZsrXuPlubea4ngJQyCPSTlI
d4+BeYXo4vd4/OIwxKxjC3k9CxilAKvq+142ae4tg9u9aTe83ewQDZSvKC4y34UhmaX6fWoOch6+
HN3ryY5IVG6Me+1aLcNSqsyM40wPh/Lvwuldey3h+c+7vdiopbwClEI6bs5bFW0JCvQ+q9hnNhQq
vG69X6ZxcZmejLDyH/FiyleEf/HNcmNCtjKI3+vpaNg0EBdBlnoWD/e8UHDTWqdXQW21i/xGWAEU
RHwWsYJA7+2d+MyCkbf4atvoSNtHnjKiTDwOb2j85+0PMK6Eku3NI7BE/Lmn47C6FnX5JbC5S1Z/
zLbfkiEXrJVc4fuBaIhYeuUPI7A4KuOdtT9jsI2Bc4G78vBxyVrDu3sDQ4HtFPsRdFwFM69e5ZC/
8+StXAlM9rHJxvdQyhxHV4eegsQL19/xQVHRpqbUymMAbFBYlm1SSDCqPPyHcXxbL3PuZlEGAXr5
AJgSpaG+MqJX3ky94VauAL90tAgkvY9iAHAGEPhi+eXCBGMoqXUgJPpfuNyflAwHzdItT7/BTeV8
xNhvEyq+gGhT39ucMx4RSBwgLr8dRWEtOXwB5p3M9eFaOwZL5P15gZFC3cQ60ZUB6sD4QKiE/F+5
NuzGebxZXozyEzEAG8L0bgRQBN0er5UqgPjX6sC/njTuDsYQltk/qfr7n6L9luzNpiD4TOb9gce3
iPwdAuKqi3ko7wBCfHpmf7wGYc74Fz34w1nCLHg29xTZjHCdhPR5hB9hVO5pm5yzXPKHXzoU+Tuf
IwJ1RQVXgl4cqnlW/SFyF2RjmmkbS6j+/Pa9KGqQn8BynGZMzDVMN/pWLBGqfT4s8zKNa91yx3+p
m+vWVY9WBZ03sTOjqBFOsz62JS9/loRKPaqqiUYxBUaGcC8F2/L1ulAudah1R7rJDs1dG173pSoO
ccLtO8MJdAE5rwk7S6DNG5A6F7e9cclN6xNrhPjWSRX6GPylnL/A/zcWVH+Pn+NWOVU7XFET8FHI
gohduQ7KCk17KILrUwqwupZib8iROT34LmqajyZIdXyiMUfAS9+zT0XKn851h8xF7D1XMapJTGit
rGO8LsObU7d5JR+KaAXEP2Z20fKLMFcb0yzEuVb+Qd5BfnNGV0lTuKrpU8ksNdAOsows1rmR0iGw
K87DFQZW0e9eXkiaffiQtgm0COd08Rt3z/WKFpL5VM+xp0LxEyQPXYTWl25ik07V3XbExV4B4mr7
kjD40gdlCiYhwZhb0iCg6aWqR643J81+V7iJr33jvCrEPHEjEGfdq5eMfRXnDyXd9oVffNxWIQ6X
/ef2/c8GqFcPXnBYDxmhKtgZbfEykj/eVL92kqF8JZOkIisqzQv7vUVuT7eO9ZXv6+Bf3K+5ouDc
pJNbt0+zGRUPVxcd79It22LWONCHxuRCtUfjCQMNa15esCOpj3ddJIz7l2iL5xs3Htt5ADzyfO6E
9aa57VRx260sz2mYneSg7Nj4QV5bhEP+cf0O+uuxAugCwrCQ9OawEC2S2u1VSEgoyibIQFz3eEhp
cKGRUQx+ka1L3KNV1QZQsff5GJ4OIGNOOeZUC201XNGQdMDhjNR26o6t27iO6HrCYR6Yq4Ju/Dbp
cjT90iGymlLbSylDHLqEI8/CbT5Fn7bqTNugcme2YoE/CdZ9vsUbJfQjkGFmAfOA8fr6BX3q+Xww
nFz5e0738ggoKTuuWqHuJzLVGnHHiavnLDJ355xQTkltr3gk3wzkvItUNwpJDM/fTFGQFLKoE8+y
YJqeOCV0efKJvXK7VmiIc0zYsn+OVgZNisIyvjKD/WKkPg0C2sNkhnifQh64xLHVscyqk2BmJc/K
Ct50R84iV8bv1G2xRctfGsmvPSnklBz6zkps3PwCBS634YlJ0pi6PP5JnVSeFLlX5Akyme6jNdtb
66u1liAGlnR9RjAu/EFqeOmert+ptsx9ArWexLE0iAPvM0rO7RnV2gptYS8maRdDURLP2frXHVP0
Q8wZ5C3iG6xig9nkfo2KnujmkE7ZJfWtk12nB6E1pOvtaISh3hPnOf0d35tp206xLgWfUBEquexL
g5O1lKQnxyAVrAZuJ0i+5EzzbIB9Qvhu0n2lwb1AFgHv1jUQ/zi9uyV9UUSE5OSqcpz5005/3v08
KyNYYJAzsu/UX8Hg3NdhtZ+TANygk/ASSvYcgzo5Dyg4viIUoc1rxFEt3m1FepxD3RTIuJ0lsnB4
xotNnlXz9qcF1xqBy1deG6tq7ovJPAAmq3zgPK23NcJSfrMvnlnOZb0Iak7HcP4OJ6GehbThtrsd
lU/urh/0pL8NEA3Dv4c8f950TnzUXO5LcCEja0TCUT4MRC69Q9ympasXoV/KH3T7wguXs7CBpMoq
uZH0mNwe4o9nWnpo15IeR1kLnkoo4YaEnRrcE+ymQkb/8EvsySG6wHcP3mJOlQJn5h9LIyyF9Cab
+I2HUgzwdL99RC3yAr0LKi2bAfi7EUeN6INVfsG97LsVsP65fL42JGe/UaM6S4qM8F/MxJVloXBc
t9d4X5oDvZT+SUge+7bjSrDP/uUnz6dm2TUyQSAm40PdeViB/JkOHEsFy10t/8bqZZELajlZRSYN
6gM+gKja1/C/R+Un7j9r0aJk/kN1KgJrSG9DTnH7UTtTLzsaeYdi86kdYDPMb5yzi/WB7+T10vpn
jCDwOe0ygRdaQ3VTKkMXmzcf1Zh0SqqL25gS2hucc3nbZuPTZK/Ev6hNJXx0aVb3FENgI4Cx4aGy
skvlLbBr0ZId9qIW+zeU+UdIkP9eHl34GBEHY1MJDZ5gSxCYlGrilQdIfuQpDwm4GofOgW1oVErB
XThxS573074Y5Q96/NsFH8VqKcYR62z9U7r0uKp/6OCJvYJxI2Xoa5T7zHlKEPwP4clegxuV8Zl+
Pl6Y1Q==
`protect end_protected
