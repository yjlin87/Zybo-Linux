`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
pNxifUnZNyi27SDw754Z0NUEh/bEW/S28QnLF/lquIwFxRk/RAkEajhgHHClobA0ZjeKjbskuL9M
syCWY+Ui0w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
kWfW4MjXNl46BYRp0UiX+O3Q3o8Y2YfdB3qbHc/woZrhfrceZ+ViY5P5W+MbiY82kW/3Q8XT9phv
p1If8sGTvTeLJ5bKQwAQc3VG15wrTg93d2Elg/VnvGcdiDN5I5CV7lBHSjorVTxNf4qOgK31Fml0
QYtZiPAqHPb/K2x+Tpk=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QtaisdpSImUyyAvxxvPYaBFq25ACsqrIEq+lP4Q/sDpMmSUtx/TM/UBk3QRIyUQJ3GFIQxXarvm4
vrYPW6G9gaiwJq6sZhgBBrXunpZEeNTwvqkJGKkrRSyKOF1oVvMaFOgi5RnSreCj1QIc0ehcvwg7
pJqBHfuZRJP5suvgLpsSZMmqX73pmcSPQTJWMtRF737hyxXXF+Ty9X6USTWt22CJMbFXWbDtL7vS
aYVP/QZxh4JmZucArYUOrP4qhcRl+zY4birz2gLqG255mv1IpVb5hc1AaPHL+cOK1BLCfdYt4zkB
bNXvjD/vGu0LklilHfLT1o1X3/fz3qt2db8FIw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
2imtHlkgkECzMG2gtZFmFuU3GraMB1FrSI2cKfe8eE5slMq4pfjioeYDqR3TnuVqOirFS1aIvdmK
Eg7eNIi09YFS3zS2y8gee5W3QFgl4wCoZ3eKRgNHUDfL6fcs9ZTNTGcn/ZTMvTMkJcfPa88nK5fr
+GelZTMq+ZWXeF3gyj4=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I5u/QQ+B0FES1BQjrEFPKqF9t6jEoscLNrr9SQrELSfg/d2GJMFulJAY/5TSCpjvht86/ckxKcBp
+XhC5t4yLQMBv+f1lTYDsGKNQGr8c2QCBpI3lIZtjqkd2XEJETkKFI4KoK0qqUcRAiNgqLLmNaaz
FJAIFUKkmwynihRv5QIRXST/URXVsQBTCG0F/5BjfmywtGrtrTTuqyes+qFnReRn1JgxgGcNcY29
SrGgqhN/eemgjmZwEB22uR10s3gukELIiSxXyhggcT4k2Ij13ztuqGK2NxUFa2eJvne3sL67M4+j
uLIYTIVQjkgXJ+oEBZSk/qcisJa5eRgWdMKzDQ==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
czJ1wocSJ3lMyyRVofnzACuXtdf3DLO7SDt8VgCwV4h5JWuZrvVuRHN747HNuIoVEmrqJ//ce1HR
LhrgVM+l4zpqEDe18exS9n7JnxnJzBNyBytfcMBG44BUeZ6SpCniBg6aZqFi5HNgnhr2m+RS+t2D
8GN3MuBK1K7PcQ90dLlS//kSSd+rvcnKJs6rZ6BA/OA1AHCp7o+HYh/Pt+Mjtt+GW0ZhWxYdZ7Jx
V7W3V0VtejvEOWEeOeFznAdIm5cJ2IK8GvAEeAuUfj5h4SCbgv27C4uvZgQWdYNud3oHrUi4dwMr
Rp9uSiHzz0m+vFSTPeG49RB6Y7llHD4zM3acZQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 637968)
`protect data_block
38jMOHZkC+U3imE/Dm2JJYymr3t643kafZztrEl8hEcYe16SLHUOi+pwqy7gM16lLqnjJukaqbwS
exyGrVrmyvoa8BB5PXofdNpQjpmWBJ8pyIoO6okOD3u881E1iAUJIWH6jEYDdxksoObNjw8qveYq
bCiKdCDy9WhSI1nBL2H+XHfhd681iIFvsdWoLH182ayQF3ZPqcQsguQY1ZKktOtow5mwjlEkRY0G
a1lCyoJP7JlYsngt8UCOEEo6QuDR/vmEcCOfoCjWTG8aYsIXP7+96Cg9JrPStNCx5iO5ckKr8uig
oo4q0RJLksUgLij10ds9IlIUu5th+nV1ekJWnTHEdDPNJV/i/uU5kGiGIiOjtduq2meGiyxvrSJq
W+qepMhzqvQN3yB+Ozco0Wg7iY9NY9JL5iWXZNIo6RL0EfXdHgae0apwyY2p+ChrRLBqLphzakNo
Eqp1EaBpsS5nb6xbwQBMCtVa31zUA9iZB/qJNIcs3Da/0Z6ElcksbQ0jLMl2VLQFufyPAp4rR3dn
ED+QgtAHvePzO9crjmAVILKfGAm5bMLncgN15vNX01FC/Kq4tu2pIym0FRVOs3iJZAf/pbSl6Y6I
x9FbFdHXEzxmLkJ+SETi/fEK1Qeg6mlLPNWpIlTa1rV4ruvoTb4sLXs8MaZvuZrDxs+uAl8ZE1Ix
SrNoN8pHara8XCSTdJ0/WBWOVBId+xsiDSheu3Pt5XF/7icxmzx2ywHR6N45kNksvbB3Fy7m5+fM
6XB3tuT30owp8pA5RaiYdP/DBqbbWxie5tZR/mu0LYRn9LIN5oOEABNISIv953kfVhcpC2URtCA6
t+Tb14iIkAuHPZok752pIXMephf3plCFgMnJ4nplF78Br33cl97wX3oZ3RjdmcCrYTTKWyf5P6or
NBZ62B14K19T1ak9L5SyC5ecP6UpKR2/iQVMyEFnsXqWVNVJXcARr385gKMMnA8wXazq91t7n6VQ
9RI6ateGOL6pbJxKWwJKQjpxvuaJrRT8db2p8RTWq7K6zZ4sWEirowmgbjasYJFddZxWQop+4zSE
R64yV8V5GzVXaH5AsWP+9MeGt3kohRh9T1h0YrvEPpwZb7ftA3y/mfxd60OC8g1ysj/gcB1+GHSv
sOpx9fPDmLGT0D5Yh61P6DOcyj8F42b+lGeEbWsQI1UycblVtN1NxCYt97JwCJoJaMHhQZWQggpR
VqnsIMG7aesyH/Dd3ogQ3WdmiJlaSzTHC1pQuJsXgtyXKcQuwmj/Q/2M71Y2RT4KhhvHonI28dPv
DVmmgE0VDptBrxklv4BvzaBSrT5ctfc3ep1qpF1IYCV715HOog2CJGadPIK+hjBHjG8rTYmXzBHS
yUJxos+bVwYxUMHvmAsOScGsay/IKdP6LSg7g1HE1WKmIMpkdAiUMSWyT1cvUD/jkuS2HgC72UjT
MUM5iKbf2aRtLjlzAPVN3vmfitCAD/S+tTDYgxPowVhqA2WfltQGB2G6pJ87it5nNoV9EMBAn2Ls
fsVuGUiM+UEGNwp05RdNEJg2bhp++TcH1vfZ66yvqA7VuXciP+Z7LAShqvgX4jaoRgXnD8zi1yO3
PEnmruYgE5B+Bb+pJRTN2CJUlQRZcWUoD8x4Lcmn2lzq4YnOHhvZ2P1QvcuftvxyzuIxWXUHt6x5
K4C3Cm6QwUnWnknC6tPomvzEOW3OcYIlTqu5kSz3nzKyjkZ9dHqJEgTY4h33YshuI4A89/loxYAf
qRTn6i1R2RCwN1eP+vWWCIp1U/3W4wbBn98LRgQvF+WhElxMZaF3T6G2hj3f36cpi8f5zCY+0RK4
p5oc+Y+fCCIMpnhOiHF9ZIGBS5FY7u6uHx3ljXBpGiEYjXFwXVyfMHb2SD1Qz2fmjsys/d936H8n
JANXO8r4Ukg8rlD657YsRFN0u6YIzn368z5CvE5kFxQBWwFBCz3Ltjkv1xQXdeRKj9YgTGjg8Zze
11UvvlGi9ibHjV1Jx3KudjCwQdbVx0XRy/Q0iqF9/BJ3CObXPzrsxLPD79xCOLT3vsav8ceD0T0W
Vv1PCaf1HqgLM0AyxMOHTfO7mSLQJD7ziS4ZIRKEoY94+oBnLoS03ZZ5e6zrP2rEDrDinCusP4LY
S5lvQ/qa1NGZGCTOE1xcArrzbuH+kkwAoDY5bZPl7D3wLBAPcQst85RXCJ0DjJnKKG66CmfOLCxG
QYdB0IFdL8soZSRsq5CvhnofYfkOhI63FyDo6dn2FrBDoMpb052qCMF/M/hKk2WmUcrSZRRYvzhV
61LFe8k1WAcZUJbMZwizAAMmOcp8OILHAGonZ3qq8MbCZHN5KrPkzr/Yc7cUYe1/lMpViO/xch8a
xpfHl+ZPsFN2A6kvcjjvKtmOZkTsyezIiLd56DA0haRW7ZlAs9PT2wUW1E/icF1GUE8Tva24pkDc
vITtzDQZMFOOuhADpGvdayklW2F1f7iZc9i6rbdiRZKmazPKqWeiQioTEjQ55GJ+cGhe6LZs8/YD
1n9Jm/LyxP2DyIdVFsRowoeENSc4o89/NHqRmNk+5rOIE6VREBCpVXMQxZYvk89WfH5NrGJh+MG8
BSqszKPqQMquLsPXyFtEU22esG02FskrGm2CrVOdwM7mWmOPyYHrefTAx4W+tdLBUKxqIUcdDD5T
xFKU/a9yTeh0mrSDohzJWqhbkttDeBwky8LAWansKyqdV+ncfjJZQ8R7VPaTnEJ2T7qelR2SNSMD
eTqxRC5OrsgbncdPKT0AOgi09s5Op0lrQ/6FHJIhf7jdexRhUQuCxJumi8+JhoMGb35RkUqhpZZZ
5kgMIR/DZdEqV+g9kksVOEqInRJ9KbYNcnk7kgMuv6bBPWQU+JsYf+/K1BkQ/U92uXdl3FUbCXWM
uFb/LvhR6ub+3sOCqfCv8CSPAl7xKr1CN85CaiaRzmLeF9cLZ4X5apzj6WXgUSmuUkVNKCCl8QYy
2xsH+DQyaSC3kCS88dX5n8ypr4GGNbyVAiGtbNqJbkGuWdnKh4OfwlakUYuO88/SUyvXmLcwdrdf
ZVu99J0F88ehbtQztorisvykJcyOkNuPJu8M128ZK0jANsBZN3nEv3z31NoQFbuMcvDaAmWzb++P
8/cWQBn+jLDHan2owojYfmVKxJn0vuod44SSNTf63wsOCFNTirWUNr2cpfVzDxv3wuuHHeT9JmrC
iiLnZK5OulKIc4yBqpXpdSUpj1v23120gp3efVIdZpqki4d6RvB8jtDahSFq/Cmv2l7x9ZXNRsmK
HTvPcozYeat17Lhoulo5Il0UxaaGXBUdne6g1y8Nc/IvRY9P+FE6B+pAQI32v7lxJHdzlW7zqFUw
vjaOqWa3rBmAnBcBuIgq8BBL4Xs6JlSXEjgFDPejKtAk5+GqA+G9htBvHdoKQaC9sbXutahh7F1V
FJG49gj1ALiSKOryOGRUKPh1rTsPR6VDaYEduH40FjQXgjLxh0M+HFqGGRgigC9tAwTnDCYZMU/0
gcdDGw7cRa5XcGLh0MVaPWV5mEfeOuQDFftSLE6Kv6cD30ermiLAboqHRiOnnYo5vm/aluRmRUIC
fIvORZe7C73F4GebmG8X7bFgwYHdz0gc8jpXjr4d7yFWNodyVehOHAmSD+58a02bMjCJVYB32V5T
BDxSBQYDcA0uxxGHMEDrddFJ3mPOxVCq/6dqqnuR7YAnuynaMy8w9SngGMiaGs+BmeJ23CWi6osD
D4qRzoYry4Bb+hXRz7yc224XxsIGHR1YBwrBb3i9NJR85C9iCO+rkZISoPTbhd8loRCet2wls/z7
/jqu5ampKqnrY2AjEO58WcDF7ZUPhpyux7ihO2sfe4wRY2lFP7M2M+OowDXoJyejHYinj7fz3D7b
afJgJcSc5K7BIrhiYFFH5dPHEqQIaqntm7EkxQMVVrJVpto+KFjDLu+dz9NfqYoAFkB+1YI7Q7Hf
Mn4eTWdQG+EuYbODKrFwPE6o//TLJAuze2ngUomovLXWPiFRo0xTJhiCFi6/frAPNr2HpNP10jTs
vXubucw89baF1csNgk+hgWKu/Sm6NwLMOrw6ez+hltMnTsRJGyg3Cc9ad0nIr2yBdkvMRUxqpBBc
dHznI3s6k0elt1Y44EGTQPMAqb07kljGi0VBM9bvMWZw9ctKvwaOlOLID/NZs/Du3P+1lvYw/HCU
/ro1PSo7L0fzYEEC5Dley4JL89VfhYFQZ2ZHFxpCWNVc+v1WW1H3mlADaICPrg15T4IcvHpsWoec
+qY7N81jyu2qasWCC4LL0bhiKxLRXlk6ZiFBOFA1ixXPEno1IpjxRsDZOZowHZvL3NUM5zhjiCbi
6lC7eoe4lszIhULFFnRJ9BW2pgaUC/16GMc6u+2HzkwcJ73GiCEsD0Qsqi2YaQsStZ9FJ/mSuySo
seITuGaPhNiBDL1ju/4dLvkumtHTQZ4f+a/nqXYpbp+ZythNbV9RLuZx/88tSik/nkikj+67Pbbo
Ksasx9WQIDGCFbziuWvWEKntFdJCAy/xHGNtqmcYbMmVLZ4rbtNEtXHTEHsqQE5LLEJvuN3wRYMc
ovefeyih+bs8krzbE4zTwfg1Xg/Z0J6JWS4+VNX96hMq2PUvdB6BQqi9dJu0MmFmEhWgVgl1p28/
JGXMNFB3rSeIwwNAret8lHNHN93fsyoDPNbVTGWrTJMMQwQ0qJyChHG2mMSNvWV3+q9vwq6zwJcC
WIVa5o2YchL6B1GqgfdomXHD9hWxV39WpIItA+5kuJnQD90A5UD5Zq5mQVEZyPVrCxk1N3xa+zLv
TjQ7QjB//Tc8xi6UJ/uAkr/e2AkxQX9sDVcx9twG+HRKA0/45fOmrKtJy32aF+0FgP5BMQ936vgb
MiSz17Jy9jj75KA4fI2EjceBLQnW3VSDAspnpnGdhp3/GnAtVIgoLF9T+GBOQ54CD5E1wOJEjZwA
dbKrFr9sEd8R0JACDB8Pg62W4bPJqw1J28bPVrB3sfaPQOz9e7IAhW1IlBA6pDYgZMqxRC0kexVM
NHj9ZsMtVr/dWz7tKjn2OOgvismMzV4Z9GTi0RFcuaZe9nlc5+s1lhRVp7BDo3cs5OocX4xxBthz
FK8KVG7faQjwR1IwcpSjjzOlXzVKe15KJ5H/15hSFtkeaPopqlWX7BKzMoc91Lujwvucc9N+wyKE
rCf83H08JomfN4QpQ+vbUQd1ETh2QAjgSbrhFzFW4EwIWBkMEjnMoJi10Lh+j1Xko9ew4SEQvMki
ARmohvq9yvfdk579s9vL4T+rU/Q1yamCLQ0hT1VjrOINtKO/MQJkxTuWKi4/N9qpj8VzHbnfb7lx
66zX+6TztQgrhXRKYfLrVqpdgHHI3Onx5jjFwNfd02Ax44Iwob6IcAjjI5uQ8EEU0Yk8++M9Komc
e6hyUI4PB0C92U66lx2qty1vWWQsxJhgoUF3qLcFIQHxtZMPT2zctNYrRmKbM1JLt4H5jyKtgIwx
95319xIDW0i3U1zzTKZWSXIyWN1gLNb2/8M9e6XHSsJkwn0RD4jhHaORM+DMVJ58P1oRGshulaHt
Yt/sgh6XwOCO95ZZVde1PJ3H39RkX7orWAq5j4yd5ZVu6oFTLrI/5LZ28bup2Hahv3Exif2Rzkz7
Qtg3ys9pPJkffLuWTJZjC8pSCxEpYlDbLGW92Utaj9jueCEvVbCM/BUCvIyL15a/96sW6aH06x5U
aAVN9lO2PXAI7sJwRyN1R0g2AbDRZPph7XrCIeJon+Fg7+liKZnZmnBpfa2WQ3VCfkdYGrY4Q2aO
w5BkO686tbQUa4t9GBe1xane8Br17lOtqniXKm69t5Mz0cEQ4LGZFB+MGpbqUl7FjhQvUCwKVzYd
7IMBOHrV5roXYchBtPzuNNpXVSfdlqJAANxlKw+Nv2m81wATzH7UuuwIe/YCTc4SBqfshJikq/x5
Mbl9/CrolDe80+qKrPhoDhnItMb7q9N5w6ZKVeDLaJbGP1OJGSk5uRTdXSnxM1aFUMW8Fjsv2FiU
tmfoS8ekneqgNSA8oNJKLDM8mnMmPoxxDIyNRLQMo9kTkd7zxXcSDEecu7EuWfKEMTKb/6WoIdTw
x7V/nVdK5ZdUaAJ4gOjqpQgbDp10Jeg3dJumrq8QYNR6NkAQL6kxvc1miKHdmGTucSFuGbgFmKzg
su06eEjDTev9P/DeWdYa5WD/SIMhsOWB0cKPAWnP2nOeQfxFUM9e6bdOxMTuuzK1DGD2zBlR83XR
dohSRaKG00p/+0MDE4RKumgkhynolm8apItkKjVpEJBSu8XGxWd/dV6qv4diMhprI402IbZ1irRe
lr+m5MG7DfNvtyvxqJv2DZ6d65ArnOHBtu3Iu8lNRwvRWBVOMGc0Em30DwRDCDnofSTNXVAay60n
ll+toVOEWJn+OmhLJZ2GiWrKzHikIkWdnie0C+KcGOxxuL/WoCC78GlcPzIBDFnUyqYVZUESYhsz
Ydw0dAlknV91UASReU4Pf8SmTYmaE2wlN2DM9KeNUBLfkpk7pR3COLMQqEey6g7ueTq9ElIBBUpl
arfJnlX73pt0LuI043nrZGOf7wnaE7/joCmVTXwoeLJKmpJ0oBfrwElGNkDgvmehZMkW72dLe/SE
DMRsLmpB8Lww8sV0xOe6zcgmaaDGbizE1QKZvNc1PTo2Iqk+S/mt0q+8jbPhtxjXyurAC5pk4gS2
7eO2EhbDfXv0S9KnED8u4RA3jvhr3xSr06GV363UjEdwPsmJYZhAV6pdVi9Gy4gcfqD8hFoK3VB3
kllUR0KprLACLHBcGcAVzmZ8g0AhqDDdQBXUuNK/EknMQdXg5WEpdBpXWxMqBIV2lqBU1hm0jkec
gQckx/4EMj+MdmE2nnAkL8EhaitbS7aZs38S6h6+jQPx6ERUesNC8GGwuq/77hkQqzGbqbg/Eg3q
YQrivTf9ww8zz0dyn1crS3u8FrEekR1XjlqHuB0gqPUlLMSLWCGsdaueHYIZ7RUJxdCotuthLStU
dltxHSzS20Dn8Pfuy41qdP4tNPBQycWAeHRUepPGt5nVckb/sTLd14/WCVn5xksOnWk0/y+f1WCi
K9qUw2XZlU+XfdljcYJYyfsrEfBXI4XScRpMi1z3IrTGLp754eMTbsWcdLPY73+sSpAkmiPsiSMB
cXrcwqNYSGywtFCNeOb3obc8FiRX7LOyW2Q+NaypEgeygy3lifZ0At4MwZYyrIDBEzliM5cEgYTX
wyTearKEutgc1PrPUBq+g9L3zyhLzgVZimdjAuuCKX5IefcTfwxYO7+sj56BRArujrRg0Wvls3ya
O0FGHH5PYbO4i/6cHyWHnTtNROpLYmgyyhK1CtNjPKQw5YNFMyKpoTDTT1qSk/qZrK7TH9DtLuGc
TnzQdHqiFw8r1uyVWwsLMnBWQrTbE00r96qBtZqpNIEWaBbrPEJjCFI4IIPMljjgdzdbYr7o02TD
mTDuFBRqFKq0BZIPq/zIl5LxSPTmeaoY+OnpZn3/t5En48cvKAKYuvlGy1avjtQioCVRAO6acNm7
B/l5BIljwCVqAjFE1sOlLtIKxPXAwRkYsmCcBOK7cyCcmvTzXiqzsrXVUYdU3s/eINTvGXBUz8qx
+fjy/SwI2LjhIJDaWdCihSHwgFvcFnRHsDIUSAKG9UwJIHHA+9Oscax3yjRPv7weFcM8R3kMhn63
WPrqbpKLlMCbOR0ILzSyDO6UHYUyB9a+1EA7G9HAJRYg7r7SLfz1ktKHocL9/DPu62J4NSmCLr4G
oMSFB4ZNqhk65Ef6fCMBMCTiCexdJDyIYBjLlSKRCBXuMXBYtapY+Mz7K2KqpFMTulzO7afjdpUx
Eb47dV079k1Z7KrIaa4SwHDL0kWO41Yqz6dFnSuGHCBTIUqSaJm01BBLbxf3pIeG85MwcX6wAuKl
P0mFCPg0md85oJKbo6i4hXzGFrjXttFh3uuNygK03XdKN9jEjHh4BQCB/bfwpqvJve7bb3NoYGye
om0wosigPB2DmSgzvMVB6X0Ea3i538kxRDnZGvGRBIZGbFjTxHHEcqf0PjaEqfpfrdHpektzvOc3
aN/esTfs1yWou988Pia1An9/eUrW6o8l/U6oWfwrXl89OJmHe8AbdKY+QXghFQrMrDvmADj2YXNn
ORdmW1uolA5Asx+Xwz0sTJq/uBIMZ5Ooqv7kgwssVc3HOFoDFQ0JyuNC1sxByntHiHP1T0AlG6b6
9+isfCTHP0IUpuieajM4BQPRbI+DHUYKtpElz6uMEsaLNeGoubkCQ5dDouUNs9Z+jqjPqWedSBvN
8kx/de7H9mwQMIGhdGh2/G5ZFpQ4rnx3XGLV3GXEOOG54wRxXg8WYY1N17Q4IfSdT3Z+q0yl1boB
qQTa2Q0+BFx5TvkTM++MbCMpi/Ye92OTfAnNG9iXREoV3eaE5pPC3vJBKaiIrXahpZk+WKfhgMYg
C9BNzYPCieZ9Onp2nImQnCHvlwpY1cr3MFQPlVOJmKpGscLPPDZPqR6hk9H9JFZn0bcDMQy9pOWr
recsGxfW/Bd/fILNhNgbAYilToA4nJnHRPrrUz6qeOfRoWrinWFl8cLSsEC1aF+GC48WgLh/qGQg
QufXEE/VEt1tqNh7IdQJq5eCTaZVSL72iX0RUxcmT2B7DcTphydZZWCBQa9YpyqvQeQ850iScAsN
zhiY+Mq8LcSLzxtB/EaG1VLHcV+gnOciWPUtLPHGnZ7QrSSZuz4btKt0N/tmnDebnI/sXQ1Zl9ol
rI7YM16WnMF/oRIfX75qLObgyhj00XKh7a8Zzihq7JBXxoNo3sDsb5mdM3BFiP8PdxraJb3B6paX
qhsnXLf+QGS/IFcKK9LA+w76TkJ0aNUKIqu+L+7FG4ERG2QdNxdQtJ2M3VoILxMCimCYMvG23JsZ
QOFDzLmpwVuVSLHhWxUBoikZhXg8be0TOFmnf5XiZ97sCwuXF5F5sXU6FFos8TC2dRUr0mxwPTB6
QUg84fL0nY5kjivSqpoFfjkGr3Vm4EWZBi7R0zMMn2RjdLoEPNlp3n/2ERaD7I2vXSMzHwOv3kJP
eudnV0FKyeGgOiHhZ1z0HzZ0QiBc586RaCt7PI/f0rVLvKRJ4n6rOntlY56uQ/M5H4CbVrfHeWGf
pjrLGpSzk+zM9TleVbwf+mzcGZXFihT5+wf6EV/B+yXuqNcBKC7lAO1yYvED0mtS3CIGbX1BENxm
O0aSmVwlHhtu1IPegMQNzsVtG3R2UK38hWFYjQMXaciRt4DphKlXZYxmHKoOlviHdlD5g5KY+rss
8GK6FVpqzdbL0hSwHgzbnKeej793T56xDgQvXqeOUS4Rhn8LSrdW9sIAtYTDJqlVkDr/a7y5wPL5
I3Z9LWN+QGxt8n9uabqOC4Um3GtCIqao/U0CdKcSlQKUadZeTtiVyg4D97qBpUiM1KbWwVOk2HBu
j6V0QbmoxDMvduBzvcOrW/csNB+TFgNEemuTRI+bm55SDlzBNG7xQvq2ta6U459tlziqbSxIcRZz
SCKcQWWX89+wzS7rle3vvBql1DVMuhx0jvWKxCWGh/BzWN1bZqELdksSDJ9HAPh8DPMjdmV0YelC
3XZNuTJLmBQ6iY4IkXzFN4mt3HrtE8yi535/cCyPVzkQkOcOKlQ/c4ZbIMKh3d5AmFEsJmW4vg+p
h2uk4jhKqYJkUdB7sMYAOMlPRMEASBmFtAKqQ9uG6Jmwwls/P/tz5mID1e6nxDHSDDFgLYYwxbMS
Poemia2sLRWHaT5DYxcB3VoNuxvWC87B0D1PohuohEWmqOc81dFxtwwO2KfMXBJpLGZS79nmc/Vt
RJ2CaBq8zPvTifYSmLcGcXqZntnhLmWFsAh97fX9BRtSm3rYbxoaIk1hnhLaOS1QbDfE65thDEkC
XlJtH1AsmIwUt6jIGpq69G4TalP4DEGyMcyklkp3wWNFF76WjjA7WPp+EnVoIq0gKMZKBYMvBB2O
QpsnasJe+GaTX9V+upS5vFfVdsq5B91IQO8Ln5EQfkPcQeeVAloKIFoRBUi1kuUy/aor50Oyu/QH
H3Ej3CPWzqu7rpQcEkOWIbY3QQ82Dj2VdrhvmWZv3DewSaveW8q/htDyUy5whfJT4KOFqM+1Rx0O
1p+vgzMy0WvqTlpP0GADpSc44yXtf8LPmlShtKMlrpUiSJ0BC4FeeQ/orhxeakusBIKvoH8DQYKu
N9n/E7xoOz3hEEG82M7NxoKcyrH2DMbQUcaGVU9MvrMZqHAGY8guIXmtS7i4AqMZB3tVB1/MusMV
S8d9440BGFchhxXCKda78SHFx/Whg//R2c3QDEYcEGZSUNniAUKTejuV/8x3gVr+7eA8Io3WiecZ
FLBSqZ+yX1jQUhigyQSAwKI38rwCnZYy/rztsXu88nBxHq8rcBH4ln9lS2SKpl30cAG6w/4haLMY
OA7flt6FK13uC5r4HNz+BtqmkOTtsCIJ5b991wSilw/l3SPWaHrctQta70K8E3l1kCZLPYfoTlEH
7UeowxLwRH4qUFH+Qe/0/n8CTYV56ysPi4m3/zZKsnsNrPV9/8uq4TTaNlay6w3yHn09mNCwAdvW
vLJaA4bm/W/3gcioDxb1HkB6lnADlH0zTyPBdiSR2ccEp437fmiYPhjODowk8BhXwGv/Vctnr9Ng
PBln0ah99OllHSfpvnNDmGlBQofnxNg6d49I8TTVXkAHSYPUG8yAbP++CUXlzVjgd5URNCDtXXPY
TIZ8J4BbLJ84xBWlWDLq9mRnC0jpUYRIcdAj90/13PkaeN3tfg3COAUbqj7VbU5ppU5qmnZrYazW
mib7+rFC5TrAuHqX8K1YKOz9mlHsMubGNqs4kbOxcwJYa8E1AXR2gSWQ+vvISD55U0bAG9qpod2D
TbVapup9MlpfkLMKxNXhq4OlP1jl1U9DeoDqT7rBhbxqv55XVdfSrjvL1jtLrVPu6XacsrTViv6O
5Nj2s1LT+pqXeW8CVTYWrRh6ykNUvkBQIOsyaMqqBcAGGc/nPs6VS4eiYdPZNKJzeUTJV0wa6FXu
hYHZF3ZnuQ56mXUz98g/MOaR+7SU3KWDyZia4U2vsFPVAUO640z0oAq2iG1zr201SQJgMdSz26+K
DbjY8lqFGRFZudtN726Iluqn7QBOC6uxBYCDBO+/++hrvlTy8MEVz7UtwRwueqnKGZVtnsIYXZ3d
NAGdWC1ZJgHVPIrOiS9YJ0ygB/HYL4GcOSiCcsAAxafTc1+05pogSpofDJ5sJU1fmrXGBwfk5lna
X5///NLUrafPmed5MBOgyyF7oRCCh6fBK6ZAMxDmb3rPbyom8xcr4RO1u2SFNKOInGRlvScpSlVb
CwBzl5A4w8/VeeHy3Ywx9kiT7bEiYf3K8aL4gFlGcdAq9RudEELY0QfDx50VHg263kGSkzPbPttc
r7T0lTrofEVluSJLqVDP6JvysZabRFg+CKKGJ3uUNnuh0FegLMENJjVeTsSvOoZTEHPXuNMIonfh
c/6yGCqtu2uhHPZjeM+Ddl896TUvZgwq6HFC9S8JIAOeQGNQnJFE9+n68hDOkB3xxgbBHJk/Wzt8
85YIq03DRuGt8HlUAa4BzUrEzLffP9a6ob/Pq4kf2gb9JPfikqgw900WyvxLgaDTO8HrPz+8sd3d
skAuX3AnAe0Sd26x/Vx2n2z4ce3Nb236h+it7dwwBRwWZOoMmK4PaJtRIgkz1O2GueDmaQeKRwX3
z8pbfbDLZOiDroo22FYGEeh6anBeMTVCF8dHflnDZHtMURxeZ8kBfVESWZ4yyK35L6t4Zy6YHXlJ
OKR0Q38r2RS2xSZIlo+WivWxvsBoBS3I8PJfyhlo+PhQloCzOetG7oU1uuZZxP0YR9sBHmG/9z2n
agObt9E/TnfuAqRkDjASZNhYpvzFrsSxA3mCA/xaYKuDkl62g4nRuOgrMoxkW3DSjrk0fohqb7PE
sTUOjiz71r1dW/VoncSyAtSolAK9/RsDalllhw0MUwr9BHiQg0SvTDBx4HIWHmShrNpAEVAaJy+X
Na60M+JvVL38GdlBMpiJmxi00i1bSyUH/O31jK9bbZ1TZDvAGhrNIw4rt0+2FKmlO+9wJ0WWTAWn
9h6w1IE2CyHIjym8JyavYXSq26QqNaqMW7NMjVPfxpXxQy7Trsin4OwNxjmJQviNFD3ZbziHnF6+
pHFKqqs/ie90VvAQXwyCZMshxdhS8FVlP3GqXtAofP0wnkvRrHaYAOYr4Yu+5PwvuMkluUf8NU5B
DcfWl/Gl7V93NW4slYTbwkIwrXPyV2bR8+fCXpKX/OdKwfOy6EAnRGSyOdyAB0DROtRdeOcj5nur
QVZdxWzAlIexUwLQT+BYyLv2JEuITmnU8QJ5JsXng/Q51ypwRRHhpyvJzcRY3BkA+xNVen6Jvz1C
F0CTdw0GSAjn+iat4TSD5+9Ny5eefEJtxMg5wR50X3647gpmAHq8gUNVcnA+xiTwkfbdjmLPXDaT
CsFrbaaobP4vRUNF3PylF8QXKtQ54aoSjPUFSsU4O5lT+nriHkaRyAzJILndq44rnKRiXPYvGt06
Q8OmRr+CkjNlDyIqUZt0ywo7+3469n1wigekpWizoASOkWbD7s/JpQJPs17+weZvqKn1I9MJEUDl
BPscJnqt9SAiSqEblBSR+nuFBtwY6WR8xxuP1VBhqVu+qQ0DCBHdAgMN6HrGpYqVUFRUsjCLZ/72
r2ptiQqUBRNaz3bpAXbtuwGgsdB15egHXFckfWa6m/HfjJfVEtw7asiHC8s+VPrDWt2S0ItPBVEf
RuvuZTvOgwtKhiFpY8YNhXqPU//QznPXi6UEDdYGdWXGAfABal7bMhg3wT/qu+aUQImbwKFRmR7z
alp1pZwIDJ3ledTFTsnxbp/o0TNmvmPygKDakyC+NTxRnaOf6ZQm/878J1WSHpjDDYhC2LZ7dMI5
4pubyGAODR4PpoVHOLXt6vmMPwI9wI7PCMai7NuwD2d0A86ZuhTpSfKnquFV0r2WI6nXhz9z5Xyf
mui7IkPMMwc5KUaVabG45XljO2MH1+Hnd264vShekBg/3WKIhImgRDkzrf/NOv6leAPB7vNgNwav
GkTttleCcMfID7b3ig3no6rGekiD+92y0pO603Mrh6udAK+qU4Vx9+V/UDoeKpFi2A/rwL/NQhQD
13avOm9BgnZAYrpAlkcOlDmQJdVSkJB5xDSAFYcV6IjVV/IYwypULfVpzBsQPixUnYU+S7Upbw1C
lsYLNfi2oHuuxLY86qRwFAKy2FaUTUwyBAmW3l5oShWS3PawyAHtcSdJ87KQPcf695fecX7yGhgy
V0RT6dSOsY1KA90yoPsl4nEd6VKYE2sjXLgoVuqYLexQ6IwubDMaV0OhZ8jV+lAMEoWYlYBgQ5qP
sCczyK+EOPQP0mxhF5nkjEWDftXt4B0k8tcwzCenB7LQlcuaszkPkjnDUFpMTOCMYwO/B8gCuzg6
amRfn2VyZLAt1NJFYguSMG6alpDScmlbJNiixNG7Bch9u1TTG6ai1Hm4RC0/pq46K4rhwfoWXulz
S85VY7cQrB23zpi+d+u/8mAX3Aj19vPZr51Bi3F7VEoVYD65CCISmakkW/cZtHjCw6gr8Ko9++Uq
P9swlFpAHejMnXglc+tNAe9GP4ClTSbobwlCYVeHAuEMEr7NNkGnXb+cum5HVK8CMfzGFzrPDV1a
6j48bkeyqR8PfooSeaTjPfN86NPOXyR9TFKJtSckCanfaKSgNTFtCLrwq+n3mvMYVoamSls3Gso6
pC09SBUDPEftG7e6u+0OwUMx8XwTXNWpBCqodTpP89Ut4ITKcAmyUyoVhG/jTJIejyLyGLikZ32O
+yC4+KNUofDnTPtsyEm0/rnofuHeKewYYjo5VzIlkxzRe8NLXwTFzug9hTI3XBMdY6x8e+c6uGh3
4OH5Nh4s6xTY5mjxM3qEztakZ84vKzh8Y9DGId5XZVCfz70CVh9sg3AaFQx2CoSqPJ93oE1tF9Mx
XxaJojZe5T+QD2ZqbBjPs9512UTZxr8dIKkX7dR7Ij5gy9HrC5rk4G9N4UgWY/TC6C+j3w1nQG7n
N7TbjyvbVXw8hyNm/fSpIrfhqTXA+aNb9+/IdwaIW6idDbUGOseijj7S72EssBDv1VfjN8gLAa4o
48dg8z2jfRlOqOv+BdRQwKGWN/9C+asRHrEg5yc/jgJ6R7LwHupJABxMaxLjZ16yIi7zyDjYyxk6
t1cTCmonm5I2hJdxdbgdK4si7c0CansEAm8/1/62Qz6xnhsOElrt9s45zFmL9jlz68ZPgykQMqKY
1KY7LKswZXIEc764GaVfaEO8wh3mrVAr8Dwb5ByX+ipnfA5VvD0zWFSwHLkyN1GVTvZg1mdYhDcL
+08/E1j3BEIJVCfl0q6tKmSkU7L0jrR0xEpSCPyZfK33hVMQhztjKzAb0oKi5M5PshhvTnh1pCQh
tIppAKgQKsoymQxXr2/xWxlsl1CaNN64ITPHu7A31PUSkTNjeiqjjttJPyimbTKAh9H6AbM0d5RC
DQXunKAl7RMjwPVMjpEiaDy6pA9Dq8zb276AW0RpSdeQ2F3Y4sqqYiBukEJLsjbNg2A8F1ys7e6L
T/F06oo9mLrLTzVDeQBIMJJ8SBux6qjkzY4JKjzsLkgtZ5xMK9+mYkK9pv72IyVkNb8+m0ymT1by
09AD+wGhdbH5Mlhxi0lmlNouz1hJAU8OS1Wq53wCPR+nllMNDX+xVFPHWl3fIehcqzkG/j91wr6H
0Hu8PW50H4SpiYiZxB6/IBMfN0GzPARb+3NIAnrQ7HLJvk0aKszRioQUQf2On85Y6baQlj3ZoGNc
kF+LTGasHQvAxpJRlsa2+XZlIFUijUda72ZkDDUvebK+OuWGQ562PlXIJ+XCOBgr07UBsyDgS/vP
1aF9iJSvuUYOQu7EVLZ/wnbPtrstJZoQlfmRLbMut/okQrkK8iHgOCmHNtRn3EBk+q4Kof5ffcOB
9t5flg0BxY4d4tdryWhe9ys98K9B8HWW8pE5h7pbFExL/ESrXMf5WZIgYr97/6PD6X900/9JkqBi
IS0wL5BzvfPA5VneR2OQyeogitdjwc87C1+kj82lcQp4iyDf5AO7481PJygN+kl+Z0OaXpIxdT24
+S7kSknAsrBcuPuEScH4RkBEe38txPen5gTf2d1sKjfcOUMMyyCvIFz5ua/AiwTykmAhKBpg5TwS
QIGuhkPRdl3ijLydIK8w9knSVFpYr7GMSv4R5I+I2ELT8IOaxx/OZFa9qM5tOHjIyWrkbO74tIXd
8TN3o7CWZ5ZqQXRC+1tHm9VOFP6aIcmuoGRP8zVvnJHdh5sNREVSs/DDfQlMp2+1jxrLuVsoEMdv
eXzktToxj2CT5oj4rGCJJFUkamd9vRORDB7Nk6YoLSMeh7ZXAgTFYy9WgLTrN9dOA47tGn55Bm3G
hLYe2P3+1lpCgbRbEufku1Ar63oLBUNDjPSLyYxdWd9LYZ+ylh60Haljo+wPy8yXhLxN1cwxKqUC
VNWkPCzUDr08Qcr1y/0QAfAXDhDGbH2LVFYzl0inpAG6NLEZtbyrzI9xOigfSlPG53Ihl0pQzMxG
DoL7XIYggT+x7BjwuMdC3uVR7IlKYeRvPMVifK7QNVO2NrLpqHw/iTBJFjtiaXcSv5EBIglyOufN
Qx46fMmy5nU59hHyR7FghOUhsMv+ErNZbq3WNIuAcSi4QFI1k/woHif0YNIOmjcTZbIA6+lM2Nfu
9GODYyt5ma7b+Bn8bO54JMtED81vnmvBZxr5iTKTP5u0D5pwkwNMIfyFOXm2444QLmVoTYUyO5Zy
7eTx1mKl5aOw33upfI1FwfUnhnccERKBStsM3Pl5+N6lWdvTyLGcTesekc+pvBy5Dq5nMY9o9JKK
koTExxq/CzXTRJzIep6XJnmSV7eB365u/RWkjqs/oWwQm929k7QshfPkW0+lt7Bev92oz6U/HO5f
o/XYDSQ3wGQONOtEmGyr+kWv2wQS4JidmKuJJihyvwp2lHEdd6MdiL7AudIxAnO0nKXYf7ezl0jy
BANui9DQ61dziPo7Wo5rKGE/eWYtbWiSamprC9pqSD9gyrQPkN7sn+qUPvn7mVhuKC5pbdDv1VkG
XNbqGPKF+n19VMEdDhsHXJnsQ9a6HwVbowWHXMFW3+eMLXuZ25ubCpbH20pumNlM5SqBuFf0Di66
YmKNyHu3etP5vaawnoXvHNVI1ZtF1gs4Td0AfvaF91hN0N9Tn7uNUM/lvsOjKRRGInnA32dH3yzH
PI7xgNbUPLMWAvyH5YJUL3/+Gb7a0iIQBy5DVSiJuAISongl2HDcRTxu7QvMBu0SCkXSHNkBvoRC
OEsLwg+HH8xmjMlMyJIcysxlzG7FRoeI5XGnrztw/HmzfydrA0ldGxg87HGZylFDa+mEkxXu8PWl
5/VgOhThhSUN2cHECu3Ksx+zbiRp1yfKZuhfWJv7XRdZ/sShry8rOSn9t18CaytVmo/Nn6fdAJ/r
sWXixAXsd64WxqsIw6LEBg+mKdmhSCNwJPeZaHnQN0roO6ACo84zqZBXmiot3obQzFWs20lTmupB
OEsLHp38gRL8ZmkRjoQRlMeyts10kKdSKl/tm0acylrBlOqPY3iwCDViXmIocAkdYDFVWT3J6usF
pk4DP28rRVjpwMWmaS0Ye5fguzRcuLfY/3Fgnz6pUTQzTmdotP5acojqZmU/oVn70h9Y6oOmDVKs
4PGdRp2j2FmcN2UX9WuFLScvc0GFaWlyYAQZBJdBEhcBkxrxgHtP2EpIvxdmMVotSOsq259i2jS6
DqKEW/OImknv+dtlJl+maFNAjnRQdqdBEr7GIU03UDxx6jQlpK0/2/4Z0KCgImgHuDFCJqQque2k
S+h11BsAV8tw3XiA7OSbYhZoVrHiN2P//JXmergiHUKY9FdRudOc2ySOLSrbV5EVE1TN4AzlJbsX
hKoy0KY6bmSi8B5BFInRcV4mFpNc2pL37k58BzM1uS54NDukhcEz0J2SSvVD5t4G9Ha5+jikNNMk
7hFGj7uwpduFcjOo/YFD+NTzECL0wbM9L2+3PYNOnTD4ayPBuZ1rnmIR7Nza08ZRIxPvzQXLhjZs
BdxS192t7t9UqGLR51czp11dElSF/onv60baaQBkH1jz8HG8SR18Kmh1u+j6y9Lh7olhJ3DHuhCy
PX50kJUsRp5/BClUlMeVOxp5nj24lNDET3Xij6EkDWKqv2Q7wTDXhX6sSdE3JR6zw+L7KmBSEWFi
zsydOBGj9J9N4sriSB3ZcC2aB9j7/Cp9jOL+DhOy4CwM6q0s4fFB3axpml7r5UxS4PnhsxVerDfj
Q78gxACpeMRjkmrty2c9U0Z7N+htmuSEwj+4VKhjGMY/vbp7N1t4Hz03kQ421poy3ZsgCP9N9B/C
8rQ8glWQEJyg8gbHSbNJlrkEqsJS09GW5MtVEcSy4wZMDy3+SPp1Vj4BDPFou+1piy9PtVvpM5id
UDWJhry7gmhxQAxruhGX8TTKD5pem+CCb5mdrMv8XvChxzxa8GPgiLQSfMmMJ0eW1eqX/B1I2omx
AimLD5rDMCilfpS/qW0dVEfiGNTksyJg8Z7DehVve7/8cN0BoXN1z+X7XVY55/5owCweFrSz63lf
2HiWGHG+6RK4Xlr2vdYopj7rv6JbJc0bsTamB4qcSQLjpR004EJctequhstTwMmzDEv8YPBhCdxQ
g7rhjDGce+8E4XkLDF6z++vQ6ugAXa4lhN+kNblxjv3Pt+lNAaI3zkxlAhVkZfwDUg3ruNw0eOkh
+8KOzeRR0wtFA0crKKjcOMo0nOaI/7F0fFfD8p10lGWwhBvqo5SNxxiV49JNsmv06pAoyrWdSAbI
jl+RPXchnnA3bBtdixo3kPZySzAgNB3O6FW7Ytbyilm4XN4FkN5M5YO852y6f/sWsMMQ52tuottc
qJ/RDfeiLdgMYzlJdftwsnj+qNI6d043z49ERBMna5xmO1enP7th6eYx+aRQKLn/2nnw3QNgtwI/
gT8a5qHGpt9sWPQ5Dw9BFO3bObgZiiXRl827fBXps84Ego7ZU7fhIt/s8ZWMGTGnOAq1iFhu2sY7
UlJ5jAtNDlxylVCTdkbs838UTwXpPCGiP1TvmRS3JKQ3TfOzNohsx8sCONxJMZOAz/8etpMgSFbs
MFbD2OR65+gYE2eO7BO0mEv8ymYGTs+CXeOoKRO7oXrKk3EOsiDWSrUGMJpEc7JWS4Rw86bWK5Nl
ZqUYwTeDPbvR0PyBaF3lDZ3Emb0JLj6SO9G9dSjGbLPHO5zno55bkHvogfOSVBATpIRhAXqyRGNm
W4rrMPSh4YxDelm7Gtwq4HKw6sd+Uv7Sm3A/yvDenIEaDZZP+8KundW3BjurX0i8fkiTWEczsXEm
jEoUELCANol7/aw1jqmivnMb1RgYMr9IlgacoeTrSxZokj18eavT0eTlJehd/Q0CvOB9OhdVeXe1
cpPFK3FPko4HGa6JoNrW86xo7poqEeEISqL9gugghTt2p61vIs3nBuI6DB9fyN3/WDAcD8hFWKAL
zRG77Wnycl7ifJFrLTFM6DEMq2oIM+9flUtfhIa1Xrz1atUWJ8TjERm31UHZEaJRsev+fDQxHEQb
kji3Ew52f1hiC51yPSD0qwB8i/Z0D5Pu9ubj8CwbguyGMWHK91YAgpinQPIGlD1C+kt5H9S6iutW
lIlJ5j8qVRpuu+F/3bVmfxx33iIqREGAwYCqNgPpFXwbGpetgu02ww5NmBSOmfqdvs1pmxN37Krn
K3s/EWn3Y29Rx0QCZIacKNZzkclGn2jzt/rPDc4J3tUBqImgiztJSbl/JFUblj/H4HqdmYlE8a1l
c62wj3VeT1iKW2aCaAqrbJCPW8C70zHNBVUn5o+ogkLV+Nwa12KJUMfPzyFp4IBgX37Z1BFY/XGg
CguNnGqwADr8KmCA81fWQ7VKjeqmqBUoyz8SfN8HzWk4NwOAEiy9obRRGbNQMaDgtH0+NdKyUEIG
mLYRuD2maczJKEeQIJ5Gi2QbxMPYQ3qMuf7Op89HCAPsYE6tc3UdC1o25Ndt9x9oOUPFv+Ldh1py
/cW4JuMqD+Y8HV/9HBb2RJWjb5Tl20sSUCEtF4lh0y4h0LTE8afcFw1RqV3UlyBysKZt9Qro8IFv
KFSRg0S+yRI4lHdjIFNKJXnmy3OE4/oWiD6Z/k6iqMNvKbz9j1/nmufPZjxYPgzWVSvNGXOtrqYj
NK4WkMGqPqP5AF2qK4ruBJh5nc5IWHgpBKWfRa3o4Nup7+j27B44QJp6LVe3+MvTW22RnsWds11Q
8YU8mT8AmGTz2EYs3HqacBdz1vFk+KGD8EC/0Zb4r0Ii8iuuwNpMK0/xd84Om4OnCi04Zi/j5G+k
wTQahP89MZTz+ilZZJUsxK3eE2KROYTC5rphbRZDoLwVHBU8YxFkH8kOsmlLMQq1Cv7f1FSYdHT7
M6K1kouH4/uuJQuvhOsfJahI5FtvgmNN6dOaJhmd/TPLjq/Q9lpz2HtD2oVhNUbEHDjuqbjx0kmW
7b0bM1exsfu3bnhFLDKyJPTEAtFCZvNC8kOEksjUh7CafDfWvAfpve3A2vhdGznv3JP8/x8u38VM
/odm6Azu6q9ZmDeBGjnJu2iecZM5a6GpinfkMv0GS8Voyzm1UqBVTxDWDUn6OaTv0NKOr0pFKSMx
NwPUGoMbrnI9G8jTrkPbzch6C1tDEReIneLtDiz6T5IRKZRF0LWUWSamW5nojpp/Aom/QA3b9qIs
qP2Tcgb0mUW9XQ7OjcibfGHwxN1ATxXi73eyouVPqEBxTDABs8Tewc5Q8f+ECbnT5mnUTd33nzIh
p+MLenqk1mJzktuubM1fuDJ4Pt/P5n3qRMCIFDQIqShF3gKTjRHBshJow3/hWxQqQftdD85VsvJD
0lpI4iffI+ObPbcppyG2B1hAl4Ho7TZQdZCcFeDjOVZM3ysVoLsnb6jHtiBZ6EvqVBkLLYx45z3o
Kkmd8qO2dw4UPIx6JAA7VX87vTVuasBo/FnqSeDk8sqvudatfs9keSP46m3tMRvrHLNAHcGLYVZd
ylvrVYLmI+eWaW0+a3/TnZGl60Lh5IOdMdJmWTEardu5SHTbaAIRRspk2ILFkHgZTmoF5nJBmsQK
esO8V6pvX6FMBP6gezoCg6JieGUdCZ0+ztYlspTk1nS5PW8cyYbUet9FWlAVjgR9H/Rn2U3hVbA5
JO7OOpoe6MmptosIOwyQdgZjyrLFUf+DRhbUq9spUt0w5AEs2wtDTe1fqZVYyqtMtRjndL8nE5LH
qV0x0OuJUJ29yARbphHg6U9jBEx46c8mxYuUPJ58ABOAVj2Lq3gCfMXE3ryYEExdbDnHmARrftrK
YaJ7lYYV32SfHAytaxVceoOdGXMV1KDfdJmelc+c7r7RhXEG9ovx3Xn0710iMXsN7KY4SlloSrwm
s0CoG3Ymqey2z0IomoCIsaJsmX0oqmNplPFeN14RlMXLJ6Yj0nC05Doc0KTczJdkiPrXm7pNhWQZ
pPdPX6Sockk1xL3uPPjIuOdOL4NQ2ap2f64bhezLoGIGgPyMYQUY9Ud4HzPguS7jcy49rsDZQuUi
z6XrfeVNrlHlH/9hRodTBsT2lDrUNDPYlrtm9Okl9bNJ5tGh6Bb0hLzyB7M1Fo+0YBxT8d2y2MUv
XSWxCskjF1wmkADbzXCEHPJIBd2onYr80+y070rJ7+t3rABMSgWVSs5e0Xc+mGVwWF8IcvnDHSGJ
V517gihX9vu9BqGMNE9WemnAGEfWS6h8KE5sxCyIRhqhaRi95Td+gDboM3yjhFYcJTyGBzaFogH1
94zv2gumMhHQAjUXuw+LSmDGatohvLv85UcNo9WolI6DrolzdwVKOB+L9Y8baYsPmI4atDsLumsC
M4d+1w2Q2iUXl8XwAc9tJOnKlJJy52/uihxNZ05OSri2eRlB2HVdYkI4A6Ow23QOrmqdWE/GqP03
UmUuWBxxWo4jkXTVycnxyMzkBp5psPpZJFDjwUhwbw2IIel02wKBK6s+4UoyKjQzdTFtUSzdj9vc
FOlw6YCvR2jP5jxZbqNyzKvJJTouLBgkHK1keAgZNIS7Qu2H8SCGEKLdUBQjMEWxpD3w1bk5xNbS
dlRbKKfwtOOHeDefpZQaEQXNM+/sbl5yzslnNvrTfHXj6eQo1331p5GpD+k4v/IrcX3KHI873kW+
jTW1RJewEwvqw6Gf1/uOssmrbBvmmagAw8RNLDk5OvoRKfeqm5WgvyXixuE3tX/sCFjg6KxgUCqX
mGZfJn0fNbR25jb4mpcifIKcpN1hLXG30G6+QMtuo35xtvsdi6XHJza3LY1KPMlSq1OgwTtpDuqm
4jKVAhX+Z0PiJ3AdmdkH0InIVkjk2Yulok/YQtwmpStVjkRqgxHbZ4HAEqyntCIOsz0L6y3v7gdI
9MZhkGUn0T+VQyg10kTwrOJTPLLSseJNL79hpPTvCBTMP8Cmkbh5Ig7BPhzl2WC7DgVv+fpRUi/P
nH7FLu+34XfPbC28DolGL3APHcPAIQKN+isevIwz9pIBgNYQCQxoXQLwfiiSTGZaMEFKwFCpGhZT
5pVfhaalxsC5TYtGag2goG6IwMdn77bSkoul+0OpmAVLIw9VX4Q6nC+ybkBoAP73zrwwyfLNSNR9
56YZyBWnUf/ejRMMBnEDSEoSVYnpiXKVX6Cy6LADq6i/nIhU0+6IuUooNWq/9FcqbJQ3v3lv/uPW
tBMziwEliKf+XT8aTvCPoKpYZFzdC32opye3N7fUT5RKyPMGjVGF3bUIVjhtIyIHKfjvF/WNLdKx
ZP+7HvdIWCFNG07rUxNfz9WIVFELfT4e1P3GBJGqNusekcfiYcVWJcyJoqwFaop5LHlSNWDIQbBa
xo4Fvd6mtp4j0l4oZAn3wwr9xjwSwocckynWxsiEEgiSsegaz+rweJSMu1ASLxTCfACZ7wsgyDj0
B0VuHiOYzlntbmlG1xOjsbB2IUjT0yggIWKXUrH/0h50tL9Kdrj11fOmYawAjXHiE+b4jdwhhV29
jZrAs9uC8z63uYxGEZ3icSMoVcbTHIAk1GA/9GoeuAY13OiVMXd059Ls1EQ7FJrPEEtw+elfGXcA
sgAPUaevmSs32orxbHV+mcDMXHDD02Zr0yGX9czZtpXP9m/q7O8FK5J9/JRwWxuRFo4PONs8Xr06
T/YuVU1blPW8WyzTlIEFR+Z12ce2JsZp3H32k5ZihJbCewjDICnfs7R9S7ULDgChVAJsxSMNSBPp
S90keUuLaFaZ09VIOF3dP/cl6VIvxCc/tWXz+56rpryBrGJQu3pZK/d0qX2FRVfNy9xD7whPFrdG
U+mfPuN0jsCpSf6XD8l2Y7O/c/XQtLXLPQLfAauu3B3xjRaz2g14uzJrrJfVhmYftgCRsm6efOL8
L4O2OotS6pjdvU1bJdZHHK7XKwnIQJFs9XC5rgd7hpOwwQi8mwWGF5QD5s0ieCsaj+CyJnWSS1mq
SDQSG1+VpKe/jjPK9sje5rdWPWqJo3bdrrRm9WZfj7v2a9/Hkzjah4GzJNUK9LLf5YkiPjFR6Ofr
KYr2PoxESJJKV/nHE7EAYfdQtW52E7jexHAM8sEu69WrGq7fsMgoR4ZViMtJEldtGmSncenXfEYT
6/V8iDw/C5/UIISfImYQ2hncx3A8WQZfBu/mlvBMTh3dsQ2g26Obu8/kvC0Us7e4GnjCqXHD7HkU
WiiGuf3Yqj9WvQnadvrA6P9MNaEKc4q5ZHJGmRmUJ+iwuNxKseNq4iy1uiLTaMGm6SRNJVHiJZpK
M/6l0HfKbAyx9keJzpz3b/xFDvY2U3i6RvMg2rCSL0ALvzlJU6kIeorDZmY1l83RU8VcrhIfRcZq
zmoB8QcBYXGG2Bc/7rlSBEkKBohx48UCg/zGPHyl3vNh41pfjZABKsUAIMt+6A24mlEYfP4py/yM
zlg+t2lPY3nbYx3+uAIKc9zwW0mLrnS7kknCeTR5Zx6X1uT1H++qaVq8pTsQIEISRkyj06ikRqkV
nWPCqQmWc+zHFXiz3C8l915YXazvk3RYOdyjRtkWZTlGh2u/bl3qemSAiBzZdbzx/FpwqWkPa0Ma
EjoeWmToOlhAfRgkBuccEF8PAgJzzeIc1kelvLmP/dYsyjGpaeRMZSEkHdu+ylW4V/+oDJFURqS2
Lah72CmN2gXNVhVDaP0U78LB17ifSqTP0iFuQLXai0rckLNW3TzGxENC5kyOaH70ScnmRBaE6yG3
VimSvEVu6JcJnDdwhbD8OEdYx/EujMsGI0wKVXIRvJH//HxDY4D5Hg10GpJaw62tqNrsDvReqOM3
hnBHolGq05tZBUNv9JQkqKJUnGZW95PgSCVW0pB/u973MqRbvdvm3c6As0y6sdVj/IL+0BlGouUX
b6JWRF+/3v5L07gGwCl+wCi8iaY6HWyirCZmJKjoLdQ3PYZSWmL+ErlCsw11xc8vSwZvEeAf+Gul
2MLMixKO1E/tkROxi+vHJ/LlaAm3x6LuwhcZ1QrpqvhrLFcZUr/Phw2xyWtzSIX4PcXSY1hqb03L
Dh8QB22+WFx/LqJ0xFLzZJESxrpYrMQXp6coVml0FqVxmMxCbcpbj8mqAF1R3U6r1xDWgEHyXIzF
Skchh2uj16qRnvjRSPaL0JRZXyOvu+NANSuDXmBJMpekJa1LmkJ44YUrNhddWOeLwew+QDBy+f7+
LSyCDbz48+/9dFm2nQyVizG1r9uCG3HFby9XFIBgHLT43/5b29fhn4q7oX5YJ8ouhr1WKmltH9Hk
Inm7LKLAYy6r0rmqUj2C3oEDp632ZFqah8D4oWaYFvzLhSXAfgwRo+cB4oWTNMiP3UZ6bu0OJXVr
/3ga/fq+tULFP1y6lpvfSvCO43XJhmSgcZWKnmx1mmeVO1H+bwX9cKMbfM35nCO21p9e58FVAoLH
SOwNx7Lex3rXeTUt1cijZjUuZjtZu/Mw9TzdEpTL4d7agcZCQm7ZWgit+DRf9mvK+m1P49Ctho+c
FApDxKb3rB8ve8bZ9HlUcehOPhi09gxQ9D0xsbL3oKiKOpqfGsKEaCBiLGGAwvb74BssDOVZ8l3U
BDhyxQzpBhw0ap2mbn+7U/JlPDrFidlyCgXWxZwujOkuYZ0b492j/xFOfZvU+NGPdphkP0D7rBhg
ZIdb1SVPXaKqbTM68Kqhg6EGEybKKnVRvbesJ5dpJ2FUcbGjXPIwIqg1TEehcG77qMfn0Ug/AeQy
6CwF9HT+NjrLwjcK3w3sQXfqWVlmoedgTuC1qOIdPoqiUKD6vgMX+p8ZerDzdiapN7dX/4ppuCAt
oC+Uq+y9daUjRwUShZOSixZwmaLE3ddR50aLr8bDsslfBkFdDvyvGojuCRYQWI6WR9luCxZy8K7B
5uQ5eh59HzWLtOt15wEKlvjIK63dxDzHUfXz869q8Qi9niCr5vgHy5HE30n+VQjMjJM2RnFUwiGo
WhKmZXnnjM0ZRQrsvRtlD2AC3E4OzkUWQSD2D+6Ey3Q5zl6wM0JHuKIQDS5pXjqvhiqPPBiXrjbN
sU9h7yKJ80CJVQq/C3Dq22KK50wJ2idL3IGnB6R6tIOVulE/K1S2duL1NpM3zH+ec2/Gk17ZX0TM
irdulQCUgAnnCpZhN08Ez7M+8nDwEpbloI/88YM0ldrRa+fZMfwnafeWk+VAzdnyyRx/C6k4P2ko
Rx352nsFbbvZXI6/eSfy2ZFKTKUmFBX9bY6cL85e2kmPfj+lk8wO9d2OOy/5YTmbiLmT+nANKKCt
tgXUKb62O0MujFiEDfpUXpELOOJGIdIHAxKbF9OJIaBZKwZDS5FSG7lgBqbvb8s5xffCywCBH2Ot
sA9OBTjjqoNDoyfN4c9D2wECl9Bc14EtFEj24bYN4E07OYvfHSCNY3ts8BhlYNIXzh9GMv84qaqL
kvgW0udNGUVxNuNX0KQSDgumCEj5S4rOhKwCpaprIfm8oJe61pfEkoAqp7RO3nvptWzhoMxykko3
XBh3NxlNbIYeJeWCRTwRfa8bapAYnNjkJXByuhH3qiNOAAM3H8oRt2dAelCYt/C37P9LU747oQs1
u9lZ1W+qwbz7oKYcLtaAuj4ZppSurfF0dCSsgfz8EljUy3yv1qlgZarMP/Ride9Kyx4+1j6BnUe1
3TscOOeKH9LbpIzp++0uFhFIjjmfn7EnQKhF/1AZ7vx4+3QfNl+2yfNOKvg9TYUfnAtdbrC0hIoE
IwW4WhMrAvBNg8iEdA5Rro9S1MoPb/xyErOub5JQBx4YSjNEpXbt5p/dKrIL8dN2LvtH10VS0Nl+
be32UnJZKOz+fI7Img0xDRi4ogzVlbuAOSg1p5+uIG5Q90oUwu/NYrFuhruZtKyC6GofZbN3JBlG
tbAAq0pPdO3wgXSACnkTi6wP0nSl5N1cro4gCnN96S+qzmoUqSHbuXnMiaMmhzwwc0Lj+LPNODt+
NPeWxWktqo1SoTmfq1cQ8OKD3V6HZ9vFegSjeBkJiWP/FbR04tMhTta3pNQCj3JS8bD4awFlvR6r
Dk8vxXOX1HfT233qgoL1vkrSIoUbFNTCV010vbtfJYi/Kq6gRC21vf26Jr2wR1wDCg3+UTDEcni6
G5fZPXxn634GUxEYQHNzdUeuPxUwKv8iwTDgp/uwfDUfvAWOXIwbzNXCRpvl+DCfw2nbgNGy/p+E
OUeX8i+vP5uc9Cr/URvdsUYyi6J0V861rVseeOARRcIx1n0Fo5XYzZ1fsBvsOfPF0uCd6DiFO3ZO
JIUg3iZQ7xZONrRdg4MKy2dq/UBYv9fACf4n8oPrURopqvSR61lAQ+XjW25jBxsRvYcJiQW/fzzf
h9JOQO6f6wEH4fnJiF9Zrt75uB1uRO4t9Z6mVgQMH0ojA88QIPrFJHXsGHoze3kUYd/7q6/xUyil
qJnljHP7AevOcnDOTREEdOqZosWrfTPghgYFCYaXWVMSxd0Uhvv2m1H3s8qDX6hYukGEPY1uIG9e
2AEtadj5LmWrBC12HwkAhuQ+Jx4qqbQRm8F+1y+F4Jf+Lsf5ZJn9NFnEpQ/V2V43U07350GwvQnr
XxNRPd3OOJ7Ciu8et8BBseKnaEvTwOS+qNi5//mcoWnHhKUyLf0tpS/kCeOX5Vh/lyyHw1fklL0a
WxyUrVRv0f94BU8T/AqII/xadTS58rTiLddDt6olS4tSgE+r3DdvIXyV1PUTUI0SYNwb1Nj7Drz+
cHu3MosLBTzRUiAOXeatOzwooIdBarxKWQ1ylxL55H2EM3T0t4SnWe9UrppOeUf1vKHZh8dEB0NE
o+QgEgoiBVkygxBsztiMCCi78D1GsFiMXpyAvUnL7jPJqUkkjstmnqM/yjbCeKIP9Ib20fzaxU5e
4CpCBs2SLDY1Z3yW94/TQmwEWAH88NZj/Fe7mqVCklqfnFau9SW2gxLK5GZo8bYkUZKZVs2IiCaI
Q3YY4zbYToUO53/5M4EmVBpmb6If+9ASR40SUjDs63ngItaxzTuN3J88l3snWgrD9ZPivGrdDE/E
mwZvjpElnThbOQY4ZCF4KAjWM/VZruGAcNhUfZVvVaPcvCg3i/GJYdUfJHW9/TKFD7mw49SdCdPm
C0ojSzDRUP3+XlBWhO2QOUjgp5c/GgEQ8y7T4gxqNfPeDn8hIrlfM6gqsXCEvZ37c1wtPo+PHmqF
o7E8ZyvXsfOCpRvIJk2HhLJMRhheVhdMZ4uHIDYPNn5t3oqDE2TYpXSzrNuBz5N2Q+Tc6Yx9QMSB
PFtGAFygUx8Z1XERTzG2nGBGWgD1oE0/Zi4GIsO6lg1ylLkJ73ozTJ+RfgcewhrlIqnX7UY5mKMh
1Eh6+s9MjKgcZpxkXrIv/MAHko2dTCwuB5kYWDDk7KzihBdLjkPHxCQxu/X8RNS5mTQL6PdWdphh
Rvbs/2sbojlNM83ktqmIR8jmQu2Ye64FFybr5JeHvxQD8IPXTR78Z3ZoGn4pYIe1EW5oLW0JHLdi
yFIOiwyKk5yrRC6+HSp2fG+cgDP/ehiovqpHFJMBOSItCTt9jbRHh8uPxn9HpQU4XCDa0bdRpWGs
wpm0hEJ7SUrg1zLlYSzZpLvjtHt5BD4y0d3uyDALVoyvbbBg9AGPEjdLyLmAg/O8a26HzAxORM8x
DvW4rztUEvRvNpO/w4+2H6qVS05TB1J21F64ehoaLCvTAbR4cYyzr0UNvllRCsP6YeztjW+je7ap
LI7HQMzlcizm3tYFdL+TtlcKytmIGIsUdhJ0QhQ4dNeHXNY+Rkkt1D7cVG0vF4St59PgebgAl6gP
75HIuXQxQwwCrEjQtugvdd5djGaEyN+dnebPdE+wdD7uzyDji0il+f+ILGFIJr0a0fSfDF1bMpyt
djP2HeyUiECzkGuxlxkhPxyfO21epbJVQ6cqrk40f//Ft4TzDyIu7WmZoIWoMrlDWj1WjeaqffVu
784iepQXzrLa8NakI3ibhufjssti2hEZFhkkKlpy+Zf0o2aStEtIjcYFu5oukqu24+NxGbEbKiaf
i93cIElbSYWdL01P54L8shW1GIg7mMOhguOf2DYrCa8S2ekG6fjpmFFlov7yXTan2j0zCL0ljwqJ
7AGtY6hjRMi0qpkgPm5FRXgpZEOLDb74g/16OO+mXL73yiuMWTd0Y57Xxagis9bDQjuRgoJgKwmB
pCcu0adCc9bSZVCLqIsTU34fATPT9906DrfBhnEnpwAcDja1YNkkZCwWG/YOQL3m/b68u99RXIZJ
IAS88Dk7esbK7dP0VwMR7tR07i7EyUkgGFzhcrdPpCWyAGm4S0nmhkHsvsNoh/Hy4zpvi9moBSU7
IZc3J7yJNcoj4Gk2LZx26N85iY3KrLrp7r/Ii+slD/QJS2foaqyBeVoYAOvVEtb2qW4cdEiGHLeN
Gt8FsVChc+Q/qeVY+4fP72pqXu+7jmu8RgtKaqgnFx8hG/D4537NA3HiKh6LBHC/sVDvR3DN08mB
iGdrerlrSOfxTkUlh5ZTIaAi+VyWFu6GrYkDpH93wUmfshiEyprfNdeGqq4IqeKvDFUAc617ZsG3
HiCxsPUEjDXrewmt6mfiC4B4Wv5ke1Hh2/TYn1y+UQzCY9Hv36F3oUjuuyA/SiKyygE97wP09EjM
ECqkSyo3bUfsEgvdEtOiI6mkCgbSsRAs1lt9c5TnnITw0aufbUIfqPc6On9TQevk0e1Acllic8bT
o5OHB0y9NZDEcyMaaZ136w5VP0QyuaBUi80SiKWC9HCv2krWvwMXPjMMF7H/ro5ip6VktWeC4x5K
CAkMruQFWch3smr1tV7ZDdADtbqlw1Bsn3++QlEEA5m7ZaMgYoHsK2xlNW8R1hETMG0GVx8tLWHc
E0KCn4TRMUsrFzRkmHYVnsPA5uwQSYclrdY5uWRVfwp2aB9sc2h5an9QdvTYzRPW4miA6bmShm8L
DcwTEzTJHjt5acHzlJCZPuNeqUdqN0VRMhLUfeJXspURZqp+Ngtb80F6Kgeg1jPe6u0GXXGoJCUw
xs4rKR4zKZbfPzGEXf4iQP6FklRldwu18tpYtI2eicDazbri8cfIFc12uQPQEAHaJgHsV+SPKwnC
/8jIpAMUZsETH43eukWnOpYGVvlv55VbK5fnkfH+1IJOFp3mNforbdEdMdRjXygrR43G09EETd14
X+LCCS7Z6As4Pbx9GGVU1g/YSvS7mvAc+eWnNVtG8aFHe9HFqhluucrpVKytgBD1DGhJzl7jpCUQ
8QN1ub6QuAbxVHwmsno2Aic43goZWorI26tU9e8F40i6J34/mpiI1SHQsMNQCrmTZ/MrGCzP+WkW
+Kf9WoBFKDB3REX4g+MxQYXKbtc/wjYX8xuFqglYg8FyZpGdok4VxTq7LiqHcS0eUkKT5I5yd8af
rGlIfZ+eQFELNTVnugU+n1zT+VZ3Idn7wKOPhIxPnCJNm0ChPfUtcNK1ssvekf5vLhgjIrBJpexO
etB8sxGbvotcBg+wvO1+WpjdSCkZOBs6KDpk0h91EvaMhJsaEysslMYD/xFHlPRuZqM6BXSb914h
vDYNze/Y+ki0F5hcOHp/qtTqbmJSEg5FGtBoG2wc4WMV8beapC9JvHb7WJrZ1zOW8FR16Rbq8MdO
TBQIU7D4bnRiQsKnmLu/bVSfv1ymgf2eKa7PvLQf7st371QkoLNNH8WDtnpK4RflcknVkyC14Ysu
WXRH4lc9NnYK72CnNE1LSDWerF5ai/r02p0q/7lYpw6BoMvHAJcdQwpYbkiJxLKTZxRBH6qU7ph4
1KXYXouSffLXf+oZU4ygDuRiGIqCxMNQeX5ehVJQvqUS9VXvegwoRZtjMEzwHZdAn5j5gYFws4Rq
ziVg9rIreiETHNGDpeeQ0ep1hU2tJMwKkTA5fM/eY68CPZNvdDgxXMCRz/QThUglQ2wOGyJgjW5n
78qrnhSPFtcGmKfY4OSs7IbUa6SE2seziHEUSz0zc7mgJkCt0s1VSaSHlgvDnl3CL1LyCRSUqmF9
IV/wGlt2tFhr13vi4Hfj0mMwdCsVaBNO09QJ+YmoBDf2VA4NSa29BmtfiTuPbqa8ocwLh1giAf7g
l8ve4cEF+iZcc1/8wqP/fgE3SjGI1hxkx6e/48yliL5xo30Jf/L6EuyDz/97ebyknCgJ27ir+HkG
UVbCJF3kR/z/hTO31uNPYEJHrgIx2+GLzfFbqe5VYDfth3D7MwgJpGvvuzScahTQfciOApfr/Hx0
9+uxNgq98ynMpb0YAEyfumD2PSlH2qpRUjL2Vrk2G0Au4oQiocP+HtyuxMYg2n+Td56D0Y5Kf4QG
LjgsgVgtGdf7kKEsqp9lFoNtW1ElAdg25qc+OmyspwUAmgDWWkclKYUmiMVyvYWOSMMxBoIdS062
qigZNRqWKRnN9+sdgmBTzYp4mo7g4wAiY9lVEFR86TAat5Dwf7EktXWXuu61d4KjZF77GmVOpST/
kLVkLAIsS5JhBicIrOUmJRpzZCUapfHvsxmPCRUuYgENLxKH7r0ltfy4eji6Xfya4BrS//dAh2Hf
ys8ooSpF/JpWLL9g6oUGsIPWLWtY8W6ZGZZv5HIogxdcM6FoYyIw/EUd5HNlpH4A4Rn2vJux2HCr
d3HN/KEHwmC7jG7alDlSNuK08wMMgyepULBFRsc5qTqlcrO5T8kUDdP+HGv8AE0DWGgrmBNuztVu
B1VN5XzRtzPj9qdrECNj5DEyetAVvdrl58164Wmje6SxNeFhRpW53ljFZzdjQt3YBt4OpQn2d9um
5oxQe7zYTkoMlkMtuu0ypS9iUT9K2Uqzv9JMdVX/6DWGzJIqPKcnYt+Nzdjzb2yo97trt1k/R5Kn
byzwiSszVyv2PAOKp3y9Az/y9QTi9SxVRTwAhBhQPpFiY25F4lIgnOFjJ2tq7cZhdHh/4wis3Y7N
13oyqvPxdsxMYXhHgegjiUc3AVNQDV4ngEE0RYS0mysWwzF7uQ6XV42KdaJ7Z5BopXYnlt0BCMou
Lncu/c66HO/CNflYlywa23v+mCYZuW7EN2afrwpP0LWE85UX3W8K2/ocbs4T2QRyzRBWhr34nCBD
NukKxeYLIYwikoRzN5bN6JszyG5LaJrRLX6o+JH8eTDeogwl9GHc9OILgozGWGc8qR8+/BnDCIgU
eh2RBCQ4EcpUqb/KiOpZqIUQR52tyevFSnoQIWsgCg4H1I+R2byJjgAmsZtNVwxUSu39GviXqk5a
8/BScj7D1HyazxX8D55DUkJ2SK8ZCzhVTHRR/DTmnImpMW6MRxwp/Zk5c+VZVbERoEUnluqSnFm6
XAwwzmA5Rb61xv/jeBKIn9jBXYWvlYV9i1UKhtC2rLhrzQikKFgfKM+1vZXVCR5t/i+g9Jh0063d
oNhuIRBGa4nMLzMg43wpZLTxnOXEwgQrt2wueMso5s1guVnmo2q2KT6Sepjc958T8lh/y6ZpT5bh
MT3AmXWY0/pReLT3jaqkgr6EkpVvJ7y3KQ5z6Yw+3macS53UGbM9VwjUuKgaEx/zD4X0lJ7IS6eW
4SWWQVpjJY/4pUeK2DDbhfysML6KO7A1jmvXtJQ3Vbhf5rI4qlQkRumbSmE5qo+WF1Fs6qq3969p
9N/v/tGqM6Cex6jAz+RH9NcZ7yYCRMWEfyvDYofPl5vM6hbdbhBIWOikFzuetK8RvDm2mBGcplii
X8f6eOWwQyvh9zcnjslcXt4L8mVU1PZ+THg6yrqr9veN27K/E2Ge3uJBXha2KCOkPzJLce8409OQ
lXfofesKrQjA0ca9r8eZKrALT6k0Giy8Sb89lSk9bo78LUFIw89qeWuQyFO3NUImZGGFNoq4atPk
fbCIT9TrnO16xWwTAPnjmbJ0BfL8yrTKDi7+JeRWbZr6MMjauFE+3n4Ean5d1tZ2nEKtDLvTuK+t
A38cfiOBYEhwvP94Zf2EZ5GPUjdivQxZG/QgEgz3hYboU+YLl9FwHv0+GeOZ6DC4irDxWi9GExqa
E554aF0aNBqjdN+Clu8mxFJlgXFeWIpi+zAQ6lXzksELRKoGJpYtFWkDre+/0pi+zx1ZrVVIIE83
LqfHAYpPWtMIKHmAezngo/7xV5DPMgJo/mh0jv1btH2R43YkK7UFpaD279e70xgR4fBL+Nz+4PTw
TSqOPtuGvnChKsk3nhW4BwV9rjkU+7RgVvVm5BLLN6IgI9RMp2THIisWMY2eMxf3HwramZ6Vg5E7
vfSChhLM9D7bQVOs22NQQmKXXRmbukuvz/Gt7hi5rt0j3JjPIH+NZDZwHlosFQQImDeglx7WKqYw
OA3msKcKiPwYoedzPw+EtTS68DV73L+2GvwBtQGNPTnMOWLlwiPefwbtU2+9aAGlpq5iG9HNas4+
qX720CP/FuUHBNTF0u+Vx396e80IVlGBYnX22uuqKrxmaqmiQ1D5mYYvctC+eK6XocLjB3r0weYX
Is+K4wu0vdDyouxPo4zloeFBoww7Gms/hr8tzN0T4d2r/H2Pa9/E14mxAK/lWSq+xJyWYckIiUuc
SYiEFbCr/9TpZvBVj6RgLYpUb18B+8f4EdzVAjr7TNySkPw+NksNMbqzzkGdaGta10+eQgchugB9
osdmEalfYRKx7ZQ3ualZYrlKCRkH81teua0mz8LASa4YZboUPVeFkqZy9sgYDhkwSGsAWL6cxac3
j2GZWii5Ux+9qVru8pNxEk8igXZI3PMWSTKZm1wAancvFVdomqqZ8VsS7jGl+WkdLwc/lo4FJJPx
KKNsrVWRfchpd99Zxu+NRyyCzpDsoNVAbP/53oI/wprluq75Pz3tOYuLt+uVwozWpf92Y+JbUTxZ
TJfmRMHW5SvWO/zyyg2dkae7pXxwzbZcbfvHMkzSs5w8S7SyJX0E9oBZBqZf8UVPhgH8UuBcb7Fa
flxRop/ZLp8vyKXF8cKYo7xAxV796G7FSQi7j5n7L3O3uHm5U2ZUbxYZX+V795ApbZr2GTIeBX2Q
AZGkvdIhRQtTGz1yEGGyebtfYC4nTFEpeqxdys+8km59+iJ2fTXkAV1KqjyfVM2dvb1uBv6Ix5+t
kd2Js6Kp1pYQ2Jpyn+w4syoCNSva6fY69IVBPM24uhOgeLcqnlhL5S4iQm6W0iNkor3BpAWBaMZ7
LFh7PUO4mjlj83HqCX6ykCMxY9oz7RUTKPI+peH4wjTe6ZMMxgA+rwCswCDj3D7QBXpX9meZlLjg
kuYO5LImF86aX80UISHomFOeMpk8oxPpf4LBuXWOAY4y+MPAyuptMP4WSp/eheq2X3CQM38f062D
S6pngUAmPIIYUKfTyArowazKJrdXvT/0u7TkURsri3z/aEPSZ7bNfhdWRaui411IsivBBvz0hcwX
80AIKY/0VZfavo7eAi9ctKVNy1S24K+5kwXnpOCZASjrq2qkaWR8LE/4ea9zEiopZh/KjhjOkXNv
susf1RXlef9KuLU8JMPUD4x8ORsaYh4WBdPa2toWxkaZyMxp9rNKVJF7Tia6B9wggEtiChQf0L7f
paNidbrU8iEY++/DoeQf0RlufJht5WdRJOVsBteH3uQx5Rs5sl3i2KWSlcBFiUpbq9hFRNz+2Gan
wt3P7kM6yqPlyMvH1wk7fcHuJtXQd91Sbk6yWX9SLK6eFOVe6vACc/tSAJsSU0KFTrFuWjWPMqp/
r3c+RoOmm5J8uSuboBvzvMPl3o6kR5D/3Db6CrZYspk2nNkhL/HplpCGj7ztmA5lywJ49S7UtZeM
fcF9b6piONWFIzAxpGD5taNu3lKOym23O7/R1z+CULhhQJFBeq7/15LwHX+5YQHWXdwoqcUiyJFD
qLEbWf7nWMr1UZSBxCjyyq4tEsctM8LmMPVDF279vT+yC4VUXM1aeaz5Hq7NkwnYhJ0Mc9SIbvle
HMBDt8WBPtzLpfFFxQErF8eY0GVXgTlQV6Sa1MKOpZTmnZDEBEJKT1ByvIoXNm6Gk3KkJ3FTsHBy
PBwQk0e1xHjc2idINeu3nIILmy5LhjidVMVq+P78HeNk+bTUL4VdWDNAMAhj0zDXvLLkgRhefApV
m0d5NFs/iyy0RfuCYS2SaWdLCRVF3BAQB+qUl2e/vsBpUPJ/t2BH87bBNuTrFY4SqYOtWR3VU5GA
BNKGEi6OTfz+sih2Y+5EGCIyxSj4uGjWtLS2Tn/b2yoACvSMTybFqwsF9zaPVGy+9078mC1RGbL2
3V71Vw57yp1JWLDi3S7doe3DjTXRK8LRowqA0ITjy6zKra/WKE6mG1kGyBpcqz4E7pkz9F8O53sP
at1iOk5psjtlmsykPam4Oc/dDZQlJWi6yNj1+dLvoha3veXp9b1YHum28t189VRDiEvGNjlmT222
xrLgG7JI1ucVT//HjPsowzChSeTvXEsEMaCwf/WplMkSq08yQ5KN3NtvKoNTXGsoPu2l7VWsDCQn
abhEgLXSk5tcW3cOLOPHAxSI14Ec3hvhNLxpbhCKfEiNe7kIynUQehLYk+ocFVswkmTnEz1PWBsU
FzloqUoDRnhEzIxI1xdgiA2ZzuGFTZyptLDjRcB/5tDZWorNpyC6D+RQX164MMCnzDPKqkIaVMBJ
bGgjjC6uJHS7moOH6nADb0ZI7ZcvVaPyPsyxYfldUBAXC/N4JZVlj+oO5A7+RrYiaU0NKn7COE7L
/R5huIvnU7W9Mj85IVMxgQqCyH6RP/rRFllDvtzdl9zugxmO2YnVU5U2D2rUtI1rUchrTooCZ3Oy
MuGbB1HI1bibROhZzw/U9+BRqwGbiCUKzGfR1YwQFrawaPxrYZhWqGspZ7X8XOLpDWZCvGDMVzAY
YR8LnlmXiCuHfifkdd6AJUMGoGpK8Q8L3+kuPjipGrSysLYUm59c+zaCEe3YTPafgFi4b5CR/g0q
O8pZgcS3pR9CzCyewUJab4LxrPBZc9tE7ybB//Zt/u4ZZ1yN0DzlurKtMyXVaG0KoAvh+Y+1FKXf
d05uHy2FtZCg3W27e4tqQNYOOYWG8K1cKf/KPNRlJALLMU8MNNtQ3WnMYUIoRgGx7N/oyDhzrH2f
vITHgXsbyuBE350aIJP2dlUikQ9L7OuyzSsGW/BNpQTo4S4HBep3VGzaqF8smwRy7+rvO3LvjnFg
Z1nRmilyEG3fwgsIVA5+mJ+XDNRxTxXLn1tQ6m9YwzxiIK9q7yDvt/M+A7x0td0+eDszMzCxbfvY
PIbNAnTv0QKyfrC1YJL5H0txnwdpVoLb0C7b8PFbw0R/QrbZiULNNBOdYugsOv+mYmXwJcn9Ekt0
akgZnRmVDjzi2bOHVazzKTD78EmjFHQ18yYyRgcHnpNsUWLaVfJBgQUYOIys4TwxajoFOyfGQmG1
R2bEwxkCq7HXhFZSJDRQl55ssjJByJ0BGHJ2A+cXIKk6b/cpV1tlwIH0qPAZn5zkHjHoV37Wj+AC
uOEls+pToaY1C1gxFmFtpJwWfghdNXQ2GGsPbVeMBbuGYuSOUH8EDp6l91IKhtFoS8BMXOyGu+El
Q/TuIhyFU/hb5mCyQPO1/Xs5h7DF3ywpPPS5HRrSMXNiFhct1ExKv06h6tlfhEwPu6MvBI6doE1N
SUaPOdQ7ggWIIQi4uAICwxPyuh2bwAWa17UOPI9OkU40kQWd6BEpXeieeBzFDSKvQbMECV5dMKOo
FnmLisbadefHEYWXl+0npZNlyf6Z2ekXCWAufJ/wgi9jy8flszFrViC9BvyExDy8IwyTkV2tyg5s
eJ34so80ds4TgtswuJkzkc8UPV9yCeHh6++O9ndY9JbsOMLF6GcvoB8XdWTMW6BA4R4fh6yg0l9F
wrMf0p+5DrCS7zo4rSPPrWfo+MJIJ6anGudWcDuJuNq9m16qHjDZ1fTVB2Q9LIAJKHecPCnCfwjn
QgujZ/6tNfmgxBBhcIQqvIJ8WGV0pH6mz2CLH7vtxWo8KNV3gBbn6wKlU5WlQv+/acp9SSeci+3e
647AI+7KgmLh1CQfSKhS/BDoTTBUo2QbwZrjFPqcOqRzxJ/b+q/5u8u7+V9qZPmmFFooaYZHCv4p
qyCOKQexgIifEz8XO8+IT3FHS2XrV64vPVPVIRHbtpaZ0WaHKCFFRdyL0Hjq8Jevj0B5zo7VcsKX
KPBF1eM4Z1Bo2YuxKlko4wyrIqtAiHicLtEDqgkPU+DJj4K1eCazWooQrioOPRoOZDYpDtdRYl7f
DeZip3maxl1R8ipNETjcBBW5e9NH1UDN3sVq7vZ+WyikCJ6Rp3cc+2wGf5iQFIN9dAocvf7RzXxp
DKo4sAxyMWq4XcpN4qQmRQInGdhutr7/Xtrrd/yYPSALETG2rTPSy/Tr5fA+sdIQ7wJFXBSUdR9t
b5vJFMmv2UKDQFE52DyR7paZ9Suj2XvKC5NZyVMsfvluDoJaxT1oo8K91Ica0DCQEKj4Kt52OAhk
uFoB9fu43X+MK1F83H+6A3p7fC9B/snJGyx42ZlE7PSfoYeoTW0jVXAdVjlrFUxe6iKAkuxeFcPG
sFlt4Qks/d7pLq6a8ZXMyw7qZ7iCflXy5THLK6mUPhJNFdWQl0UnxZpIh83jsggAdJ+1SKywuzxR
8Zc0XpSo+lgY8svfXVrbfvreSfWOsMhut5biWaFuvJeT2NX9qOEF6Ox2h8Pzsy6E9dmJI9in7ZJv
mxxktl8U0YIHxbvfJCrnToZ0E1UI6SObEa/DH8Osxn83WmjGRtCgq0f/4N2atLYw/gfdDhyGello
4yOxXu43zbGXxBljZ1HgKJabhRaFpqddOITK+RvVt8QCB2sDNquuskEIeKC1/b1Kf7JAPr98UPCP
MVMyVXRRYnRr1i8VUSu88WlGWNmT2X1zfyUbKSvDrmBJlX3XQ/cqb3mAKlkglStr8dHwcWM/qg/J
kAWzTtFXwHK0DRbWnk0tPmFGP67RaMd71pzveBB7fVp5iPqhIzL1NJkoneNiMcLkM0wD4VgTv/aC
w7VhJw+mFP4y/HrNaiFydzgaBevncUif/+Pv2NnaYid4W78JF5Qijav3QgKy4uj8FRcRvmKe/djc
bU/wMK8xvUry1vBoo28gtPLrvTp7cZ7hbKQ3Hsg2G24l6gMNiUCqK0T8v+kB4ivH2miqgIM83VTL
QAT45mdt1iLlTX5lGbf37utXBfGmkQ43fbJT5LsO2JPZ2haX+uTHCmv4WjyWSQiywFA09cF4oK1y
vmE89G9d0AY4SSxGFFzk270QcNaZdnx9A497u3c5Uf7PqpD2NRxFJ4w3ibG2P3r4iD35IJgSZaMF
TSG8p1MhFdWo4SbSrLH91MH4IsNTVqdmFbHOZCvtk+kjWWV1MdlgUvqRCgYN1J47MjBFuga+mMP4
6Rdn0VV94sM7rv0UkxAQuSgNL2kNx5qccktXOes0NRYlhp+YvZZMnqErzl+Xu6f7YAaNojHW6GeU
sghXngrZ580YFlw9NW4xye1QWiKvaWoKNxyz0bream8w82V6PEAqBdxG+LHqorVYMDlWnUVYpH0v
k5HurKMS/5E09r+iOBmspRm2xQ1NDusBmTvXJnaIRGSL4XGvIgcatAq6G10go8/ePAzuTYSY5zj+
6o45gMv4yPSTkLFjAJJAyMyxiDiM9k9mjBMNoLRVihWklHqpM0HyJTNPlVhkN9oNhS3KM4xCp3lT
7kL+u5GmfiDo7FlRJxBiIkorLLtbYqcdHY85tzmWAJdFDEyjEbfC5RCyqTKBGB9tDgLpw8hELaj6
VwiIxrM4Fq1aKRIZ83m8642mdHIK/dljGvI+0YEfJ3MdOWjDE3+sEcuj6VyWBRjSYaW5NkFMAIq2
PX/5mKhPjPg0UEnsnqHgvUM47tw/FVrufkrhbKLu+g03qwzJi+isPOADYntRBe389GA0NJWqwL31
y/Fa9rX3+vmBkJWBhr7FQoHqyov2B3VOZa8kjOMFk4BnQXhSfedIDIFLd7snoiihiYZHZJ7cbDn2
PYzwOT4NspPyQLQcqtRbJd49Z/1WrU/Z4dcmktr0O+jJeKEIDMTtnBeKccBWuiZ0qrjsBe1OptgX
IPMLnKlBGSziAlWZP/FUOYnOjg1yCIv7Fk23igZ4PNMaBaER0b9vn+hNITh1mGwy4MPRfPjo5qNk
x/F8lJBGOG/5BjSSqp+R97WT1hlEl07qVCo1ydgNzAE94Enok3Us88uoP829D7eYudSgWdSyqDL5
KRDaraSPcUfx2NN0PXABXSIBxiIllGJlq3SvtLO2oELnIzbnNxkSqn1/246as1zpvUztNFqOXoK/
2jaVoDWkDXirZy9/q6fmXho+U4VjqZliQx/TlDMnaXhnUPli18wJuKwA9hDuSkp4HgQGI+YxqfUF
gXTHRw0h9YsoNJ9yF/dXRUdZoQEMq7CCmZOueZ9xH85Jj+QwszDUjtNSv/VZ2bO9DvcL+LDoLNKV
rXNAtMqVO5a+NkLQZsl4PakfjkughyEed7uGQv5nbRZOc4qhC4kUMOgSAtfgod2la86LSc/r4sgH
lPGxnUxvye9s1xKFj/BK9THoVwVDqBq6fOWPqs4ets2O7Zzx1BDaGEf372L2jSWQ6ro7uE//J+5o
eWu0i2wkkV0TKs/sCYIv/KMXqmnawkfm8n3HKVZx+EvWn1ShSG5eo8GatiflwczqzS+tjxpX08d1
EIeD72r3Nbpk2rYjoaHdMBMbAQX9djhxnZy+bdlHIiIha6pz0pJK7Cu9djGiOo3UzBEyYUpAI+2j
8NDgyb49C8tTzNBnkhJmC+VLAhm0JXvD+oyQP641TwEDVEV1X/VcRqvAXIlWTaDMSRVaFkTKi5zn
9P0srqLvW9KxCryzaDsQOpIdhHCTtW4ykQxiV4Wc9QI3TBBLNCVuI2SQTNqyHa0jMkJrjAn08mNN
x96Z3p/3nvypem65N+LHG4EiN0JTtdKyv+KIkkJ58H0kvdv9MccVSO9NCBjq1+QjjiZG3HcorL6c
jsu9oDsTjyazYZYd82X/FMsjmFrvTgw4CRk04dPk4asoJJ2WERETql6sEUFJ6Xt9nmdGSHtfKtI1
HPUexPcGF4AR/XkhM7wlXfYRc47TRCQi9DwStu6VBl3YaKx54MIFbL+QWsAGEJ9tOaFWCMgCukp3
pHrjmg488cIxASjezY6i26AQfCSds2hotW2eRTovp6/qIXnxRsucy9j/r3KI8sniWsbSsQ/7DbKA
CaAloUdI0T/s8XKNu3Lt8h5geh0ABCGvw75G2dbWfyhRttkB++FznLQlF4f0TbnIagak0jtJBEaQ
HS2Skf8RY/8wvPxbBZfVa5GMD6mpujfEEGGnNEPQDPrsNKPywE+7+pFl4qXE143zuHsFXT3AjR6h
3HGPPvvjbsSF6XeUH3g5qYxcWZZFIgx2cf4805Uy5Dsj1J9sXxSk8OZqaer8cXTeIt6hobNpvRbb
JTg+JaPZ20jyN1RseF101OZ5IxzXTEXLnA9LU8FLUY7uoooBT20Iugx70JLLEYtBXl+6uvl4fqOh
DMHUS8dA/7MAfS6grpdviwaVXfeeOLDBuCnezKaa4TTGFbKYKSsaeJ2ILMSeU4xk5oveNHafF0Px
Ak0mLnzP6PDkcKETPCJLdHCGKA+tkRgAFzRaWhq+GAB9DSj+QQDipoqVZXKKFWbWIzlpFIsMsWKo
QbLq0t1F0Z3Ik22QHMdXmbC3g2ZDFj4t+6wZ7KMiO1eCCywqo4R6CnG/JAlQxoKilSMvAd0Us7Ad
Ho1eE9jZNKjoTbVo0LH+19fF5jzbIIgG1d7VU99i+xEZxA1pf8KZWDU2mGfGSwPYJrA4mrUfgoCi
bTjJiV145wh+0AJUUc5NYHC4/hdambmocVGW6zWcTtf2w/YbLy4X+2SK0rudvyuPPNk5sRTRnrrQ
PAxLMqEMlsGAuqa+YKcko0YeCqY+W9LsTFjSov0zSDOA+Zh9Em9parWiNfBRcXl2jcJzWJ4VmxyD
jDORdgrfxYNLluLN49yiVHwkav3HnW1D7bHvM5bVpc8xIdE17hsXbO4rmJhOM3cUZ6iuqSD9cLQ1
qZEVDWk8AHYNgVSwnGCTOlXY7Ychn9EsnqGW2rb+MmNU//57iEmMg01aIs6lIbgbVv7+IIJ3oxUI
OX+mBLUp2/Z1to7Z5QlS75BnrU0Z7Z565p0Gf/MwCo7f6bMEuFNZJSdPCo0YwYXSRIg3XHu5FnQT
Tlq1PG4cjWA1b7n11uFJOuETFAKJeDeK/z80CR30qFiJ34bJTBEDCBO1kSkm1QgBag+gxwq3EL9Z
n7OjgRAmXef1epwt2LPl1+D0p4AvP1fM4MDIwlX0/6DY4Y+TB3FpXs2I4NzSbClrhjCbjd7rwy9W
I/RJr6u5Kq8j8VmT8vonjoVICLE9rGJnWTYT6FFFWA8aNw0QEvXXcO40KwPsAQfKsc4jjitCmr/V
xAMaQIvQ9qaf5FmdDJz1aKg8DKQiGxlhNi+NhjsX7w9QLXlkdn7D2LzkIL/hLG/u/WR+gS19ALkR
LwpFrmvclF3U0jSt1VQgdRbmcL8nnegW6lAlMZFb9qLZuH8OS5um0q47OAzb0hVyaThFvuNvvG0w
06HmJjLoA6Rvx8co9Zv/UzR+Sz0XK+S8s+6R9/BzqNW3i+9WypIXTYLWi2zEjZ5pwQE73VQke/n+
SBzPL4H7U28Z2gHEdZCkJBIKyJBt7KME062+bmlaJdbx8/gGcCerQItBs3Ym6FxD/rjVQfJnRN8X
kYJ1+xEfwVPpMriqQrK19Iu1UZvTN3pXYCcVmysHusSWHkiAn7jUbinRYuvdCzHKtmuwyc4Gt1IZ
K/kh96MQoOxN9GEbU3xCCaQ6MZq9Btf8v7iVREdjVBl3zMVAS9gKOWSLosXtd1703HoMEgNbiX6V
adZ5YuArwa0E81bl8NwuUFdLyt7nqRfz7reia8KI5dOwIHrVvX+AKJByVPzB10rBRZ+nfSvK8wMb
YA+F++LUvBmvxKT4CMYq5kloXs5/1hPBMeMZhTM5zqPHbZ1ZdQvlXkl/3px3sh4Mg5k9+VgiHilw
JUu5Ip2FxHor22s/KYvqZqq6o6JpX+owNXBvUM2PlJLl9nLfQdSOAAnfhus9rupbCBAYyvZko/ZB
SwXxQIBoVWK4OH6rDT3gMM+nSDpsxNsZkhHr1PqMW7lRYa3ingYTOBYDeZjmzJzRssGL7wbbDUY6
y7cCn7oH67UE+W4r9RCB2uuMJCZqTC1iptOjzJgWZDPC8L02WIZ1PCtOQ0v1uDGkJOd7thV2k37V
m31wDmPwj/0IyK58orROlPedeUkayLxHe3aebbUCV+7X3DLOZBqO65aZZ7dUpRbguTyweL24EA4g
vk5/KIyaGCJhKbdVvRnh85BbJorVq+yWzucYhW0BPD9YZj5aOUm1oS7lnXNB5flb9lrRNqM9BMDb
G+Qt6+sVen6Xb4XC492rq34R9Qp4ldfcQzsjluWoKPfnkiVAvXPGaFuwOBPt82Jg9w2kKMMFy7mP
ESNMWsmw4DFD4OrhHyJu+UKX4BH3tIlrwwTaeeOD/yRE4iXWlZylULUt9k5e9wZzsuAgkw8pj2/h
rix9oy24deyMceMP3CAziE+KtU+8jf0CXHblMv135tb6auAPWyEvsFtbouHuN1tb65RbWLcVUlHw
RcUDlGrmgYB2A1SZkMEz+RuWurMmkglRfQlMSqDzpywYwHJ1NRloVqG9i9A+If0MMsrspRFKHiC8
rPUCWfKk1CZtA910RuesmpFVeGiJq534z5w0WIrAWIa8ogQsjUMm2BXAknPB87JOsuH5mX58WvYU
3MXjomRh0EaE2ILd24pFVLI8S7CwN9yXZNMBijY++wy6Hwr8JGwh4Lb2V2yZbJTH0mCy39K+cQ8B
Wl0OB3BM2eI8lfJQk94q4AzPlmMv5LatXx5cKa8gO0t/5AfC6lC38RCA7LZ+oF6jRzWWtN3tNO5t
svFIIcbPv0g5ePmuAagRknyqyprAQHidmp39m8X3sYg0dstDmetud1cm0w9A+LnM5+E/xkInPyZ4
dHW63UcN5zoVBZykAibbMuyTOFcXQCQwgaOSKYCcg/R85eLNtiGEe/NaVgoE2n5gElgmH18104Zv
c3S/YtXG5IrP/pABB+mR7Spu+d0oMn9y6Jx3cXgkmkxUXsNq89L2jcfmlwyiSZ9vpSsXX+6KLS7m
Gz9cnsDCtRHlljL1SjjxwKYDBybWsTEzoKl1A6mittHpwEwEChagnr35IGx2e/OTkb9viyhYZIE1
C7EhWkn975HD8IN6e2k7HMJvWQ3sXWvxoH8PI6lI8gPYIpAOXiyDJ4C0GTQCMT+6V5Vo9IlXvB3I
4y8S1L6hknq3bxfoSYYVNSzPFwragDggFSMRzP2kvlBXgWlJCHXD2B9xkbJ0jrmC+4P8fWHSG8ZK
Pi7o7MgVy+12UyRdYzlepw87DZ7e//VKlRgkzS6euOP+2uEMKjo4pSRpKov352IdaF3clJtxy3dH
V2Abenyj4TD8xAyLed72q0Gj8VU2whty4WWYp+Jrno7ncinNlPIFC3Vghi7P0CXpiM7A94UuvsIv
stvjoma6Nghh8AuGCFNGHJlYmPxpQEu5l0aYyhHgQh1YpyLNsKTiZk0R6YzWmHa4UAYW9Aevuzau
JQ/2RrLQGxvhdMHDYhXvAdQlxr6SSNgMKdBlrMQKvEoZZw6guUYXMFnV614PDOl3fIbk70DdOp46
zImZrWAIWGKUsoZmqxZe/0/4pkpiNpR6v/WKAuJ50xz6XdHRxVElDGa2oKNBuEL5+qDuJMSi0ChM
1eQohUrXCXaSGlZqK4BQSTuwU4xf3i/WopoMEj0/y4/SMQNV4e8VY2J3s+0KLjTyxesIZR4LuQmw
oH0XUEr69V7EOsL6EqvIRCNhXN0N2dWrtO2pAsj005Oa31UakE+Guzw85f8ol+0lLSgsK0c1HzcO
Xv946dLZXhKjStna70GvdAh4d6ufye0OQgaya7gUfb4bt2brR0ovb7ozTl6PKt3HpCrmWJDIHeOC
dvtKeFrTpyrwsja3HYfu6apA9UCwFV08v6Zljuew1WdWT33spVs/daJHn83WP042T/opJ3rK6PPA
F2CcdtUuRVwhjbRYkGLp9C0VqCeePOk9nZZZIJ+LKuIALGpvMbv2Rl48E1OBCYyXtuMqqh+CLEqJ
tTNBcqSoERCvHDCAqj9xVOLn6VikjBBCMd8tbmIPVVmSPpcSR4/DuL8iBSuq3d52kJDyS7/5w9Xm
NwbU867E8PsZV0jL06f+KcubaT9X5U5d0ZUSmqp3nBVxXzZYEyoDKCD+rsy3A78cP5ezN7o9iA+K
vxzicG/ew5aaubawvCIRhEjgiMQZ6/XxVKXgx0fO+mcV/ngcpBid07mrcrf/Xa4GCHNzjQ/hqkNV
VyNsGjBziHLcpol12AF+vgbh8JvrohWjgCyKOsg1BAKlUAmYLbO+EGp3BqqobIafQcp0/5mt5aAJ
lN527eUMO5QxVyXLdD7ZaBBaLCdUr8FEdGVof1nSQv86w8ObvF+d1zdw7ItoxqtJzevaMxAMzOPF
DJorBspZFxQEIxOWSQ5kJcH587ayTyzIqDYeJ7arh2K8k6+EkYfa/D1c5ugds0q7VzKVIpVJAc9o
oFAJ9u6+t5GI9V6p+FRi8WQOB/1GwaaVkv/tMQamdI4aCquaaTVZ0HMUXs6wGNu3ekDPiWGMaRk8
O1ukcDqMeDyeQP+pJRxiPvvbvDXchjxhhAWPi9ipLaeYc3hD5FvJlVTqhQmU93LNy1bk0p2GfTW8
G7Ghr8I56DyXIwEr516zjk+zu8REu9drDb7StfYqHX20EMJgN+hGlYLyxWp5Mdg9lIictsBZd5dq
HILezPnoKGCWxoC8x9mcAmFHc9AwjJeb2KNzGDP0CNaO5qmtDkjop4RHE36yM2c4Ev8SUBjT1vsi
yYDwMs3jrrbFv36TdW4ddCRMkNR5UhDpAWKPVY6kjtQgaZIiqx0eSLTRlmybwex3QJgs1/tElar7
J2acgqrvScRN8NGQN9/81MuI7T4LQTihzZMMmTJjx1yp+eYTs+DlnOS1xCcnVS7jpWhd9i0HX44s
TxBE4yl0bTN1FocadEpePXYnP19UMhMxIEwI5EP3lcg+BLYO4YIw/YuXsGv0JTIS0PdqrBeaL895
q0CrVsrAZtkXlFoLOQdqvLwVQ2/HququD0TXxNoPYlUbWV41BbU21feRJOHUog315zy6WQofvi0p
F3jX2gUIhXvIeQrac3Rk0Ubx03gEk/oKZA6a2t5Es7uDZVeDEceqhvkUGlQsLavCSKZXPF3PZQan
sgbk4dIT5qrVZGaVrbUtWB6DM1JQTWx5U2ciZWYIlVYJAb6j39tLgcw6aPM158E0nHRWZpg0b4Y1
SWPo+Z5WFHjk0So6mRSyrTRptCsMNv9y2MS2+NT7ezeh9Y+8A2ygvAMnBh0GIx4EH0psI/Z75oRd
WMbrrhJ46CnshmJ7qVAsCxD8MYGwYUNPoOkTztR0p4SnIqcZhtksuGDijINV47gigozBdrjVYpMV
eELuOIkklvcj0gHsrwoJDDr5WsbCqvK5lMMgPdCO3dxeDRvmT86N0kOuTzUF/8w3lhnTk4jYmxEP
UL/+YQtkik4chhbXJ5r06WitE+VaN8CLtT46HV704xoZP/R0UGqXixRuD5UYJ2gRwmrIhyMQJWKy
gYg8fgqQYIJGdjISaroiKM8GlCuse6d0JCRUJFtA8PogYvODMRgNKC2VUwyLXKfftlrqs9MtRtXp
5P4gAHYZKaKJ6vrDofMCx3asiZQIBO6j9pHUP+cJSv+pl+6eww03v2cn7LmrFqpcqdyvzc0mNO0S
2JrH8/qvt2SA92YsesKdu+LpeksO7Q5C8Qid7q2nGCvYO6rUP1wUl4iTpE2tyONSM5CHVk6nps70
e7SnEgxhtet9fR5WB0kRsbBJb/3hm/vePiHgYRzqL5b35nanol8e+lZHRVS2XWl5MtCaC6A0H4e7
kllfJTd+f7hjSBNO2HJWWB66D/Rt1EOSL+7SP5pawan0fxRCO3wFRllVrVBDgj4qcii8+sISABGE
fCqlrtMZJZQ3IyVQ4A6HW8svmSPK8xvoJjiflRSsrcMdzQKVfSDNtfAdqi5tuhtv1z8X02EXlN34
nijGjhaWPjDn6ESGcjYlW3SG6ss1UHy8+405D6NvyhX4qF+yE5JCwedR5lsqd9Njckme3wz6j5MB
GqFsBb/caNn2aEaf7meGvkrObKazbvO4/XFhHB9+il4sQZDHL6grsnNBVho2chs4lvMMviAPfl2M
tqGSkDecNNp4RtpKw60hntn4eHJf3moZCuezGvSOjuudO53qlVJb6+D4QCPJFjSETnXX/dUf8Ejz
EMfM735zNzbkwE9metN8ugAEivoutxlX4uuGsLzNPSGJpTS7ckhLJ71E44jQl3r84O3eFG3+/g+E
icI0XKczys7Sx5riye+jy7mX5/hN7syAnqUiferRPIezGeIl10nApC2Md6W9bUXnCioKlMqQpvKH
d3J8V0JyVABt1/O3lNb4jpzZyZJ+B+sa2TcxFSoNEpnX3t7BtLH/wXyWoMed88EoWNaF/Pv+41+U
6+UXVFJlbOvHQ4AGrIhxx/6/WKNjvBUbVtOtKaXnrz94iDC/Zutgd60wDO9cY7dyWhmZ05rHOGXF
qcH7WBWbWr3oMtHsS38xkEjOSp+702tYTHOeFD+qXPsplZY50A0AqBUzq5q9U7qavW42ZurqTQpR
pxvZ9ynZHpnA8jQPJjoOlqrOKF+DtnoK0RSCnph8FFlZQrH91SbstMoTgv/gc9vtrgF2KSp8p9jQ
rpJFbTwmo6Pc5Tl7HcZ/LbWxuqRAc6lBsfp8KHUqEX+4ZDLkpjxyMBk8kR/3Wk1PhMZ96UGz7Bra
LNJFTr7/vO6gLr2C3zd79I9h0K97Z+ZU8ElvOl96rcxQi6JgVLOzJMf2GnqATcHzOd6htjV0G6C3
0tfH/SKunJYjri5xr0eq08UIXEHCQl2NiYqxta7j85e1/IKTpYdJoUvw/DO58q6ek/4LiOtwqNTZ
vGt5cRdCOjdYIT/J6rsM9ALVClgWWZHX7ZZedcE09isQ4jmK6BT3JkCWU+eO3BJHQlH9Hg57rJGW
SAqXPjtA9nR/cwFI0bhe+7KE2GuCqAtWoNu0qfXMjTOmYS8/XoWvveKkqG9InRUgph6sHEb0lviw
BEyYfEUe26848R5VnKNBpZ6gPz1RjXN0qd/TdiIiVbsYO8xm5GNjCxQNcgYnqbH9cq0XJB+j6Ser
pffDoHBufXioGHjtBDzG/wzwnrE4vzsGveG0HZ6awOuI8vl06pfOmEuSZuChJ8fz955v46Pz0gdI
ZHTMHCZqjQaRLbqi5ephtfjyYHsZAB7nUwrDbd29zZXj498CEWKQXyJgHDf84tWegQlXioCmWsXJ
a54ytXIxQqwi/Aq3JN0RybQ40QIdYFaELNjvY8thgDLImtk8O0WjuoTcT+IGXIT6kCysEhJOzOWj
7/P1leKq0V+kCACkhLrVh8sWVS721643lX+UOC9mo3ZgJZad9RcdIbRbB8UZ9IabjKQayBnokkWC
sktpDb8uC/5q4vRuOxCjRr5IxBkoi7LnaLfxQBmrbzxT+A5bQ/qL0+DogQZFRsUfMJtC03kIFBNo
innD1U6H06kJQCKiA71e67NltVWHdcLzuLWXlveeCraz5YAokmdGIX0LfUw/XKMxO7H6g/TkPyVd
WKpPKkmTKmK/u54CvRTeMGeeXEgX7z1qrLdvf27J9/BqT93T8w+fZx6dTFzUojGHUfGQvTnBxjz/
l2TfEB7Ku9rgdaYdeoqTWjuMUigb+YDAM/jDgVvxpRLDtCStrPv9h09KrWTmbpkp53fKyLZk77eQ
RuGR089gIQ7fJHMo+pWp3s/UW5k0pNoOg9zPYR00/yOIihN35CAB46gMILahIaVIQxSU9ILbGtWJ
lwrEkFsBXd1MghNeQ8quFPtAKVL1JB4fh2lHgvBxmhmqAjYlklE3EOGfLfHGb266MVs4LHp7QEwG
If39kjZ3etmJCA0fNWEyJSTqXwNN7n+gC69hJp89OMMfU2koABv75JwV4JSsFk3fNqBRij3VDAo0
yjL5rKFLh5Kb/w3EEpcihRp7RCU0t9qNWgo/jrJ14gXVwF7nlxKPlhIFtdERZ9l5OAS0NcARr3XR
QnibZF5lO/4y+Q96PYV5rEl4UqedxQNe9CU4732pI8aiyjY43U1a9I5qip9OqztuHsyiRz49CG9j
jFKYUYRHSJ+qn3mrAwpsiUZTCmDafFhXzBQXq86R2/yR5MOVW84EkVTkdV4HWuCzJmja4mXtThYu
tA+kDC7t4c6wpq6c3Z1pFomlIlLgP03SFwZtXRsjSeKbSli35gdGBDfj2UN0QSP3aZj4ew+82ILt
gBU62NDV7mB81UF9DJarraBDMuWpGCCL9U8LTKqvII0QG3o4TLPJmnJpcHp+jDorI/oSR4pGpzdi
qRJPTkBBbuwgBQ8MhwFixKThZxRuGcOtSwKRnGxijCMB9P0WABorweD/jvgaUdEOc6KPdPiM5O1t
x7ID0Y/VhjR/jts6+LLsfbvkMbOn6G2yeYRtTyjh6Vx8Bjd6X+LivcWXeZglz4usfeY5xHKiz9ju
eJD5LB6B8zQtz7PldssnQpd3fdeT9KQwIcODlc1BBZs/w0k8Iwvy0kLOnpgZANFI3tBL3kpTbUPe
Kp9DFHYKeiUUnCFDnsRai8jVZuum7ySR67oDBhU9YtvU7whp7BjkpAIP7QyRNqqmN1QOhxCvHj5a
S+WlfiOCkicd2i/3AGSQ4rk5WGy8ahEBSHWBRjkYQdAOacQTYMJ9mojudFjok2iPpBt5n4VmjT3d
uiYn1v1HJO4ifS+bvcr1NnNdrBARA1V4g88EjTGpyb5uBcUSvVBCN4vpTG6Lt0Y0fBYyQHBKBl8k
hTbGzdhe5wowVobGmvhBRna2s9UITUwuo21DR+rdkA+YQh9HPpt67ARV/9zBr3v4tAS26QoZmA0n
yo0Q67Cp4+54/bOyIbtNW7g4PMhKcnnUUp1+bP4dxd5kpie0u1/jI6ddDRc/tAANDjZBdBINzndp
XCExrHihtiiKWuiZbqgGtfui3wnqYzVI+eXUNX8pOXIUBG26UA1QOTTqA2YgJMhsBF9uTl1SLDaI
DnaBzOzGBABWpBD6ErLUcNfhtnoqC5EGhbgng+/CltI5wLWfEki6evaXPF9voRtrXh2dO2PyM0yu
6Rpf9WvjkFHpAeskZYQrnJK3dmv+1+IJkxoVz9hl+IisRIbc7EjtDkB5aX1Ha3GtqjJGELAA5DaX
KsWxTaR2+iztMxrPKAbsv7Ny/N2TcNS4wMQ3RJZf4EqqrchtW5xnQCsUEMBT5vymbgdcwatWMXsA
NQSUD7uEf2Mkqp+btIfpaerY6xdwyHdCb9WiZnZcDJr+v3EFGEVKyItL/JTooKeEqJ+Li7nioJpy
1kygNMEhZ3zCkafrFLlynV0ZuPoMC8/1ix7CXPU0/auinE7GIr3IK3rpHlT9Bb4mR9Dn0of0pfrU
SyDstZw+/GYyyk0H2h3TPOwCpqkTMVDaEz8BoC+czQWfzAUI/fGMHgRpU21Zj8Jr1HFnAPT207jZ
EUBhEw0IwteZwVKxL5M83DbkOe9LxTi+/ZaA0irjeX88DGXwLSuw2mP6e45p6m8BNfM5L+AaBzX8
5ckSGEr8rsbwlieUWpw9aN8ZMT/4qI+0I8CnyrrC2Uas4D3PmiIeGM6H98E5MPHWL7g39FK9qMXm
2wgfXIaQCkk93oKa/Rzo1P3M/+mLjR5Qv8muFa+G7y30eJCvfEzUzgAx5HcanO1i4CHAMwyGpowW
q+5JGyGgNYE1lAy1DpQW95l5WrNBh6TuAuRWpOPqvoui1wPZJBSL8jQFOAHCg2SXpNM/cpsbJHRu
8IJuXOTMVIH29hH5gHRWGZEwdedPBjedcmE+jISPFOQ+HaWSfYuARdf6e30wcCMpz3W8uoFd5gq7
MenJ2YcVkPqYdg5jxIwMj4sIku0JqdRMUuQEU8pCBIR+KTAlPe58gLZelUFrlFYdDAlQEG3kAdDc
3jojUzGln0AcQwS8NQww42Vv5S1vjWZD+k/QEH6nHvKWdF/nkgbF4uCmX3xlL70plDoEEkFOuJ2c
lJ4qVKhpXYVcFRwpS7aQSYjhqXxKvMdWbW+JEsJ0xxzE+AdLlBFbqn9mmu3AQ3S+u1dKCpvUtxWm
6rTzyAFwP3jGSb9X9d3sOijh7zOY7VeG7f08ASbnJNHLNVk2FfSES43Tu3oK5MEsyCLD7l9CTFMD
ftFdxwcgwHvCSkW34Tl6svIjooAQDmXE8ettYJyTIMse1exRYbbkdnjb79+vyDCxLh85oid8PoOH
iPxyhrSHAThgDjIts+dxS7zJ0SdEnpjqhxqZjs4T5ChPp8IwS7aVebp1god7rW8oKv1B5xvvKLdj
WtWeXYb4GKcaYp7M2iwNUiS687pNscUeIu98LXlU09k34ozE98cGm1bKfPCS7lxQFozf2UD//7Cg
mmhj9pbK1g1tr/MsEhju2MBA0zwEbBxg2sRUN+tIP3vx4s5xa6mJrRY8QJiVq52LjYveGLPknmEv
o4T7dus9DLsIjkO0yv+bWWoRdDzzRxZcRRmwzGp0LnJso8n6gA42M5a4oFD6FMKZ2GuxOYZiBNTu
7sW9J5yy6NFwiHSQM9kmFnd7fZutIpV2DoATdR/6lC7crfE7rIKHhnI2IGX/b730aQhjei5GFv+A
hXAh03ct0JUuifO6BYI+0fL/oL9Tfpp/B79hs4K+oXnuuY2TjmLt7GUWkd7/B3IUlcVNii+9XSp2
bKidl6x69LFSoHAjF38OqciybHLoqm1T8YYsMoDvsMVaDXrZUsnC5OBNznQDR2czgKd1lzvoO89w
NL9Kphu+sLm9/X4DRvm3Fl+v8V5zvYRwbW5ardHQHGkXHjlZhgy2lkfnaF0Kw0vJFvS0glJdyMLv
Ex8Eh4pI1BRkFt14W8X1KvRjqq1F3CklbDGNKvMfLfGYqcqPwKe2wFLsMvB37InSBfIRUmBCXjQq
zCDqWlDqcHnTQQuwXdDRSpIL3KTQyT5vlFKf8K9taUtqspzGjhWaTGqfm117s986Y0PIQD4YKnHd
0gte1hFnDD1LKLI/yUNhLwO2mvDeGzRT2uTgcMYvF4UMC6gYGSMNnd6BHE0zd04vv3KMD+9NaMsu
q03lY8NB3BmqNhW8QDhGPlsVET9+Mgo8pW0b27NZ2ntYAfgn7GLflW1LOkqS9II9NrmH4S7JkTiu
Bndy26RdDdRJO2BJ5pPxYnBVtLz7K4sBuwmsUhW6E9Zd4YPXBPSQneX6ytD+FXRWVDZ+QHwXeCmA
m/Efie7NAYHCYEoSP46/AAn6TTBTZbgoRci9FVHmvH0MVgwpoKAGyWzwwEtUsRIskYdUIydBRd1U
DSnfh8ScNmNg0oz3QKTkh1Nbbt4kJiA7+wgcQyxtiYC+O3I0J4ZbuGFpDOaomEYfvot5KDXAoRfv
irswbG+Xnp73FJQg5fvH2toCkU31Q6lFbqhyTrpJVRxSLv/8IxuRDkae7gqfoWshHdT+PbUvFwcF
x2F7XidJFQYm7mlCUMrTMXZJTnqUCyFMCZhTiqdG5ZxcclCwOiBvDu0Qv8LADiHekG/SvVGnBt12
3MTD4SbI/Aii2RhRK3ZHWTNpDgYexAlauAhf7n+rDXsQGb9q9XHYYnMEt/zIhwEEi6VKmfPWcTGF
0ef7pMx7z5Xhpl2MrjU8qhB4VCD60THxMMpj4XdfnPPyOny+ma11SX3KGkYGUk7yAqvM2Xbt0KHw
KTePVR0V2NFmlzXVlOTqRC0dKePfFpumYI1m7OqbVo2Dz3aoUZpRfyapQ0LJNwQlrqmURfL9Wugn
0fGjGQ4o9vjhaX9tE1dXmuy+8PDt8M7qOkNXNTKGH7wDmUQrElE1Fg04aaXCr3tAbLmc/qatlFIN
1UzecoDBrhGTZWM7gozaWiFewatEjrUZf3rzrmBfhiKSHzIIXmc4C2Zxelw89wVUM1UHUWCvB2sy
m+s3gY5qY0069uBLkq7DtZVFo5Q3xLNpR5ekZ6NSKwDonaK10rXsyReBMjwNr5qGWP/v31E4okut
tu99lZo6JewvmjSOUPLvJDJF31srpisZjIP8K/dLH3W5Oz73OKLkhHHyyEdIGuMrH0cjxHkB5Taj
8aWIZIVs5yKpdCemHK4dsB0VS72vmS8gqX4NfrkI1jorgTbiPa//DMqxumzBh+plpBwAcl9I04Fo
XY4mnrO/3G8/4aVItRZrVRPHLO8PdSaNIrgE3Ijbf7RHiFlVZqdmcGHfbBySrXJDtRvuNSTZliaO
z4/d6rNf2zQSPn8VhgF9UyP9SE+0G5x2a50WCuBDk+pz/W3JxVg+4zNaftQuPy4sYUQrjWAVohWS
5bp72wWR7akuDgwQlQSAh3r0ycA33fS3jp98B0OMZZ7UMKccwERiyXOzDrWbP2vu6okMpA7I5Y41
57SzabFTo7X+xzE+z+AK5VLwNtA9xptYQANl1eLNAbkWFusWUk81AZz0bb4Ruh/fkOPzJnHntpbM
Nvgo+vzyGB6CX6qrpFF8X5nWcbT7HslP0kOKfPOmkh8zORfxdoL+ukVKKMuKZ4SjtLB8PUtuPdJN
6gyihpDVLjYD+X7rdMhUIfr3kMz0P8BzVok3r/p+dA4Z6vI7HfIx4qJyg54cyXYQua8DiZ6w0Vwu
KR4Maszy0gsn4Rovp48T+XW1G54+CqiXn+hdmpA0Nu/Pccj65e091bnsjBnvvaxXip30l8Tk6rcD
OawuBtASLeWb0ZI1mSMLk11TBLEjrkQWFr332W5eDQqZZUQMmipY43Vzm2+uSSruAuNCQsVwGQge
YeFFfoSyPVcEaK0pUTself8NX6HMS6AqQUwrOw/ra+XV9zbPm+JVKLO14bSiJtfRk9bO/nX2UIYE
H7aBBgewTUBP7qXpdTkQqD7LhrpgBfGXIh7W/7EDE//KGwDIq0IrH8NdJF5cqamo8FHEsOstrmvD
DNhcjEi1kd1y2B+EsluTwjjtklb8xUMczY1cXwr+juH8t13lU7qRtd0Udssdmrqdu0sHelLsz6dk
LgRF79AQZi45NmGF6x24RT8UvKHCxdJP254YGCu+mDpJgasJLaBPWohdN2An17c3oyJ5g1Tg5Rju
HR3u2676ZK1xcvXm879SYPtvEhrrg5yzTQr9gG5sCD9UXUhZVFRglon/pO+yrtprAgQIrroeRSHT
UD/M+z3H5ckPHIegLVnVsSwayNFCx+TZLEa1vmQESLSOdKUHQPrNL7sVVVkeVA/EqG4A7NtaM7Tt
ETD3Q4pRUJUvEFzlX/rbgn4a/I3knjHASzWpnUkqKXOAh5+J04CXRwuUaaBA93yVGCbm7lpMGxkz
BI68f3SxpyNm7h2CHGg0r6cStq4BOdZa4ZRXFH2esdB6+5+tqlfMzaNPVPuBi2W1OYLnWL5L3Cam
OpsnSpDNn6T/EWLohWjWjZemq4SjufoZyFZgGUioNOJn7Qz5D3lIDTRy0Ds40cuFmpUaCLvr7c1f
9JUYZktBMqOP1xPqQ52jSIJyDpNKlPivkdz6CJKjjTh2ej42wdQVYv63OQPxlEjivpOr27Ho9KuO
g4ryH2zGR0BEryw9THGP9tUCNxPn2NxzzC3dbs4/3bDcMyYUb2YHn2+vykwNLC9KwQlv+wVrruDk
dt6BKYDaZrJeooMiF1aItv0DkYsZ3+6KMg+7OZ3YwivWvImRV1OHeONOUn+Qaoxaw1beB3hGQbYu
oyoVHa2/sCDGS0l5RAl1Ur9BVyZl0sObR8lL6f7KDZKZUA/16kZQ/JkZJrI8eXnmX1A7KjqRIBDY
BFBs6aLhc/evp00Hin3lATOABY3pkU4DGonE4KmknRKZoLqwn0Oq+R+GSaVizD746oXH2/JgrCHO
+z2u3NV9XHBsgPizOvI9QAcYt9XYxGzxAGGEd38JODnh9cKNwItOvyG+4Hvg8TbLRHJhIyr0ITX2
E5JPVSXzEKRGfVs1eJWPmLvOA+jjlHNzwCjWvqk8WIXagoIRLt0rpTgw6oUBcK3BP0uzr7OU/39/
Pd8r2qMQPDlI1d2LHjThsYRQgVufZ++fHN+v1q1hC0be/fSYKcIGteSr+zieHhsv7ROOXnC1GeIz
OQZwOZS2A+JRqXv6vNBd1IDVNP1+8+7kUSEKRIVR0ukdO9ydSCjP0Zya/lvAxcuDeoMdlDYnmCUQ
F4HyFP01CNGovcMH61ss39Gy7cUflE5ZXLo9yfRHTaTNdYJB4lCGgGuHKwtnla4DOgVLMZRyTyaT
Ovs/oXm8zt3sk2DMbOkR3i1Pg8ivg5pVhW2uN7PfKm3CSiw3d6HW6I1CfYPbMz6jVb6txuHxBnHn
cxBGWABZAzKhShX95PlYLZu5JNcJQyLxqyrNlErk016INSjNED/i2LbfXulCf5eBzhEuEDOEC8mv
HJwcUIrdenariin/i7940nlXoZNnR2Td3sA6/cfbnNrZ0wXraTKB37JullvQY7ZqtuqKNFwm3xDN
QXwgMG1IFVHMeNtn+fwJe7Uf4mOjmjrqBePnxifDOlPFGg94574ICaV9xYNL3PoZDGNdzsMS2Dr1
sN/6WIuXynywG9rOdc3q9d6y6SffUmh9WP2MiBA7bpy9AeReKRLsEf6HQcSGaFfbeoIvmF+Tt0hK
FPVqL6dzjJb9VVC6DJ2Ceb3gs3A49vB3Ii2levM0mQMhGTNnbtRG3JXAkeGPTK/uHDlqYALu2pan
fyV3YjjBsxR7k43vws6n1bpAWHfhbYMPv8RKQKV1onHNTEQEAsF0AyMc9I5Y70iPwGUU/RqZPHC8
c7jRjbCWDN8+UquYUsp3hFJZCIozGNepkwtM1kwvm8t+XLDSBf+0eC5EvH3eY8YXxFYEFx2a3sst
etSkLMoQpuDb9AjAfzFDc8mPwXV+/IKqITHs/F+NK/X74T3RRnwONjbemGpFi+G+Qg9YXSSFnWeZ
EIOhgTaq/vndor5V1FseDZxXkcbvC/0w5rtNf342qtoBUpZ+j29NC18waVxhScocF+npjuexYcrB
i1fdkTGdKxsSSnupAKcj9DPFQhu/hRdCI6Z+NwopvLo4DftGnH0lm7mB3rCvakEtcUcVgF8mY4Yf
I+xvVhGJG9NMovuc+CnBtLZGx95PWsjrSe5WvvA7Ol9kxDl7sizYYXTHQOUlbGf1PLttm0PTQMu5
bI/9xslyR47mJ6CXxL0xpBql0QHT/4iSG00slggOq3iGVusAE1pgEE0qSjdMuW8e8zkMDJINAfbP
dVF1BMrE1N+AzVzX5KpHKW96BLolnAv3I16iAynuxGWigqR+GkH6E9MYkvJJRKVhjAlSVh2mYMPU
QOzIp1enFRb+8tNHrfqS/dK/WEK2Hi25z/ItfOr9gm4JCQXoA9v/ZTAKkE9wfmP4Cm7besDyKUCj
5FnjDsQOg89D0dyegK5uYWg0SQmzJN1Z5OVAqc3wDpUGNpEdcrzTzmd0eaSncxD6hgkaMUPjhpqu
lby3m6ryAW/lurHsBrS1Jv6bnB8k7dzXvW6U6Tq/DNY1NQrFt9+gqONyxU78zhf0hwc5PPja6lpJ
BVSsQesaEsw5Zhv8v7faYSCs622iZnxmtJ4+YJAm1ewqluW768bPD+nCfb35kqoM1XcfWCQIhI5B
qqw5XW8bzYM95wr7nc2zKuoSBMcCmsGCSSVmL8DwnYdABkntEuTKnQ51iKkb1ry5W+oYA27gPCv+
BstJjaSyOLBw9XLfAPlVpF15ZrwkNnioWLmTdShGLUWT1hdBxpbFb3B1lzFCdJE/+E6rTSC/626T
NNFE63FO4RkfyifukfPe8m33fi+kQoq9qVXS8fXEOLp9b2Wk2YpS3fi5m2z0osKNJR/xmAWKOnZr
J523WMIJQMwM1RxEi/yB3qmNB1QMU9fV2fkBaO2fS9wqhrRsHYVWvj18Z0x17b6gtHASBEPTPJ6c
U3z8xa6NZWxQThuKAu+8Yk9lapy3pL1Z+aEm9a1k2gMhvfd6auWwAszpn6xCXU03jLengzcZyxaI
d5nCfnk3ELrq0G1xP/JO2RXczWWQ9C+1OF83JArsbbPKF+EAUT3KpK9L46eFuvPmdj8mMJAAGwhC
5kiHMWwK0/B15DijJaHp+7MIiPeOHHT8qQYxJEAM56bimVS4tlE4dmw9tAv4/cs/VwLkmo5xskLc
Wil5ngIHNBqor8XOwnRBKtxNgV/A2JL4YOJEuYYZhqMfhGKtq6t3f/djtPJrA3/k4SShND/0efbw
0xOEqvi7u48o7mU5SVgcPTsSmC4PPBJxzuqFhUzyHk6ucM2AwbSH/8fwG7shS8ss4wUKsrtc+0EO
WndBqqmjK9+nX/DbN4T4jsMkhBgosfNC2m/ZMfyvYP5D5/YmqsI5YbiteV96qWSuWF/Lbhx/rM52
nRRGzZS4rgCAPgE5DRauMjZa3DnhZYGFFIDyCBQTRcnjt1kWa3kOnofuwsV4DuUeT/d+H9H/9s4f
Fl5c7cx7X6vRy6srQi2dUl4Q2GECl1gFUF+V7b8a5gi3Zn6WZF6OtkPpd4dFOo0tOd4qSk1LA0OE
Wpoio550PzC786wNcPCwbshsgjAVGWTCwBeX8nyT1w7MFSV9zH4prgy++H/5f0o9AYn79dWC13Tx
t17e78M3MAS1GjmFYUrc9wZsCNkYpuFMeaWjEjo4bqxrpZ2ol7dSkWO5sYjvTx4Q5MLw5M0eEcAG
KRA0ceUX+4Cib7LHP3xTWLxleukqJ9NpId94080X9JsHBGNzTR2ydgzgmNo8T2vkHa1ooqTC1vKC
rM3M3QWzvayLgANS0sdFaMIhbN0DRj+8ndTuUmEqU4lyxDKnYGnhRK4LsZa/KibIGw6XsOJz6AUb
w+utVXMsq8VryD2QI7xDm9nHhg//QdtDCv9b9hU3oZ63Y7VbC/DXRgTu2UzWIq7NUzHiuUlNlxkI
PPgZVYVdLyIFuOnTvaajzY93DQ4QXZ2LDhKfEmH7VRlHOQa4M5MqDw5VYT3zcg++jAisKFFltuIA
NsbUm70GodE4qeKf/vG1pgrqZEEqX9kdjdQmcWq7F3Zo+XPDaIwEbKVyvkdLXUfiZ25p7XfsGJyh
9JPgcBWqIJEn/u0uQPvWsYaajbsrTtIdIcRcJUOvYG8K1tfgESM0D4sOQesi05pFoTX//6ybhTG8
t86Xd5y/2EwdyhRm5PMdXyS9qIFF8+VuDsZxDu1AEhlGmq+OG7esJL2V7EZRTJEVDxEOtGsUWvnQ
l3W5IduqtRBDWZa0mP2Fm7xq/L/jTWd16qVaHpIYytlyDVBVntqEznKEPUPhGTT6QvZ1lW+j83np
V9eBUskC9T9TdaVDKrP9kIBO9l7SAXvccNMRbD/QjqgRrPGy/M4O5ThN+o9iDy2rIPI+9NHMxCUH
q6fyuc6Up9WCdHrhntWXiEwQJo94XrN83jYNbRkpvp3fn68oOdwrwFt8if+hjVpVG1pw6uaC8Mh3
0K+5gm/ouo6U6Co2OPNI0eJAuH2+TtNWZ/sc43pcbjd/NoITWRmKAIZB8Z8Vg0Vasf7FIqbmS1O5
bQCNxKb2665WakrMnk6jL6fmwR+gmgXVDl6kk+D815WcayD6qZPMxqyIbkq5lxznesD2Sb1gm3hu
t1jr/QnkGX2shhS+5ePIpXffywhogGqXtakkUyVX/dN/LOctC8qxKH5yk4+lps4RYyx5ny+kpvka
z0JpA/D34LTJqzno1oA1oQjiHTrFA/VammiR2TqbOD1KUfG45xplgW5NscSqvfe7kNESdkqkfYZT
xIS8lKNbk7WhLIFMrpPWpxImMJDk7DA8RF417WmUUmhvGBXy4A4FTmyeW7NQCzcI99HqRI0LWBNA
R8c1nd5UOhsDEwQnK+0WZQzyN6rU4yST4M57d6caVlD+AMLoUEnqF1hQjWzX/txMn/8mXeFuqMFY
IK3e9gYk61MDP3aYvwfSqaxiIxP0yVe6qXYgMdKo2azQWY/5wypvNGGb0HavHsisB2FQIzI/x8Hx
2tKFfaq5ZC/axEaOgmzJnOKc12ycKPjkDjsz8LxL79jiBBjhxaq7OscKjZ75uC1FDFW7gDXlj2Za
AbJloAOkaEeT/6zid1btulhLV0TNLgr7WyOfZGVojSIiGhKfb6bs2t13W9seyY8vaZhe18JWRc7Y
gZcpnUkTcGgcTiETpML9sSYJaqE8tJQ1BcNp7jHD+88+BLQWeCphRTdxJCADjSVgYHpnUjd3I8dT
227OVIBb0zFEJrQJm+cqsxcMbmbucmrmaxm4oz4msZmVKlHHy9BqS2eKANYh5E4rYVIbzumLkUDi
SelG5nTbULKtzxbNqSapbNNp9POIkbKLcR1xlsFm4bh2WUNbM2u0mUSIolRyJqIGwLh9CrmjohxJ
EKCC/XXlmx++dilcdYvh9sY3SVFIyc6DW5cNbCNtzhnKrCmCPmoDvX38N5R1PUQViX9RN5Rlbss/
Z47S6mdkUwfx5jdbuUrXGkPt9LBpdxiCUAeXRv/IPXq89+Ec+HH/R3Q3BH1oF8kMlwdw3Tc/W5jk
f1DCgC5zTfZPN62jrljgAjtGs+2yvzTq0VxDwZZSrKqt5om1njn9Epd6o/Dtkg8iErJDRsjqlijw
/7AnkPQfc92JdBXBU1RFC7LuB3TPo3qKf/l1z6aiKQTSCRN0Nugr9lbST7r1DKQKWMjt3tC+djGN
ltBsd75vziUAyeXXbc+MtnI0ymbyYc86TKCD7X6iehrYAHn2Fc2d0G+OXggnupOCwGemn4e/RZnO
yAWdII6NW78lzCE60vg67uSqlHo4I4E4E96zaEDN6oZQLKpJCoX5TZQOBixtUWvZ4HokjzjA/bXg
Z6q5LmKEwly/F3odbUgxLd1kRLzfMjhvca9kpTP3H6rV176Ac03NhcF2jBo2w2LMph5HvZVAJboJ
AvudyntHSbC6euhkyTNo7uLyjeAg6Kn977MEM6+xJkabCo6UfRhUNY6N+4i3w8+nCWgNign95mF4
AdiVZfN5BFU1kmPlZhTtHJFodi4ZROSYt6GvxlHI2krfgTSuHkNP3RkB/TVAMjpcBflwvnIqkyfV
oppzUooNnEm7dRBXzKATRc3+V2hwoe0J6TYx9NobQZnqdrxI9QSXxFWU/arOWCvVAL4UrYMbCcDT
HGN1iOMrllg49i3oGLktuLiWLf/MAik76Su5FLfno68SA5E9l1/FxquxYkoMJjAQctyb4D7kQxV/
KsW6gUzbOkuKd6H9Yx+pBbpuWxd3PVzHcVasnFw8o9kKNrxc4mBSQPdULYCBwxEkmVlLfCHhk+Wa
jvDj2I5aBZdwQAGYJfKLnr8UfxqS+kZLXBfKwfoNzq/h2eYrwlxulG0s5e7plkJu6gh3q9satmMW
JIeRHRrZffk4O/YeeDIxzZcOZy/VrthWY+dDtfturQCsVvRRmbibrZeHPBZcqu3E49BIgGDY8cdt
cbzyieuN05Fb3fAwHt9lSFUKonO7tZuo/BHza4rmQrme+qAniHAQMmJsevnmUUkqFpcQu5ZKBU22
NhTLOywaFm48WxbYYvvjtCzZBvDRUbZE3mhpY7kpmYuMxoH6VgIWEuCgGKl4n6h1I5TDJiZiE6f5
XwVsobVw3fS95XSJCOovg3pBSejIfjy/2tPPvhVUS6TzahBoulRD4Zz+h4OauGPU/ahQtwTpokHY
C9GlfobXZYplijO6PT7aTtpVWQpe0PafAKXYbkZO4SsGg/OBaKSLkkj8lrh8fvUwrWCyywtobdWS
R+W4nHnJKgPmWbJtuvdURdj7cH/qGWOSSArTqWzwmUSsLTDU2I07fLKgKF3pvodY1uUkQMrxp1gX
ji8XwO/8AOlBFN3cZ+r8nZl6Lty1dcTkssO6ojVMTYgheouDbAtwt+KqqKD6WQjavgm6J+06KaNh
ytNP1OJ+M8Ap8rCUE69ooJwuC44hlwro7gUaweZ+3k6VboGFxe18Fwit8EvFTM7SVHTivZipY9JI
KJbKpZ8lIjcvPCIB3eIhIvWi2PkhqN7IrNsJASwzGkSsYOiJ0B1BwFymFSNdOgxA+cFZRxe05jq0
dO/WHLlE5tpaa5n+l3jb2wD3gPama+WR84RDacf0sUFW2XnSKkATXV9ilh6PCXLCd1M78CDWBVJK
aCTdK5iEC3lv1bCqr0LIshHSqZ+vQu/EI8mb6AfN3GNFDqxeuQtcvzNg7XDcZJ0f5L1xZggJAyzZ
XCOfCSoZBbiddZqabxj3hE1m7gnAkybzxJ8dz/6ZRQqE57aCydesBFsp56wADrTJbbbXLsg7IOY+
BgN+iPtbRtfrotv7eB35+z36WBxWn5MqqaPHlYopqPDn2scwll3oJ2ygsgYuvXpIMpY0K52Dd6G5
3m3kfNKPVl3+JTgdapmbCd+5IXOSYmkVT1F35/7t4SiKk1HdUrTZz6RgIWkRlA6dXFiPhrztVUij
2extHCvg0z1vMBbrUQ3UDewJLsca9cRGE0ScbkIeXUtrpdyLCSIfgWCMOqFqURvrMqjHthlgDBY8
duzwaAAsSJDXTXXW0rBnC9Ul+Y6aIr8D+MLV/E3918kKxNBIsso9yWmYUMJTGPhgBXRO4RgzmGF2
r0Kw2T4Nwidqu1Cbp+kz+pAtfvN+GnOSeuN2ZCYAkxqOw1HsqTm+RAhsAQINfKXszoUN+2XFmV6z
QybrzpC6bYCByHNP+oqjyjwu6ohwY9EkTFKPs6Cbtkf25eaTlEJjMhEwA7CcT4DZhMNfn8+UhJ5G
UEvU/x6cDQRrC3ghxCt3JFcOwtSgRgKVxrhWZeMcIJirnmDyLVdnkFo6mRUQlKa0TUTPNQyonfAp
1AOvTQDwCPRkGQUH/bSy/nPkizZmJwUW02P7RF/Iq8GTnAQctFBBr0jS5SYdynaOVQl6UyqiY/1G
uEG0RYe7fBpR/tc510o9CT9e5w6nno/rriqrhWe5e7M58CZglDTEGLipkpsVXbTyHIahPYxt5H5U
cmgoz+06+x0eAvfP4gPL/koYLSnSpuGg6B6VfKQtv7C+qGqAaHDacW+L+SE3N8VGuI40AUVuynoO
p3uYh+/iQTAzqvK1tAns7Q8cgVxuPLh0NTjz5hXz+WIlO46BXoMPTv0RDjWhhAiZhxlAIDqHC9f+
w96VUfvqSPONYxtFxgFLdOmXiBLUD25A8sfWnK7WFH+/GA0qVwMgR8MJA5iUgQTqvKc7hmi8ToOg
SjfK1O7NXoylrZxWZQ8YnLU5W4KPUFJcMqSF9lq7puL6Al4jZL5xYohHiSrhP3D453ZS74QJ3AOn
51PcF1Mi8+u+SU9faFwNUc3QQ5cSygwEm4F/fwmrlyaZgLUzzbS1PjZBiLrPTzItyQKk1DFIe168
X02jIMmYq7WikLrA+zbpC5A/ZncVVFL95k4fQ86oq6pvry4g5AXOjKaGLh0w+oQsR5VK3gxcykAN
2ajB3oxfccDvL6LvTAuWXkAQ0a0uDctEX++mJ5hSNa8/NRkgq8F7W18XPh78afWJs9809cUgClTy
X06BcIzy4orbJEEvoHnkrz0bIFuIy1/Pn6chj0rVF7tpcQBDBpgKBidKESgazLX4RaHijgjKuvzZ
lnFu1ECb361zoo9CmqH+u9ClMXydaZzLXzq5ysrSEBMSsVu5M6TYiPSFN8nkNMpch5wf1iC9O0q4
Q3YRlp14W7NIwL4/lK4ruHjcymYSlT3bfMjMvvg7ezbpEseVHfdNCIA+l8UDL6sdMODXSdOYZDqz
olruAjWjFNn7sa4n9GDY/ewForVDfRgOOQe8UaRqJN9S8ItIZWTodKdl4pAP6E81jSybjSVR8MP6
y4AFnd2bw4YMzN8J86rp4WIq+0tlkvGx1l1IbDfbjOwukhZmzIjptb20Gd5inzrWffR6czDdddw3
ozMWB7jw4PZ7c+JZ+f+LLHq56cMwYKr9Rs6ZJEM2hwX1/qwAPZiF1C0qaD9jBIdfchm27C+xN+lt
oygk4/pW+hMQvSUroV4HLgticrlhoCHtaqG8mdItJhqPI1F8ECGexEr/wLJFQrbHkwMtWnTzZKj7
zalnBqmWXXb4KvDTMrB/AH+d9h4IfyViTMMBNG+DAWagyaTgCoRDUfsDqVpc6pIu+PdutHvx0fvw
kdEMaz7NihK9maqnfJETJGDzUPjehWEDamhyOyp2HhJNe7ec8HnRUxQGhry9p6tiPnSultahqKC7
ej5lJybS5DNqI20SVpap2SwgTBiBcDEzn586VFMaPAHvFbSwQBkhgpIRxCQeM0G41mL4duSJH1nz
h2yqiCPmbjYpM+ghaucUkO0Q2llxG609AYNzio7+JwUUcoLD63BHt5cvw4oJAz0dr5Ux7prMWSNK
Vf1tvYrgW+lLwl0XjHvs6LfmmAcF61PjLVe2auU4ClM3tC4Dy5nvvZHnfB6W038UigBH/aZ6oW1D
4eK+6qjJX1bvkXsMlDqk/HUGabkvTCY7+pUaj8AnXnqfXYlWm8QRHvEctKWyC2wpFM0C87X3OvDG
0TKwMpJBV3ZRK5KOUdevoGN3eTzN4Vr1cquBfuW4dKgB4HgysCSEvQc5uebpyi/kJHp23iw09xuU
h8EiRrxF77XVrelufk660oZINSzVvXxl5MfIT3MXqGXFvXL0F/aeZuuoB/A5N3hFMn7OUwt1pkXp
YF9oThuxzlOk2ry3bERMtBzMhSQf7tcMhOfJXz9sWGA1GzYRoB1HWO9zY3Bwd//e3Obb+ZHCSC0N
pJQzcCvtc1EMAWFzK5jZS5KlO+GmmgCDmLVUQsPqIujZQr9RGkUHhXVAERJpynXOLsAZ8oxpAS/u
t8siridjVbF3wtMN+EAd9HmEmaxeHK0Yxc0BOoetK/ySjsVX4P8rQuORrJWtkLAw2F5Uex5QwAeB
fAGzjv2vhkp6tWnVYUgJV+pojr1Q+TjFmYqP6KMh02rWiDwmGNR58kLWWAD9IBLWcfc9kNmsaz0M
4AD4WNhruVrgcEv+0ADJ0YUCyEu/xI2vA43zP9/fd7pi6+2abots1Ya0ElYWCkl4ycnHAAxNMN+6
jXd3icy2dVcTY93Qboo+8wXa/GGhFzTrod9Tba8WFBLXVmg0HYv0x4zvzneYXeIQYB1chZAADaJr
jF2hCdizZemZcl1qaCehWDIaJONlQnDYjMs20giPc7XllL7fKdM3c5EkKpJjwJ138/NDl3mnb4bd
kO8gqCl/jCBAWvhClXThsJaUdzxCUY/2TS0BodzhFEJwbornVUXN/ZZ0yhy/vtf/HpUpVUMeiITN
KMvWwau0mGSSP+Het+eifB2tQLuzrwcvx0n17yA8aVbF2pdkefDlhJpfnud6swE4r3xmG6ywNOHY
HCiqZRCCcg9YpCD3ynZ5P55viR28wxIYec72tREa/pSmrHSmJSCRkBakMpxFLGAcS89Di9HDUwVh
23Ff/2YY0gRJSlEVd90TOIZVHbq52Ji8zf8LJryhSWM1rP1JreIqSQmoHgoG6hE8F+5PeM+yrKZ7
4N16fWw5Mqh3jT2y6wA2GlTcx9b+u4Q/Y4JHdivx+5rByw9LtCbsVNwmlA2nOJOlLA/JbrkoEE2z
fRccVtZ84VlgjeZrB51tYxCiBoLgghSfdqbOdG/ZI2BRA3NHKUwFNJEruBiFH83qMSaPg47Cu1cq
1QKjFi+hD0ARdRPCMii5JWBF7tYNfdwqc5C4WTdIV5LwtbzYiLDNg5x2ald9Ay1yLyM9NMaOBef/
Q20IoE7SrQYVA2AvajpGMfpD5FXkQ50O7uxsR/dE8RAF5mDfNnV9QoQ3DR6Z1li5Ic47q4vOtpS9
tlFBwoXbCfM0ZLt+GviT8WMoEGvyleUg+qCzjLsF0jya1a5ip3jdB/BX1MZFl7O5XniSq/KyoN/n
MxDy3Gp9YVFwagrSc7tfUcaULRU3JPcQJem0bf/+j57ojc2ejG9D2YKGIQtnrpgSEm/yQlAZgmov
qKrk5jQhvzUUm4x3L+lXy2AtJMh3GJSZqtZyq6sZQYld4ka8RBqUPn37I86ukJ/Bm/S5Qec+ikkq
427XPPC/exHLt0k5H/Cuw9t7KlbtjCB91DHMDrwxLBigCGq/PKuqHYt1N30e9IlUlqApsEi25wa2
iHE/6AuBHe1P6uSQZo137Hl5FcQqXHJqQ9mGso0+Rm2yY9XFT89XbcveQP/aq5XA+ulRI0oG1mZN
Ob9Kfi6wCeM4zJddP/4PFQsUmADW+9cYSxTfxL8qjD2Hs5xMI3S5VRpS50AFMHs6Xk0S4nVvYgZy
vGGqHDsQRORxfeSaixVElmGfoophj3C2VFdjEwi9jWaqoOak+4ZPc4oL6/6d98gLoDUk4+O5RY0U
R7hUGQYJcW17xgN7+IEEeSSAHZMylJUdCGxet0bqMYAFTgJOD6zF8vfw4G5hEIw58ZXHPpP+Fz7z
swNWNElpOJsPD5JKnfFqFaoG+5LdOm1hU4tSMxX8esZ0TuC67C/xPxXMT6+J4DUKXOMDvTQIHF83
ZuJmeEXWuhWgrO6wNVnWAhqZ/MUkBmTIW+cvEGj4v0tuvWbnmh9JEauG3gVfSQ5bIV/SooDWgAna
jLhNqEKpH22o9MdJ2KzIENKMqn5v+RgWYYFcROMGBtX5PKqIYMAiDaWRybtN9RhQ0YbiOjSekuOh
Gxu6Dc76Yyfe/QT9iDE4LkxpwBAI7E8yAXqEyWSGdqhxzMeL/6e6Kd4uZSlYmfkXcaugMDnIcpHc
ufc+sF1MdE9fo1FWMpTklIZ0JnNcLo7cUwnDnYEBP0cFaK+fLTsnQPzB+BQq0zz41IObTqS4IaUP
Heq8qS1rdzDSrJ5TRDfJynpdf7Tj1VU82lC1mgdAC/L1FhU22N2NSonwchtFLBiOdIt7cX/+ELKe
QHQxD27n2t8+aDnhFVQ7Mzurzuitve2NSaGd8y9CohEv1BtF8fj/5kd0dchz5oiowUwMvss8nP4a
X4ysQ12QO3hE51HRR0vM0T08zGJMEwNe6T2BqOCCvyQPr6gNEsCvPphOEISWIiCdUrSvcx7a16Uq
BYuEXqNRhGxcHiMOU6xj0G1JDsnzSUd73inskXbsW1SIPJZYUSxe7senCXbXkcePv9hUMRtTHuiA
PbZ89RQByoLSQmFfi1bGzf8Gwr1HBa/oOVQDa2sAgpherbinQQ89qjgZUi2bw7N/jD4WacVeroxB
kTWGz86BAy4suFP981VWz9scfI3ZXf5qYBOYT0h8DiNdCig6Bi6cwym0yDF455nj9NMic8k0admF
w9OGEoipcUE6LbJ+Gxi48cq5gz2XKwSpfgnRNw1ARM+I/FV+vhd7aPZlnRkrJ9ZI8sUs8/6oixw7
HDZ+GwmyFdEaPtihP4jwMW0C0FbU9jvKtaJKhv4c2D1Z7aOejJ1pOWnfXIduHahddrFqeyIRa6nU
g9U72rqvhN6tn+4xErHzBiEBdZ9Gh9E2t+8M9mkFmz1lyELA7xQ+CAZAnQy/O/QHy4tIGRmrwmYm
YfFHJLZSb56mrwoWn6w8lAWO7+Zi2N3F/goWJT/72aWSB1eyyBovVMI50J4z3M0o97T2T+6Q1+jM
RgPbeD3XQxxqTKIBfyuv8VpfqTyiiPQAXgU4vsZ4oTL/qT/XHFFU8gxQgA2K+8+mgyxOCVeeLkhv
cbAWADu+c+nMZqfZjL2d1XnZXYjCKQFFnGt/LBvqT9nMB0hLyFMHCKiW4VT3ZuforuiLi8/To+A4
3tz4L131o4712Bcg2bqHrFME2j/Fq/zP0sNnx9GU8rVErFGoZ0N4sKbtI352qBEwN1HcYyXcVmWX
mGX8AKllX5PoGI6Zn4dHZ+vtYt3mFwDkW5GnMT13aDIgkEgeGG+l9pv0tCx0kP7XBjuzB2L1uCYU
KFde2MbSyBoZ7vo8L0+ngaNFcduV9o0GwnKR6fmgoZmZIQBCqZHb7vhC6PwFJBM2BDrroI8Bvezm
d4agLzClcohOh/zM5bW9yTOlOBzPe14M5osD9lwXvPnEJ8X6fiAEj7xdzbKzFdr/poV9z1QZB1nK
k7ugX6s4v1kLYjAytRIhv49lMO244XWx8omb04s0WAEA/hdxiim7y/po01ES4PaZMCf2axKyhslO
Lw3rK5fLlUekCMXYAfEP49K0gwoNj+UR8Vw7631v/N4Yy0D9bcNsHh1tRbQyerrFnPX4K9+IhWek
JFSBhf/ReQUWIFaJBsP6ltahMHDgGzlhQyfVTElaD1ahqbmwoRm9jndKXJn2NL3FkMhAyGIw9Haj
8vMlyMBViJSaxjtM6pJ3hHYjjVpUXc3vNC9S6O0AHdT0phxTcZXqd8OMSLNB0MJ/Gsxyk4qLrJH6
dtq5jcClbhuSqU0xEopbxvfUlxfrogG+6UjMOflGD+6yrrE/bCamdT+xlanadPBZcv0x1jwGhldS
EihnXV653W91QCeY/oCnVtEt/QsIwotJPUZmSbHJwCKHVJK48ckxFqQgwL4P37wM6dq7wgJkm9Dd
EG5E0dTrlqGHgwajhyK/U9PNuVVEo5PjFFrzZrbXIP6cGUSjBtZQY2jJXnazQIsanUkn8LBgnUgI
Po9iLykJ8bYRCtOnYb0dX5lQD8VwGZQOJZVHn2tTlBrknjXzTwaUbsb6EdjmAgSSMJR8NSHX6oXi
ezHlRwvWYo+Mqu503b9+OZuucoJl7rKFWR/2GkK8ML+jdwgF/ZtsREXZ4D+5usB7EmyIYkMX5vQ4
7IUe16m2SX+a3rK/q6W3/1n2CWZpPw1Jb6k+usFvL/vjWvHCddljmx9j4VOpErXW7EPfzmSPPdTJ
KRSABNxK21jeSn4FZnx7v0hk37XoaU2WR3Slwn9tdnR2pqrPL8ezd6KPs1YSwS3ItWqMVKlj4XO4
9JX0PFqOPch2UJlTMqTbcKYYCtAdzjS3i1+8JbqyOjSicMRfX+nlmitr3GPG8G939KWm8ZaE6iyq
6ox8PlVx7v9pquz7PQtRS+P1MaTtZRUGsTCB2rhMj+kYB1J61M7tWSElVSREnK142TuzIk2zfixJ
7fYTpUX0cK+4dWb9Avood1IQZk+dx6A/3yJO1fiplwjgubN/Efls0fcK/PkhYi09bPxoQ5KWGX9e
iJBl6/IhYHH+Y+k/wvkf6WC4pk6lfhlfho+1bQFiqZsnempQY7+r1p5zvgpq35mp1gdAmkA//hQF
TMALT3qMo+0TdWrjtOEoV6bWRUZSnAQDJYweTbKMDUbPXvk8ixobmAI25KHFdvE68KFpqrQK7giW
11k3pYzhMCEkfWe0eUnGljnA15sBs/VynYlL2QMQnjBgSjIzNscVh5VUmCc5djPsSMzqjYzubTos
o0PEwz13QLulvjCniO5xF0qBN8pgKCFI+2JyZUxU+wCNSkCUlmkw7o/1Bl52EC88B8ouCpr0SzQr
1BBfDWg6AvS0OKGDMLP/B3PCPFd8GD9xizNv0xf9PSqI9mBw5akz5zsgY8yY1m34MWwwJKCvb64j
6vht1jj+EK+0OrVTRfoQRWadx09BKpsCeaOFKou2FGwTPNSeimsW/qj1Upf7tXwH+JALerZ5YSlK
0zAvun1dQY5mcUBHQFqGISw0XtTm9Q7V9WED8Hc8RJrfpEdu6jQ5gSO1cPXIye8vrguqIe6eOrBK
cQY0ItIu2Az+GVuAFzysmrC3H7PrdEDjeV8fHGbrSYbCiFn0MQR4OLFq+xVWWjU33EFx1jTIe6KK
wZ3JgBWohsb8i7PoKAA1lVYshWvLVtyoTM5uZaYVSkAyjV4wp9c6kBDrDlr63EoirtY/1vCLPF5B
c+emd23gPdIxxrAXL++IYRFd2U7v1VxNz0G5A032ULRFYdFH+IE5DuMlq6BZEgN9ivxGCk4RYs60
N5AmcDmxBTm0ZMRBNPKGd5D8bL9hrmMRxABiMP0qDvxKIKqq4Iy929U4QUoj+CpbrI9OuZSU5Ez0
H/1sPuPy8pEekBQpgu6kYKGNUhaXUVK7J+TWGAEGrfoSi4dP8mCgpJG09NdE2x0+LUpo0bqgSgkn
zBXSVY5dlj9YdcL9fB7TcsftsF4285g3U6LlIdijziCVpTsy01cUMzxBucQhQUIK24w+U1njPnNT
d9ROnmxs2wVXBbBarM2dTETdu4ORrdNV7P88xAdxp5tugsrKXpOgwK+WXWDN+IKPF8RKP/vaeykF
mXhj8MZutlbPNSu8rI9ncH0tdMXQXs8/LyZNLGW4Fk4fne9vqsJ+vnJYOGr0ekGTQJ3qXrEqo+EX
cqDFBJwcKGUSl8mCQusEU2eizpPlKQhZtJOWOpFydL6Tbu//uvXSXIPkLCTKAyS8jhr4Z9Du7gS9
cH2ihKrGu01UFKbILfJKNlvuBKFT4lfxfbX2nnQiA1UeXramBXqr1QuMZSD2Q03YesrID9MYI8I+
TE934Ej2Ci7cxlx6MbTtFUwH2AK6MMbA6dbqIXiVFbKCa7vXRHyOImsd64MNsZRXJOsq7q3uH5BF
R6Dlm7AgyHBZIYUFZLDfouu2aL97ou3Xndv3H2bikxAiDVJRU7agD1qrdYv81heaIxOMZMkSDZyv
9ChD7XckQX7+pn3ykTn1t6Y/SQgP0CvJN/crk7ck19S/9egHpK1NfeUnTDtG/e2jaijTStyBZvr/
3Rk2EIJQN0XEhMzMdi9kTs3y8YDi/qlfGilIMqGVh9AwcF0RC2ZMRS2fxcWWtTwgWxNKiDuP1pS+
HM3YnQPg695Wk/2BgJZeS72WcymHxJFrTd5B8qqMwJskOnPwKyCm8hc41Yur3SubmKt6LIbXt3vP
TggsFYicu9OKTj8SN6/Y00FTsnowsBUU2FNrhVumVVhF2kP5kOOi+ZMrRiLG1GJnJn/u/kO9+zm4
9wrfEfb1NJH9k84eSOv8A4gCiA9nZaOis01De0cpH+nERoriYx9300hw3BftScMmwU7Qb2mIiUTG
rm69TEr1AQW9WvaXtMPs/BRzTmeZV2E+Dl4WrJ+7KgTvQx7tqu6EAeA8KKLMqFhaCqgoOZNEEEuq
THTeppETwMKqS87ctATD1iMZM7+FWQTh9nDLp6fBpFS5fNx4RMaTy7LuzeOgf+MVrHx9BNn2EJvu
Mvb4O65mADKgAGOb34pHW85DTjzO/iHyVKy5zsgOsMw5bPu/BQS1v9Y5dJZRRs9mvlhxK+J9dw3i
CxVRYAMcSNS7tA3u/muvjEbHEYj6bv4dCKbyCkqB7az+plrOQC3eI2jioh46tDZWicoOt7gqa5/c
RFcxTLuVtvX+tNOzigSMjqLIQFYDvkzLn6Sw6y6Zws0Tatgfsd1XZ3QWq53k/YoVZ9ACxgdzffun
nrfyvB53BY6+afje3OpPv9tlpFVcBiIDIox1arkMu0zwS95q4ilaY3bfS+t0eqhsqHuGMKfrAjJW
0GRPk0bcOJYeNWk0Aihowk4ghmTRYCr7ywZXjSSDUiH4+6i1+y9ytYielH9oZi/Zo4LFZVv0pME2
+niNpQMEXkUTDZe36/Aqi79/VzzK0foNw8IsOeF78oHOqhwyZb2CgrK6SwBKNzu9zCwZ0bJt8yg6
xuBsw5sBlzlbF9C59s1VlkSvux7RTHyt3Nw+Sqd8P8E/02T9Fhhhk7Z10KUejUYBdAcYJnDmd2Fe
966QMzGD8o+1JM9Rh+wO6wdxrPZWzuAVlxuF6NgHYplT3uO/BcUtBM5NPuUXywVHupgiIgA14nqG
VUU0MPdsVrvxq7JijHt8Lfb2mDPL5MFyPPrtaPyz+OMPjkLJDRQ3LBWIC6cVYSM7IGR5K5jkzQXz
i5iH51TTyjgxRjEo3TPE7MOV1ZR38QuX/ErcN+JUek/JoDmvBR5BShelwYZIddSmZGyzOJNBcvpd
43NPIhnqOTAijDkBN6FimDyXDXxz+v7x+YuctOIM+oO+TAZgq9OVTn4MvXd/ByqknuoHCFzyvbvr
mqROkkodBFnPKDw/iDtNupgbGva883IB7OoNPey3yawMKhBFccWEjx70o0h8lBS7tFpNX+Rr31Hp
6jCtxiPfCqKTzOj4sx699BHbl2Ft2Ku/HJo0pcxesXGLeCzaqXSo0SuthF810lHsbYwLkKQDyhnK
F2OBNdnwtIN+In6vY2qYikXYtxoiwY/P3IiNZZ3eRKCSeOtF0N9Ii8SBqMSzSnL/BH9TiaPxDpIo
HKOrIfy0+I8xEgVkvi0f72et4RBR6jEkEpzyAiyi95lO9X3IUwBJXA3Ri1pPNLyDTqnyvGpfHt2n
E07/Y8S2Yvyxla2PMg4/QT63UrWdYMISgAUFAATAXp8phrrzVVXMlCeZna1cxi/wR2yLCfegW3gs
VaUWU+W8dNkuFrDMT2aAWUi2/xLpMHwpLOWq2J708HmcXU3i1pVCN2mC5c3RYivv54V5t8jlI3r3
5ytUp2DT0+6e9CgdRr4NL4kaTsmaZa1rh0+CEMJmOtOd38U2K4s0/pqp9/o0jwLx/2uZ4d/XFqEG
WrJhP9eSnmzx6NjHbLUcd7yIOCSHbUMvmXHokXh1qC33bsjyKEdUeJsP9PSntcWZBlE0zWrj4N6F
xEI0NXV/CpMdDNC3M4LWnfMHaYC0lMOmzFufnh7cr7/grWy2czCevre5GI3Xv1YPfy88skKYckE6
//52BWr2fx6klHY7zfT6aO8JxKHHhNR9bjH6SwytHmZeMe5pdp7Oj2ewtNI4H3++6E5slJT7fPdW
xEoPxJespESPBN7YAKbGO/da8LXtJbaHwNy9ARRzoViaN+3iwk05ylDJn/Ib+Nx0ME4sPsXGHvrI
YZvcAvW/PGeNHjkTR4JxHX7wYiZwG7KqjuF5eZEbbJuuXHdKgJWe8PEuqgleoiM3W1cc6G6pGvwJ
s4iJIfXubocudQS6vqTiYFLq54kTUk2Ji8ViHO9W2RibYQOhXLE7q9xbBIuqSm1M7dHJk0U+pdTq
WzX9pQUKGcfRP5evVspb7/atRZtGsn79bOkOJC3rIfs3TFf5hSjjA9etrtzxiOPsr6KsbuiPv/r1
svZpxmwCA2/5ic2CIvQ6588m2xUT7Ve5iM8/TqnoPCk/83Yii805K4QU9gLA2mzfSUtNcg0+sPgZ
jOyNoA/URhSNC8+G5SzMZyMu+OGDA7vgWQTs9MwuGse1bdZGisHMV07zqy4hbEUkEUx3Zg1V7M5x
gr7OSAXXImibnJ7t06cOtkwTogoWXnpAK6sCS9zZDtFChP4rI4pt6Te8F73E2GIMTFDdp5a4/UV9
HeKYUznlKVGBx1yDTxHLit9DHumBAM1/f+UY9O835X316FpYJ/NYhtmDQ7FqrSy8Mm7uoSEmFk1P
T8AuJspp+hnF5dCsgZ/5Fmco2eZgAMmdm7YayngzjHb2/8jiq7Z3wEOfACD1Ixj1jbtv3s8XZY8d
HQ1jWY4vLtcoGVMBZ9Gw8fBRkgNkKKCKp/JwA0XSHvolr/VF7A8vk0XX2EhasBrKwh/M3MCanmGe
8hRabKEtCjLpmcsiG9XdxFJqdYGzxHIfpZF2RmUdLZsXrBZLuXgSiXNDgHwXGaf+XnMP3JZBNjjn
+x8tuY7EZbptwqVY5k17xl847KUhJg0I1uEftYYMd0KVD1NradvSEroJRvmU5czs+cTXb/DTbZPd
pR1NVn+QJsR6ciInxnYmNVSwNxW8niIuy2eFo1VQmSoFT48tw1nOGSogxSLftq1rqY/vGC0ZV/Au
BPl+qRw4NDfGiRWeLdTQx812oeNCu3bp6YT2LI2IUUvExyul4ovTRpDZX6dDxu8e1Nx06ZH0YqSK
oPwcaiqewdLe+ELu9u9cnJUGfjVKUyB95ljs88Ddeli1i7tcDDPCXMUCcwnBdYSbMys4h5YPp4jc
iEoKBS6Ifw2VDdjMS4ApnM8h7FcRG0baEcVn8QIaTmg0GbLPWysirmnYxbomuHz8/NUv2RKV0bVp
e+O82PBbUT5j+ZFy47k8d6AN1rru9uRoSOhZkkfeguQXCq3bMeYLvQkgKpjOAH7tkPwqDwGdBFO7
FlZfHpcwF77N7RsFUm9FiFteEyrxBifiKcQAEW19XeF/RKJ5JBoY92qu/fjiR8w0b2iVfV/vk16H
fBzFqDgaK9TBpDRAhXe+Mw4Adhe5AwS8imeeTXCOmhsyaEUn3iaJkzLhYFvDCUWdYEAP+4Ggw2Mk
UasOkrvGk3N7lHrTLRsr0rKc03RE+IXFiQA2XxNj0ETUWPaMatGpoPj7kuulTjekXzh3mlF6OlDi
zIvrzu5Y//RI9AtVWB7KBO/5bclNSsNGWLsx9xlw8Q0/0BWv+gnmH0eEkEcmlLjRMAgY/buPriUO
IzOmgc2xz8sDDzpqr4ikslkxuD8YSt3+/5De5aw3/sgrObfzSKArc1mxROPmsviaxpoNhEs5WRHN
+Q288LZqj398b4/KmZDL2/IKGrhren34t5JCWRs9IkZoTkFzVZeOeMpi1FW0QPYcpEeL6KTbpN1W
fpb4UaCUQ/HZRG+AwMuURSgUyyClxoESFpMRysfXd1soZkSKuTp0Zmt22dDfcw1lOYqJe384E0Tu
JwXnuqLo9aXFDIIbCN8qlcolXt8fItUP00A6dxa7vYhDYHJQ0cGmoaLYhQclh58p9Sul3mIRAD0j
YBCfbl32JNiNljlgCkcJ+NoDth+w1LMhub5bbI3AeR2LjNbkMHoqfIUPUKNYDRnteMClna+O/uHJ
mJYaIgVAesS71kYE6S38G8yL+dfbBoNup03ATaFOI/13Ds0g8jYug6C/t8OgJsyvrUtf/jpRuBad
NTDkWRJLAKAd0wDRSUeiGE7jhWeH9Wqn55bmQKCVoVUmI0wbSbAHZQ9EOQ+9SAkSvqJaU7Nr/PcE
Bs3kUpJmnf05Krmnvy7ygab5+GefBxEwaKrr1VBAo+ye9AlbK6KPJE6jfzGhM52/KWNE0DaDuq3u
p03x7TUfEzHZLfyRfPzw7vq0hIG4WF4WczvDAHj3Bo9dF3yLrNwc6ITJ8z7FIZFCd8I5HdKw9Cwu
o/HoCnMt73PQcJdYFqA0sEKGnYaxjiBS1FdF7DvOwny/xAdRE4w9LRYQtLxJ3x11DVhTi/k5USig
z4zSROSK8lUKd2qxfXQOp7aeewEDy1saETRa+lTWOzH0jDyHDl11P7QPrDycaznktWug6uFjm+07
idGoeAoqoyniCzKEQY7y4KrUOZ1ZmLT+kpRqVt3fFRr9EbjmMQKMuME6nEfSoPJt9WCGJYlv0/bC
eifStR45dYb2TVNDIlYK2DU0a614vDswuQfgJSo5kVuRxQAa4+AvpsOhPngkvQ27EinoJzVABf5t
+N5Kq2n8AaYznknfhN5Mf7ZFRRCowPp5nRjGsvckL7gKMstCz8dbptRK0TCK01ffA/xdqfF8i7cR
V/7LzNHXyL41yywFKKbpJvuqhRfJ4YERcBUGS9HRTrKyPXoPh78TVgRkPDgoBU8C/zKZDIam52xU
YCSiaVfRxcZvlKf0TMBtJRgFdVXmfmktZJHH+sBh82qdjGbSkj/Wt+iIhA36QU5F6kc7peobmH+r
TgpGPBLbaRhSgV4mD9mZgpoHtI51R9myUBYaGA2WP3lz0Zw6gX/9Wz/hk10S4hMIOtmtSyJM9/YI
24Y0ABBKafwOSowqutQ9gfXOKwxe2EJ9a7i/raTQ8GS+dJ+zoT/xjQzs/oaOFZkj7piwHPH4hhI0
HDboz/OH8MUSyv844E36H6IZdyb4S3aDQpo9J5FM5pLTRKUXKc7wStZx8zFS5fUn/ZeeRA8NwC1A
PFC3NbAHWdbng1Hay42Bj0wnfblZxawQouexcoYwU2vBLYAq4+NqtSiFonWM/jK+7A966KlLt0Vj
slCPAW5Oa+oDNT93yYk7iD60Z/ID6bApbxsEISq1+YZiJn2DvsZ+SJ4lkK5TRlzvwjIqsxRRWD+H
Pco9FUipelVpm/1v5aeLM8k0lahVIMvxnVWmEOSTh3XwdIlC0Xd7/CZExfYmlizaOT7Z/g3caaDC
wmsPgIU8b3cDZ5C1gBwp8yhx/neeBJzKLDCY2Jspyxl3tdi87oorOMmarh1M14WScmxn8AtYcWRP
Vn9gmbEWBfdhGlE1p3Iqqo/yyOkoVolmeWWDoxPCSRRQt7lgbz0wgtN3Z1c6bRNvJXlfyRrLlDgl
uJ3BQaJIXROmb3R1FvyvJmGiwoRCfMSyY1wMKbyge8S4o6OKhwlVgVQFRDiCVjl3Z5cIKQ8Mb1MG
nwuW+AmE7hq6AQkQPdfq8fJCHuCVz0w+sQIWY8q+3ynKKaAg9CS2oCrjl3ZynOwxxr8+GxjYHx11
MgLFW9t1ZyT30d2Ka7H+E5di/t0OdBD/ALC4adXX/ss6fYT2hnnHGbVcAiQL+xEq2w1o5w1PAOyo
WKUBe7EPQ6mnrPbCheYk/u5N13dIiLy9JT4UazgH/661YRHopDMxcC9q5Zvhq66KfKDUy5vTNBUM
k90/6ei0ivZJSDTt0Sfr4cNuV3cmsgx3mgLl2IEGCcSKb2wfTfiaN5sSmbzQlToHpyMCBFAJFrnN
W8naplZlA/u7/vx7CdYp6z/9brKP5KjaxQA8j6gLO7vbA4v/G9YyFVmlz0qJN3h7psY3jhioFUr2
h1Kd6DryJu3XMeqA/D3ge5Gt8r/4zq7megJfksAKK6talLYM/C98fMhDSET+cjm12wA54U+lMS0A
ys91TOdKW7dLixhEoI61xmtazS8q9JD1TELkTZ8KEA+YEDag6B4my4HtKhzB2VrXBfIUNabcAsmY
yPz+obN0cCTAdMMMqbZJ/kDFpJXUJy8grDt4JIrc8DlzZ8Ykf0ndYOXVsXTTe2uK4L/dMjU/NMZS
R04Zb3EFJ3WdKp1SD9L9HOyezw4GPfsHgkV5RLiDTXJ+K0+zOEk6Bc163lWFsb16VrW5avqpMW6O
dXxLNKU/1ItbLZVb5fjBRSNOIiF6eKzlP87M0TrzR32/sgllKv3N1nY0zUf1htuo09ciarq2zNHj
wGd89TIhKJrXIlLXrcnUI+ATncEHutJ14d6rY9MMuRPsV8PzVk5lFOgJHaukCYSiV3Fb+KXdaCUk
JVhl7+NBtK/6VD7ZzxGLwKP8ah32wNnZFi2p5MWuDBQjlF4U2JohIGQtvVq/Hs5cy5o5+F5JFjOP
4ElGin1lhCTz0M7EYVcqht1EtCuwPQgW1HSXWkVLJA7AtkAEr99+9e0nQWWdjQRzybet6rFO7cQC
a5mkfsu8If1t88S9eJDSpuAt540mLv1bml+uxS2YL2PWqlGpUo7Pxh+E9mqgE5YEOLNFxbQSUN2P
2HE/CujJnhu7AiPZh+/bw5/puauHVZ1gFpZW+u7CcYk8c6csS6X9IuqaizSxnLjGA61cq+5OVLhS
lishWovjltQJMGydN/GHRjgkasC937SHFcHpEqfaDAxj0RERMfBn37xk5Sj+m0ne9VSaf9q9TQ8l
nY2z8YijfhK6iEfgUuIXUs1QPt2ZGXzyjYJyVrUyL3d6gepeuZwDXivJIEaM2FXQoRvv+NWBXyhG
LfAFkEGVPbTGgJE8sJDLFYHn8YWzqbhhDymRy5te19B+ph8wAecDeYXp57f/Z88aNGygtL5VaZ1l
JCRLH9c38t5heLVo7TIDA2/4onVHv2qaUZQnEvq2innMVF8O1kIDVF6I4kcPFuOrS4xWaIRLchLW
G/BNyhVxoX5vhr2WoO57wM1PWOyxE6s0VmEGqQdvxBc90wwqyvjuVXK9oYE/H3GUs9kDqayW+ABf
eL+sYmjs1gT2I8ccI6QLtnM6KD85C5xqz0M+p9qjB5hp0b7GPPfYnpQ3JTMlrWb/ipzmCqXeQfT0
kvmYwlXxxZ17cn4j+O+zbq4kobTulno5YH7DFhz0cFhiPLE1yDbEEjo7Hb8yPAImMhVmCR65tV/o
5MZp2LisDx7AiuDmz6f3oyBJX5h81rLM6RFBnQpOSryVhn4JwCrz8gBBlSugx7wBAeJVntAoCyS3
UUGQIzz9FIN5Fo0L/adAZuqX8Y1oFHfwJRTiAA7qoYfsS/I+GPnS4PJkg5M24xUaJoR/slnQwrKt
cS9wo4BOgK6DgqNf/U6TMw6t7pEsU6LXGVipP5D6E+zn6Z3iv9Rc/mVxp6THDhbkf6pQkBEJ2B8U
n6thEdDBO1vo4hU2m5PvzBvCA6MVNRXKYSOqemwG2EbEYXXOKJxVqLFSlodQSOrYeIX/kFjFTc1J
S3q03LDF0QQcEqGpcJ08ANmp9EwlGgIzfgYnVXXgTGdmS/Er3/+6fcTe/BCsUNFlsejFonVaK3U/
s/bJ18P8tj4SdMnEH5FDQdqoy6oA6MYYzftWsbzrWaUFWYXBWvanlJnLBIvVoFXs7wCGJYVlTaK6
/rM+GjBNyWpnEr33+5MHQRsfcCdYwMMwqiyk8va/4CuzQ3/uNcp0LPAiojUOqZfieQnjT8jzolUo
uFBZvY8LkHjG6BhhCkxIEcRGto3FBXTijpPfmwNs/QaYE6Z5CX1k0t8lyKGZJPNbq3NTEE3g8BuH
8m/wkRsrIaPMyYqYnOcwE8mSb2e7B81R7xvOWyW6wuWW+atfIcb/s/l39v9gtALWB8+T9Ezu2WD1
4DFB9WFpA3tF7OVTjDW/DFx5jsD3wZ1PnQKdlrFaGsPuS/fiQ8nYSlIUGUvJOfTiwR4QWwPw0Rtg
2Si6sTq0heebyn+FOe1Sxiedr2PipWDSySdIka+bS1haRcVWimzzx3W8iJEMcaBAZ2LAGAsTec14
pkRZgQ9bQ4NsotqRaMprO58e+3kTmT22adgcagE8WJkoc9iKFgTwEbriPatUcWiU/LyHE0c+6ZZB
AY/CcmQjXDT664rLHcjgEAdeWXPSfokUxlUU8Cl7raE+8e++6VGENrj630MMdmiQx/c3UkL8yePS
KxbX2YKkffRwDPQihm7g79QR3XwMo4o3Bx1sFZfVHcNwZf1Adl9ENtll4rbInCKBlUQpaF5KUySW
95gnw9/8SzdVKYB3t/630djWC0xOJRP9Me5On2cM70Wble29jsxjrvYU4ZmAgWlb2rJGqge+9/Lr
oKdbvJdGA0HsOSyM7JgUkXH5B6N1WWxAuMZuDyELEdocdl6G3U/d2n1X0NHu/wdlkPrc0+PR9Au2
7dkNX0FB5vXT81tMsz0b/qKuUQ177jNJUDgFEPFG9dZqYG5FHNR3U+mUCKh6UHZsN/1MiW1Pb1r0
vkfHBFtewsmU03E/crnmI0WATgcbgVNVlQtMU2I8jx4b246Mz31fV/6SURSjho7ftBX7hq9PRiKA
+pLBEybRsbjT9noGnqc1QVQglZdbNeuhrw3aCmnzB2KlC+02RW3Ze/tM8WsXHE4r40xCPg7v96pa
8g3uBDc8uP4Qr4OEK+GJBYaE5BTBqujCgAUsluHL8zSH5SapaJqNcuj4uqy1TckZglgqcPo5OD+0
uiZOD1qm6t3dhhCwMyLHAUrOMBpUdmPIMf7VNmJxDxn6Rk+6BGvg8xOpWffAERtIBeREBb6I/a/o
NTsMSOrXQXJgKsyamVgkN55hQoK0F97ijKsxYiSMoBIZaY1hbegoySUE8QVhURpZp11S05DbdqVk
9TGmPC9r8dd4VyM+rpsGRn/PUbuDH17zkdSzBuw/iibq6KMvWoqouWHTep4+N3d+WBSEcgyQaL+L
0Ol9csTmtnSmAbSOPTvKkPUeSHVQMAxISOB+Z9B2NK9zCFLvHTodjybdl6NRBXS/d7MHuOex1Ny3
/tmrQd13ZzEOr3Zz95XFRrxX6rDQmPZKFkJJaSARZvAYHiOftyTveblMbFQ/69IjSeZCXvbTspdl
EhWXOdqztYOrwhMprQBBJtJ9XT4XxQuOGMCNEmFZqYGE3HW87Hzo3ATqXLIzH7f+CyCfbwiRvxFB
HKdTKr3xNLaqWhtCgPSCyH/3iwlciYQvPiLe1/+t/tNj4miUQdgvxiwIlPvsyb7iWb30mkH8yDII
MJTX2rLqz0TsUhlSU6wMsT0PrZkqCOLOOw8ks8uGXcgKMfKn9YfmqEAOEY3HIlQUiP8f9Ual0DUW
fPA4WeMTy7HLtH+M/OGLnwD4Su8OsWJ8z0HKTJXhhw/OACm9UYqwfKGUY2scjblXlm6e3ngP12pB
fcrfSEjqsfNDWv/jh32oZ6rsvsBb3F+Q/ruX5t9DmZ3I3wRSOU50rD4RptKeuwHdvhAomGOChSXu
6/COC1zf/4IatCdE4RuAOkgr40Kn0dTON2Z9F8TUHWa/mPUDCb7wJ4WeBgPBIqdvF5rMz56bECFG
3lrvye/M7a8IlFfag7xtX79Gcl9X+3hrcDOw0DFi5qc3nJMoImKEBl6v0mKXpJPjZp/2KAmtyk/Q
ES02OwOOmYPx4+PW7y1d2WctMNu45NDy8ATBiBOrnSDSmrF3BadM8j7T9ClQWSAeyPAIKzGLLWbJ
n7F5eXkV+xi5wz0ifHIo6lqvfxH52coqtwBE3zkLQpVJdewZXo5wU9E43oWODveUf+5E8+LSaC4E
MEQPlGRCUy1c6Xe2Tes7WUvJQSHvCVSfYBtCNqTu31oYxSOZJVDPk5bSLCkjvrCZU52USmRHzUto
XzJtFtexjMNSRQzrndSRgyq3SYkCaEyleYeJUpkN9qmTQW0+7/FUlYE1bfPC0f1uclTexTyW48F0
F342R8wBWtZQaeOKIKBMRKbPuSNkTHFMEGRIA1Mgt8hwpxiPm+h1wvCbFUiNm0L2H5SlIGFSMIIl
x8rtQg6EJawSGXvLpabrsc0FV2XpEnF1YO0fbKtEidVUaXMkZQiEUUWk3zWLQXgyf11FQtW+fPeC
6J9IjXJRdzfvBg5j1c6O40/3HVosMobrbbiIzCNSVw8pIjOiXbRBHsNMGEbxjb5iVhGq5HREtyKK
6p8KYNNM3YZiwv73VCNRa/zZLqQgA39PdGDOHNvBwKg0XGP4LMM8S/byu3j6nWKkrkhOBlV8kDdv
jlOtFXAxYPVbK2Ofob4urN5TFe55U9mOtpMVOBnJgk1M3NITmYTycnImPzjurYEhtntPNNMj0+67
V7PsVoS7FeWYVPh9h7QMbiggUH/TDmSJwgMwujMBw7TBB+CzlxsSqFug/SvHlQQnk5VpSAShtCLX
mcbq6WD0NIObvLw5fhGReDO7QUyyQa678CjCAasb2vxJS6fcMhTkW6IKQWxad1z6zxFCkoZCU+vi
t1j5QojaiogCOSV0IA736398y4HlLWQX2gYFo4nByguWG9H0ATP4QsjKDhmN+fSoyp16dSsEE1vS
83SDKGIQuKZeTXwctXPEfygwNE85giQHvScvAM7RPq+5Y4uU6ABUwkbRPs7b2on68+D33SrbEPSG
3oaGcMHm/vp6gZl+jht0I5LDmralKV9TtnMWZ82BtAVnQDFa7tLjABNU5o/Hks1vukwycQCRJMzv
Q2gaf44r3EBXj5lHrsucY/Trifkd1H5/+aykFnX8IbAQWgBdSeNBWOjufJOVdFNGTvfnqbDlwo0L
cJzUolMo77jcYrkytkl/k6qi8VvY6poUdEghKEx9xk6+C0RO1Sea1lDzSVsZPq95D4NaHrP0Z1CL
HgHHZ9W4EHVS2w2o+HVGyxe6GEv5JPNCeikGKClhbJ7QMZNmtSYUNlnwNaR2KsNBIEJVtmYC0tms
yO9ihlkP1DaVdusHACpridmeRhQYRSQdR/Op6cHgXmd5SYr1Z/k0hyKQLQkCHCHggjrQyi4g9WUy
ibmwr8eHf5lkH3YEAHDCJYKFLivnwewAzc3LjfjCa9zdmpMksfZuaC3YI5+fWWGGWBT0mJOKM5Db
DYWCt31FKRG859M5vAZyccknluXM84qGTj77DMozfiMCzpHyHukNoTfIgCl8PPK7NK5V8B7dL2LT
ncvSmuEohST124Vl/ae2Dop/1lsX1+3uLkz3AiLT9QTWUP9haEFwxuojJ9i/BwH0tLDEsvtZciux
G5ravEFp+KHsR41tvVz03y8EaNHJbyC82OZgcG8ptL9st/Lw718D6fdDlyMCDDLTlJDjcMut5Moi
OpXfsZom46GoUz24hxgBRPtZWAOG6ruvQ2J33upP9aboZkyyRJJ0Vbe17gJ0s/52XRcqloKfHZ0W
px6MqbBvM1hUmibmEJE8oUJPeVExULj+LPyL11TEONw64vnvOITmlO9TzwNIAwUudIVAJDLliFMN
Heh54QE+hwl09TIq4a62JTucVEI7QwMz0q2ArLgsIgWwrAxkTVIoPAlQ90kLdHntGGRiCJeeE+0W
z+r0X51Q7XAvCdd32GG+75Z2EzQrumE9xiT/r3Gcu/OEi/gDi+SG+ZrIHvIVpRLUKH7f1vcMpt3w
tG5x82AM111uePIA381bZj++G/hY2rFad7bM8hblS46HQ6E54qIdabopLZJXPsZ+esca/KKn3pQ8
L6pTC6OIQSG9K5PEYaQBjUTnQueFRBXBWpCT23fPc3cTK2pO9oVlwNBZzljpSJ9wLjy0yciYETV/
cl2TbgL53VoV90WDtkMx9+APIb30WawuA7hcr6zILEbRoL61OAnsF90uNcXeYtLqEwN1Ju+2X9Xv
wSSQWpZySFn23N8oaVTStrLVaw47R4gNtQZ5M+gtm+kxI7j/aLpWmltpivzzK73H5KoS+wuRy3rX
E+JYqMrI3VhBaYrcBgN6GVKt+tWVd4lQwUWQIUG1lqptddUMWW9MzK8Eft+9Jf1CGuU6GYvf3g6a
B4yO+Letnn5wboFkA5cbPTswGZ3SxdYPNPZhnVUZ0fdAvbZnlYkI5zJPcyQx54JDszd1oiuMP3a0
XgCU+lxuRj3+gjFS50X0JcENAu09J5s5iPprI5Z7a01a0fjrWgfgcmYZR3uQT3eXjgKyhzMtEFmb
6Tyq3vrjIBgk9KDPclsoNmr6qlXcZVcekyI36agNmH1bPXEZ8LnrgjULsbKDWPQQvcMhZ3X1HVfU
jKMC9S9PGJfWGis3arAONOimgvwsvoHxkCsbh+qa5YxL6eicgnuEa98PKURZnvX8G921U5q935h0
36ONDxegm0Vt55uYajVCDzMKPaeFO+26+iabVEuln6Tz/uwMS16PXisj6tVgmZ3bovixhI5khpQw
fB55p/c27+t/eFXKyW2LdjEfPBvn0c85Ianu5RItpVNqcohGFXNFCcugmPQ6fS8y8N/R8llLOSne
ck3wPG9ZmXI+2oMg1WKlnG3IgwY3ZnQHpQSSeLLPaRcNO7NzG9YNVX9HN/4cpCCtQXh36sRqWt8Y
FIx1fAzVYE6ZhxfgSB8mnW4t/SBXrssccX6yMNwEoMfKmmFbmbN0Ffqlj0/46gdJkhOEGrxWJH7T
KuJepn52zHIZdJC20SAKFSiNQnuty4p76d8HS95//IHK18LhQ/E7zAbJ4ZMRTy8gsOb/YzJwKNzy
QlPd0It70ZjCQyfjUjFNRlOQPHxfhCaCc4wdhzLr99TurEXELsk4Tamv+448ZXLLRlD1CbMHSH8Y
thcgRVT4pnSbOFHI4/4XZ0RFp5yEroc8BldMHIp1x05aY2jAFy5Tn8UrEdC/8pI5A3jGiwD4B8GW
YyuppjRMXJ8v5jwvCEemHWdTmM/FUdhdiW4IFztqnk6iWzyEb3UsqhqzHobjz9nVv/Tgkx83sbpE
qlrugUiUOXwvC9xcQ5Q7EjdfhTkc+zxnX+AKFSOIDzdt7b7utmSAeSS12BHmNkWyAS5L0KC1soLM
RTz4sDQULAeRdc1nMnXIIbOTMRuvLv3BLVZvgfAE4vrdSK/fZkU7OnQNFsjxaHnGCPT9QoUxfbbn
kwk//AmlWjkIv6vgrfVW0qERnReUqekD9NRpUJs/4QJBkMmdHXyNOXmczAGM44MBpMkShO0tmojk
yOKt8ukbEDDQw/db2Qi7+scIMzcDTeR13taO6JOJLXTZ+Cj4c/EzRO+tonEhN2g7yyTjC+0Pzeuk
tyt2ZjHBrpFOL2SJ/hRFH3xy56Fuf7F+Yrn6uJKqDoynbkzOHKn4RrENlHs5ABwvrn+FFcB+qxta
E7RBOYgU8dJsup5UKuRW9r2tg9M5wb8vdOAsGjEXg1b25WxC5OOQs24o0OI7mdhqjzqN8xubxgQb
O1Y/zISx+3oF5OAhu0dmIAt0TCiLLPlSVkOb4n+/g1hUIT1RuaXbVGSDVrpLOdOprQaCha6gIbHD
QxqB8ychm9x26HdvHOOcU6nnVr+ByYprLxuy0inzxlkmnxk4UxxM9NDOjo55r/qdTlwJ6iIrj7pL
KD/NqSWFzKs2vaZZBS/04YvK7txbiuDZ/+VdNSEQbce1Fs8El9DgdvpxV1P687hk8HWWLu09w2Tj
AEMpPtqGqKi9Dtdat1f0Ph6nMOtXH1OMivKZYJUPfo1zP1hjias0I/zGppGul3Ki3tg+S6yklKxz
K+rwPcoTEJugbc6G+VzHHk2kRP2mhTE5hYc9BkMCibpzyRcio6oqkab29NNvO7oCRsWMBpFXIbnQ
eWpPjogoGneiueYkXWgQHu2vKUFcFgwZNglVnz2pb5VejaDJedyISxpxbI1LJldnPC6K/k/aaub+
70SB5C3D/CS7+9M6ftlEwyiFu7WVGJ6X+uK/yH5byGBM4NSabVfNwAG62edCAl8Nbfo4TC7IKRDl
R+ZS+cgTu0hepgExYsLOwmxXs9hzVa1iok9zRYtQeo3Sl2cO4XfFAbtrf/QvJrK8cfzsIZNVsUic
id1czM7fekKZdKpmXpM8Z7rpNKdzX95F5dBFJ/QOzZ9tT3UASs9MphBfPv2S+jc/Mn0e4r1210Ai
9YntEqgBxbhL2JFmUqdPdt2baOq5cn8Tk8/3br6criGMQRnux6F16iO4su14yV3HsDqXmt3ZlsX5
jDlDJncOU0J0W8MYpDeE7UsfXnPtont1keCgE6pkdtaqYwSDQVglT2EZfptneyghLelHCkBHydqm
b/i3War3zvEu7Nyk45VBFCeSM4m1B/SiwnYqq6Jk/8AQtBY5MMg+eaEGTNEuhsjXovZHQAyelfLW
mubeK0Mb7SjRKajFGSB7E8n/FkkBVGIwGfmLnG+Xz/YRo5Ibbb9jIoaAzOdFudO7dqzq538UCM1o
kJCTYjBYelIFhEbMfP6yZXrrpBkm1dolMU1C7GGTXcdWK8Z05ozIR0rO/UxRczW7OySvP1STYOgO
qHW7tFQHbxb9f/gHYLiLv9p/H3Dysdd4WYcPAWCb7zXsPpirF2XFZUK+qLloFTxY5+nHX6bcAfqq
2qr0YyZ3gttDslLIuMWs4ucEwimUTO3qhzi+NxAoqMk76St2FK1Wx1TNy1oRL/JHS0pqC4ey2gIZ
55g38m7IyHzsV8xz6Aj+Bzkp8LnKr2NL6Youzb4afxhziTV2146a6fRc/1ZPUwgR8jMgEjHXc4Ko
YUjpkiotvZRJqaYMdHk9GuseAzDYJtq1NcodEBIMWKXQV2I/jRL1Vn8Nxq3u3uJWcnuNLG6NMWWA
PteWByHy7E2UQxjBvXFucFGz1Rwr38PzV17L1BjZzWYEpy/9L7rRMgFlpekOY9tjxFKs7s42vmH0
tPQgHUp2t+8yTeq+9YPDeRcUVwIy/M2NdtzmewOiJFECrkieWsm7MHh+pUfOJjS4UW3T6rVGQN1a
spJ0jPTwgH8dQmcU45Jy1NyqT6fDAfxg4G0Qe4V+utjF+Nf0q2z4VnurNd6WbqCx0HV1P3ksl58S
bPU96tgSZa0YTuCFs2Zfv+vZqIKz3GlYHOAsHbY/cbXqM6sp8eFgE/WuLu4dBQfwcdLsm1dYTFXS
XqVWvw7VTHqwx8D9ydlFDYjP1/E14v8AnuxZ0Sx95MkFpnRMZDKnnGLwmfRrG0dLRDRRVhD1o0Zq
Jc+ZfOsAELRdOn8GvpBM2eCqI+zML9PCDx9p9mT/KXmrCBnEYv5HfjMauVPPHMuHCOfed59D0mms
JN634ZvMkGwJ3wUTyJDl9VmROnr5ZZBLXgp0ZvnoXxtsuw/QFg+QkH/jF1+s+8k4PPOYAkOftuCB
rhD+7Kx4YtApL65avF2Rl9t5GP2XE2vFTs2HgJVUnmPf1KcI4E9UDMcZmijlyRSm8W7swn5U9Vk+
IP1jv47n5guygI8Nj+pQqq+ZmEwanXcqNnAMy1JjuEAEzUQ6VxhRGnNkGbR0QJFodRWjpk2NnPSC
4cAOzAPMlzb8qOmtPduMJGUF6W1omPaFBvXsswcfApqnuRE7fJ77JGfnCGajAyX2CFXBuvtwYVti
VrtYwYWr4IdLUfiU9GUjnru42h6BCWoeZv+o4vSkwKU4zwcoVdqxpCx0g7+q31pOmQtyrlysUcrn
pCPuLtgOeeHFGO+q6PsmYbojQ+5GyahPwMo4G2UU6r30y0Paa6/MtWsPw2CFQVxattbKOYDz6qL0
Qbzlk+BvdtFW2eg461RaM6rMCsG47JGs+tVJ/0iTYCokbWaSyR+Ix84EE5v73dg4xxma+3p/K3fS
pfKqWC2hVV9NXo1RD/sYy6fAFD3R4wTfCIlSG2Mo4eXtGU/ItYlFem/HFCAeTlfg3DiFLPN3wHKT
pWmQ9xi+Z33F9LxDJpgGgK6IU21q6FJUAcsDF0sYQVFn/bqMkD5ODe5WiWLERhHoT0P0p4wPmvC+
wZysk3yJLvpFHXvq27UVLg5pGBvC4qalioZq1RJqI1l2DaRP0R0LT6d7SuA24lrQEB9GllB7Z2tp
zSV+xG+BMIB/ETPPILR6/c08Ol4JoaYveB6uRxWxj8HXpaMYadzbaq1ymxqDxOIMRa2YR/DiFQ/a
ErgWhqzDCTSOcF0DszzG3MBkweuRhXLkez8yt3uNnpHFWBtLOntv/xZejCEpV17m+EW7elUOSbGU
Q+RXj90z2MDRYBkWhb6pCQKWZ7AqyGlVD9wH1EWK1CeqtbyH0wcLvCs41//Qvn/IZVG2YSJC+YYd
NnnvtjpEwFYcqdgqo5VBJAfq0zPIfVK92sU0vjZVMRNVmBSOuYrI5uhTobRo/mLDh9qeR3QTm6db
BMaymGc08yHEuExR2bppCiJTdZQMRU0u5ttsAlRXNDymPRCdMp0PP80wEuzjvtnCmTW/kNyRqS5Y
W0+uMT1pcMI5knOSW4jm6UXN6DfOYy7vcKSvtf1KqQUpbxH7F/a0eRWFxCoS/3HZ5HhKdYeT2w65
XcC6crBA4rfrYn/Q6wDsihpK3zvM/YMPqyI6PTkH7Wvg4uwpYXEk4O7MsISv4lNCzwDp9mKkrUvT
+DJ4A0sNWSXkOvzWNOyA6wKCEUSpQCBqU1RAOlsJCkckjgL7ERYbw/jiDpSWv4Rvf91wfMYeJv2H
kp3gx+jSShJ6QvnZtcHauVu4Y8n3TIjGxDPSEjXNtQrcbGOWHPqNwjqYPRCfQQuHpz8KEeaalI5y
UB9NaomEwNyq0GF1m63q3GQKIf3Q6Rl+YYZOYoER+lN/ncNsFmTCUq2k92VAdOykt7ciWLPk2Fv6
2jLZuXC6ZPyVRrkTEhuMcuObI3CFAHW6HYADY3x6DiAzttBZFLQROFtidNsM5Gc3qWodYaL3Yeh3
rSKZHC/R0DSP1Wf4udqyaJ7mqvDcTTHpLFoTNgh97XE+mRNYbk3hPl6pHYHJ3WdC+MyauCHuhJIq
R3kOmmyn6VcCWnIWk6r7aR3ypMlfjYbiViooeFxxDG8rSQk+Hg9KuZxTgxtDuZcWH9pa6CbxB5GR
JCJqp9R29Zi1hSrIGjstMo2oXaAHgTeNaZKzvR4DPBpLOn1wdb9bDHILKi7WtJI9RzmRMygabrQu
Urn2ziUH4laY3yqSCfww/qfTnQvw5G59gwT/vq/RMpRPG4Fv2B7FOk3ysRZgU5LmcX2NnaDRDYrl
iInocqdlz8oUEJADRZMLFIhE6nong48u1kFEYd3aUEkDvffa8nojk3/GfvawOizWOp3+MMbEf5ky
BwLP8gfLZ6l5w2a0YMaKawBrhc8zc+o7vv7arqKzVgLRLy4G+gYW6xwEEoo5upmxJ53P+cLRkcc7
MOw6iLuvjIX7760ESthjtgMxyTWYFCt3wvRMQpZR7Qvj+q8+myS6diZF9eG/NPi5bFnw0H0iI9aw
wGNtRCJa0Mqd3f+jB4hlfLLiPHwcFkARNc1p6sByEvN3ER73R9wGafJaACVfpbKiFxNmO1JSPAFg
sCcKHcDyPyRg0XEvXvE+QwYuLgsWhWRl/Opt3G4MUj38Tz6fJjRRvOWebeinzN0TMAWRNtGzC3NO
5YvDcjWKLaRzcKsoNp1hB+CrwlybyrNbFGaSASQIJIrT21R/3x2U4ieMoSsUW3XxIBgDuivAVNiq
IktTPEaz3hsdj6Ve9EYSPT/pJ28+NLE0NRo0/VtFUOV2HIIKUOlEyCg3MZQmurOviyPXO6+XEYKG
k5HEDR3zGxvcWZewmUEh8M/ikuwaFYUZQQ60rDvwj57P9znJcnAP9mYv5nl07mnqfZBothTvCRHa
FIyr+u3Rm8KeOGsvEBYiL+E4xnAYhZSVhwlV0PtOrtHE6r2X2CKTiClIHUUEFeRs9Kb31dgt1X+r
bS6SnPwIQNDI8YOL+6r6OjdfcWdL8pl+OCR04+qriFBBsDs6JGQzd3Cv0QxtLi9TFBJEy2WrE/4n
PaLp2wkzW4CkgsjlbaSpciHzDZZeFoMcvCAto15vUjGFnz/hUXzt8xqTosLcM/WrhqOEntQP53ZQ
fqP8LI8/ljXH6mGdjH0428AKMNEmgFtPI5ssQPE3EgoAFkmxgKQQYishVWpMK7h2nOvPufZTyDJ0
Yyi5eLFbFT14wdMsGoWOO/Thyl5cPowxj2jDw+Q3mcDMHDb7QRk2JHEvDjKggCGcplWPFiEHhpfs
gdKRM+H1zSZMGWnbJHuYFyX9R2/woga2R0/hoYlrZOLZ9jwMmfTRuTGMk9AWgmQyVUBSX2ayttOg
zB1OKN21Oqmpiiqq0IwbzFj2AqEZBQ+lJutT9jWZEVr2s492qowD1kGnptHjHj1n6MbsnT60Xp1j
UlXwTFSgVFLV63W391KMrWzQKwE9eUhYBNUmXzBi4t3JPI+TSiR9VFyJf2gqQQgta1jfcWf40tBZ
Mv6ga7D3RPukj4Tjt4xd7doOmooy3jiW9UsTBpv9n9LGXzMXIGSAqzwftuY9vjmje3OkJc++eLYL
Fq4nrpEtW+e3G3PH4x2jHJyCX7v5IB/Z1lkOLgTz0OaHPTEjB7DmtzgAfJLBocX5BnLa0cNbwO3t
pj+ORwIQihgZKGs94piCr1VwdnStyqDq17Ky5Cqc12GRR7Ncuo3iSQPBT8OQnfv43UTJWU7K/0EA
dBBfJv2Fw76UAfyfBY5H+2ZOoHtSEgAr2tqQbGo5GKdtHnCJoVE6leyiC1aaZeEERiMWWWph9zPK
n5zHAjksH1VGPmfN9VRWspRS9/z1YpUTGxHo4cs3nAl8XOsLKqb0cpsKFWqicAcTElQUpRyo5wOR
/vnCmh8KXxt9zSsA7/bkiFtfxEFH5NNd+Duo7CELlRocXknE6aNBpkLTMH28slCTkTOkj0DALOBj
aRTBxCikTEOqdumcsdYBPPqx/Wr5GEQ7E6AlU7I3go4Gqx7IWwhHuvgVnATtBYf6kFUj4FsitCeW
OE01pGpPv2Rp1L/oB3zD4X2spGoZACx1jn2GqhKJ4CkdhLsr1tOSe14VNBZkKalFSRNvAFoMYab3
Hq7ugHLMcjgUjztR6rTTl9JVAmRcOb+kYeb51DKj20TMoH2j9uPZqU3oespUDuKh5a4UpQFedrbs
TJdimXsZDrC6JByA38kxXs6lzuuvN1VyyDNS7sK857ZJdfevuYFIkqwiPtAGjllqSJCecw+b0pHB
PPHZ2T4KcrCLc4EmovbgoxM7DWy7KR7I+wlR8OinLorQQjLtJ8cffC9BCH/AydMlx0ROb4OF/M+C
Z7aKpudmJFXj+j4h1+5TGl7dXt+F02b3rPA1yvzO4/vFDvoZKcaEWsrZD3sheSHtEEXeC9rVOeQL
Tu/JFNbaMGrlscVofJ/vAufB7H27iWcBqmdNjaBjq9NqeKg8tFPB3epTk7PPlJP1j/Wgre7jtDSk
IfUDWJXHfFz2K4LTciP6hQ4mg85QRY/Rx91yl/sCkbrncgzJw/p+GCiz+TtZMSgCpQ1Emi0Ulfi8
3oX4gxpNJA7OnI9+vIkVNiVyex2GMvy8/KeBZFeHeFyeFEV9QVJ4Kw0fd1/SZ6j2OwBg/SIpOz2q
zrqgF3s8be+FhuoaW7SFiQFJ9VOblW4gWwNVireLWcoEnTZSWjThvhgl28xg6rdfrVU3PAqRlQUN
behlWJaeBlFHyId73yOu8ZAnHQhNeyUkS4ImjSK1m626J15zgmYgSYPHYjQvAGH6aUfnHaSKvBGd
rsjCYqNiT/B1/HKZd36M+bflYsZc6q6KMv3OGpHLClLCB5I5mtpk++gXe/L/zLnDhv+TiRDjZ64k
+s/lVCeeXJNbeBf6h2859MJu/zUwe9lWxjitvDwNkwZAHnK2nFV47LJbJtoZ7gENZdlrJHDAS0Om
+Ao6Lh1gXkLneCbqBx93cxbvoK2x1JFKDV9BM5Ay1UmfdJMu3TD9W9SV7kazXEv76MMhj7pILZVo
JwUl5ZIV3CQYbZwzruYLg1jle8aPuuB96VXJgnFMIh85soqgkFxRZEdsqsdzDs1GtWsmfi6qkGVl
6eyq8CYUUPHG3d0woKF0H2FNRI9Ay+xJY/u6ceI6uTZn8v/Vd1qm8T15+bQscr75pfYWpjrttvXj
DV5hXtN4BqZj41AGAPM9GhaepJ4mBEeA4BHLdp8UWMUikAelNg07pTyUinIshsowT6z1XZuiKjkn
WxROq10DpGnLPwq7VHJJt+Ki/R5HHL3TnPy0s2kB951tfoBunK09dI4+sWhy39fVLXALIFxM10Gk
zLive3Cz7XbfUqtyl1+xwyHscV10h0ouNHu9XS/6PJh5U4AoWe/zmiY6L92rNpwNsONY63nA211w
nmWHapGt8Jbi7hOZz3WvPk1GDZwWIBq2RIJvK1p6YR5pcGBAvs0026VB5apK/5mSV8HqLNLD/TBM
tROiiiiGYSGJqoLz0ol1Rtik/CdHM/L2lsPipbYbHPZpAFps2eb2iLfoLQv0pTUtuYAg81rJ+Wtu
K8Mg3GjenyzpFF7GNh7FctBLVr1qFFrk9NbgIs/bVu8U8pULA6kPSljepQdRgYRRT4vMqG5Uupcr
0s6p+TX/jlI7eb7nAFfCzMVvHaeirIVut8zdP4AwHj537XBbLu8NTM0hMuE3kIAdZ0i2gLjAd4Aj
yHJ1oD1gVJ057jUBoetH85CCaGSIDDNUkXrJsa9DEkwNpRQm0u4hCJmUg+URJ3ZQhOuZh5gZNZsE
AWqeFmIxmfkbGv3YAEBcP4uhHmORRx2sOgQ91thPw5S56Bv1T9Y+WeB1BF0ZmUyb20RUQ7gdxlJ1
bB0l+npDU/wTMIQVUVPfmvwyOp43KuoB1lOE683jXeHs5QJhh/snvJb1VleXAZrxRUXFQNknpSQu
lwRPYd5R6Bn3bPvMiwA8rgF5DATfUIBXMVisHM+vwBZIaBHYVF/XHnqhvryw/MdE6Auk2VjGCGv/
eL9sUzOZ9rMcPdKriKQzy5pFLO1GNzI/NqYZMMd8uZZJgPA3KcU+bufh+8H0EM47hNlbZnws9E/w
mZf51TqKr1QoTYNlHWOH/EgwyEyV42MXSiZy3FkkjxFIUUn1OH2U+3cAobDD8dBiFG/QTqEVQDPH
kANXBhZrYYj9tIjcLi5RvoX3wd0sXwDLxNkOw/y6htTDfGZawWD3JEtZnH5hYswMOmhHlqpY4+sU
J/c6bZDIu97fXfYDdiD3LnEOQzaS/DrR16s4UkaE5pNGcV+AZ6hyc+48tVCp7lOJ95fHpWRGt93g
+XA6fgX9xDuDfBCTBK8JSX8n9DW39MwtfJrMU61ekpUjwrb+LirLAhcbrKha4MVk3DL+zx42KcJA
/I6u9RNeZC+YWWYB+54q71mw8iLjzRbZ+siqS1i9q5cumxESAAIWrj+8/SNt2xkozVHXm/OUR9y2
7R8Q4tIVwAviXMBvyGfdiNcdEww4P7xTxe41Bsm7B99u+3Wxf6qEtTR0tEMcPAh0zD/GsaoeBOur
teELvFi4wUDWHDATFhF8Q1l51Ld+lsqhQkOQPupUMfkS+C43YskT9JWmgeld2UWpT/70ti6JwHH4
wijxC+vVYZGkeQZ8BkA5BZ4TRnQ59HZUvlsLUUSxmsN34E/5FD3RQqziHT67lzBt4JCwZMqT0z+z
U86PrwMBqxS2oDrD7EBvJpxpeKKJEgGjkOyiWVKeppEESrepA7jamd3Y984ifdtfLLsZIcWiiFo/
kCQGdS8dZCnUFodQF6Yy+pAt7feqgxtAdwb19RaPsVaTm/X3QChiWQeiVx7fLYEfwC57F5Jd14ZT
MT2RtFNCdML/YCDiAXtGY0ZRtPzQlycYASWAU9ErS1TtGY0O0ABoArleinGB08qqZPwprziGxQwO
y/ZJFVZTJsFfMYI+2YaqoUV1D5M+nwhsqeuAuK7xllinJr14yK5fUXEkuFoC0Q3/MKqYV/NfZBdg
/ZbzfZXngrBh1sOxBJtRpZxdUDHCTlpEMwhlcZ3yA4A0LcvTuCVZlLyDF5ZnC8/bdcnTkAQV4i3y
KGIIHRbxIDrHRjV/0RoM0O8mBDt4gsVGkGRe4aw8gRuqQSIBKUkM2wMGlOka4IZOiMQ0arfxaZHn
WgIojshDh+faiQk0ra0jJerTif1EyrFc87Wz+8UnVw0bnJAd+mhC70vv6sCY5z9dzGzn6+5gSjSf
evdPr5iP+YsgZJihoabl8qX288ZCvouvinaQAMwjrTibL/mmj2X+JK+oylb2/0zVxdBobgbd6CkR
SsSDdjyuzMAoN77byQsN4/7wsedvovzJA0vMi4jitbDjl8hDvq4t0l8RTghORhButG4cMmCyxDCL
laQqBj0dN+bG6cJg4ahpRNb6NWMSfTnki65VOjQCbG4tX0mJqJfKFypjvHyFxgQ+EdRzqGhDMYsU
zVt8dOuHeX+FUrIPOSl3oAA7ZTM4K8NljeAWXsUwbHe6mAlZzmO8p6D/j9SzL/kSSe2XmcUPXeBj
2724n9Gka0BGLnQ7nFelQO+eQ+1rbBp6/6zHzSKxIAlxjLNv+GFcchghMiEwNoI4KmAdm356KzxO
qeSv8oUIdoPGMlLE0zPIsZyKzWKVhU/lJeVI1tcdkyq2aIGbSMJdg+5oS9SHgZGqZiiOM6GsQ9UI
VSMf8sbfXwcJ18PNxD+LW1PADIr3TBSFR+wBP9ojVVCZg+90Ndqgr6IvW7y/mi3Pi1tk/+G5b5V4
mr4bDg7XGYSMEAe00dzCWiz7tSQCXEJddfkEVwcLZ9aO6bvGXrKIb3Rp3AdVxhISFENQrufYm2t+
N20AHv9Dp2NP5N+plbXDWkduyxIxG6yPX1w418QRKmCuw/GQ5Bs5FLpIQnBmuwwrgsTM/e5vckP6
74gPJkuhJHxBhSg7zT8BggLmxL2N6yD7J1bDzc/wc7jVtmph+hNomd3Ph/tk3P14mFvf+KeNXMO8
vREs8sXWPD9CC8UtDEJhxbwb4lt9BM74GgN8Wo64i8mnvtZ/zsKkQRJqoKtyLLViBIckpuy0fw4n
hl0X4iaT+F9ntoRwkQtHmqjyGZPbK4G3ig2St8B2p4rtzPSGs33C9d67cQBOEiyLadYun5R4UFgY
VopBcITN9RFpT+wMWFTz9IrG0chUFx3f96OSroZyBXzsDZKHK4e/eUqEQ6cxdNUi8qgPOaV4iNlf
pcPvWzM9XPC5Ir7sVPIZH5DiVgtEoWPCXF8l22urJupxpO2yVas/2/s1bKSIHgAPlx/wR4SMXCHS
H+SFd24E86GmBcPiCR8ixvZSA+RQqO20I5e3cGyRpd/OOO7KcGS1/RpnL0uwiHR6h7mx4R0BRvUY
MQzxVqnk0AX9OcprXZLZV9avgU2Ga00upnoA42MEOT+dJi1MXcBymiKXbMOhRvyRTwby7j8H0WK5
Hx2G2Zw32HMWI1cVFbX7G1hZJmv9K77yE72UIuw0K6fOa3mAr/fU1zkbaIt+94qspuB3IF6FCh+k
3SFjEcSLP2VV8iSgA0Z0aE8CIwi/MTtD8q7AYMgz5FEoDS/1LegUz3bsbGnyQE9iKCqwAjZLWAdZ
Rr8TsjyExhoGBSc6Ikszt8UvR7bT53LSqkXE9uA/G2UcKPZ/Nb2v8XYvrhRzAJakkKY/P/5x/YUm
RyXBZMaR2fM/fVIAQGBDIodAvokucl7FjAwSiMPLMHW6hxS/tVaMFRAxIKgX8r3B3edMJi/5lcs2
Srm24pnD0DR56daapyu266AzrORfibVPzrRp18upRWPb8mQx6PLm7W8+5GLtyoNu4trbpKB5GyW+
Lwc5gRWqXC/ZkP+3dlUtDlrc/U1bkdl8N+jvOwUhxxtcoYpEL+BvRmQAaAzljI9hlV1gVw3SLjRV
fSb7hFhUMBvbl4Zht+4Hq7ESMTSlWeHzUjMR/DL7I/mMuMhbepGZq1YYBZUx4mIZBJQI/jMAkTpI
z8JZNd2UPJ76HjZqeFk5JtVQA1RjIkj964dvpqNbt8hG+/iEZn1hUL+9nG/XtbNyHDfE2tzDmVZG
1f5aCC5vbZ5StulwkPF5RoElTgvdQxqVr9vI0x8X5ay4KSLw4sxPSCdUhKdFuWl2q9FHa631Uoh2
tiLJ+K1Dg9oZYPwD72sdQg4V5Ox1eBMYZPGV6FrldX7eBRVKFvnGWaCqU7xCeKUtPe/evN8lCWd+
L/K3gAh+ko3BYkbrZAs9gIAW5vXYl0WjW35wxrHyULwgwVKqPQuT+D5/wTadG+U3FQmGlUryqCkL
CW2EXHwhezwayba668vX6ZQ/zc9SHcx4qUhy/QIsxsrk7Xvy+g9j9tHc1SghdaCXRMEzx/muf0Cs
pSGSYu1EHCQVD1n948fFx9LMienPF755QVEkRV9TZoLhWRb9NJHhWumw49qaBD7d1hw3eudvWAHf
w3/Mn0IgKZnDy6AuM17JHXXfozpi4+xTl8722ot3ksHuk3fbcP25crzxyqho2XCOnclaOQ7XuEsj
E2dJ5ZH68Sl7ZOEk/AR8PN174Xo6EdrCniLeHEilwxTNfqZRYqIb2yld3plhLB+xSJ1K5hOV7DDw
DDMfb2/U4uaIeocOlJ1I0BILKxa7y/0loHiOjFZXBfLBLUIS3PCU2dvyAQ4BuTf8MvelkkGAy6xL
H0kknVPSvFj1eLM7qthN0oXtlO1VXMkEq6oXolHKuZs7c3ajhfkRPMkSrww2t5Fc0iwPcB94/Qvt
2ijVumNESRzxjPaHu/zEpHeWuLKu4Cib22S9rvp3qLe5L620lMXKgLXVeWUFf9Td0LXannQerVuh
oION3ad1v79mti5d3DU/0Koi4KrEdpeFc30upV8+lIJRft8Csmei+totPqdsDR1wYZfCVyynSAXC
bbDayP4YYhzKcnzVgJki2rKGpik2K2lMMsrj8QCvtMYA4dH3w3o3+2GLbYW3xxQ1oIP/3GM3BJ/s
1xkKUrETv6bQ2d/0pMdA+LqwupNhDvRsSOuUKiLrJHTXrjcD3uKxckv9ZK9C/nHcF6wUXCd4uPRH
ICnO9VxvXmZvWm+lhSctTZzkxHvvoRMRpoLibCSjInTmqx6GVNcIJMo1B3ZEsYk8j7C6kCVmv390
RF8YWU511sSS8ioNW8rK8fMP4YKA5SWEOUeBupAluzgyCHhg9zrxUkxJeFPY+l1B6ID217uo/LiH
+kQW7a2iSccHFs+GTzR8XYh6tI9FGeHUQ75SadUym9ybahac/swL7soefW0h8yNz4d9GU5gaSLt4
OjHklhBKYYoNd24Q5Ki4MH0/uVfQ5m4gwFEPYnw5bV0kzIots7/yINIW1MlGppUIOL3cCTMk8ma8
O6v8/h37KbBt2Bkb1wsEWqP0+K7mAWmM7x6fTsBOsL/oJDfRoPWUhCgZd4I4Cb/IHkOVzEnGrFaz
NmlvPSwADxBZPNE8JQWi9avZDCZX7rH1V0YazrI79159NR3oIRsO1yuuKjoH/TY3ikbhS8Dy1aUT
uPNYLuS0XQ4mRU9us4pGYzZijoNLTpmgro2waweTos8x+Ztu/1P4zr2HD8z/rN2KJ+nKZOsGGQwd
LAYO19iO0VoMgc/JdkF4irLg6KnckQplmCA1XpOdlGidTYMtTXEFqjGDg93k9zKrIT8bMQmKJyXf
vjKkfqOs0bI+OdhJb8M5SjwDitixLgkcgH6jctucUgVM+8t6a0KKyzpT2rq2FmgL7nn8lh4sBEmh
VA2rKDDy9vvuJI8ya7vCDxpYAT+rfJiR6yuwC2sic4eFiOR5Ms93bo6bEKF0KINteG3vVew/sY3H
7ZYM1htQjCNXNCA5K8TOH3nuPcJae+iTPsu5M9Joh3GRlWSmOqYgC15nMzS0AS7lvakJpxk07fNH
Ft4ti1L5G3eeTEs64H9zUeWPwvrhguaAklfkAnwPn3ZWM5LCynz85RagdyvgsZrvdN5aLS3s9p6O
p6Jmr7N4C+4ovOONJzn3B7l9i/DvzwQsnkoKEpVj/e4eLEjvx6irjuQFX5j4EAR8FA+/QS6Nzvzq
HzY9tCzqeqCJbWHop9lBYxrYvE2wJcRQhrFGRWtHJtWiQWf/hK7U+H5I3hPaoxYooTz/bHTKqg6I
vpA/MJnJoTD5NzAKHl4leTaBKAkmbQI/j46GF109zirQbkAqu6ei3+gjVNe2zyOz7KomMFq4IJ5k
EmiYE2PTlQgKuFreea8rzPxv3pY80rSgxso0jogVZnJqKlGBA2CaSw4xUY0C5SlwzC4z/f0Y0ykm
xkzaBD0FkstnpXRv7+sDMJNUvDZNVjJsAJWK8eIG814JPCeE9mKX+TKtc1AvWLDn8xUfqT4XSFSv
vQtnCv6a4J6Jnq1wAcgzlQzCoGDZcTIlf3uGEJDuG11U7wRo4jLar8jk3fCgPe0dwmzgKnsVVmbK
PM4Ej5SMBDVLfJkY7lGKjzA02pIWCoE1a2659vzMW7aKtAOEgSfJ2rd9MZbaLfzW53HqGjgDGszE
qpGsNRZppiWJmuqn5xdC9Sm3pXiXo84SvORgn3uLSsa6Nh1yqAkkEwIniX6EV2anCZNdMmY7HQ5r
KWeUnKUNKEW3CjhyYYoEqAGSSXXG4jk9JXUpyL1G8hdnaRIWv7XTqPrmLBj77iFw+j4ButlXBfjS
M+/3JTO3lOUgrCq+jZFhL1TfkL2hWZj6GK1aG7hMalYO3ptRhzBtGMUdpNwo+9586m/m6bKmQpTR
OrrPoNMQD+HMYuzq0aen20PD/+btwPYfU79ZH4qroCrVDkoqKsuhCVgvMeTM9t8CSDWwHrDJtOLk
lBfchm7OexNM54lckvrm7dGwRgcGTchypl2v5o8kdOxaHy2zZFMRq30hd4gJKImH6BgrBaMUpXVs
iLhBfUzClJnPyX2w3Z6OJ/n5r7eVmyyEohmnBNh7rY87ED/g3tnjE/AIBGIaFJFunp7F4ZVdiMot
4z9kZPubN3i72JO42Qqp9yF/JLHxOJBaotkSA7S9tAZj1ucsmHzJW4LKbLMDgwtn1BCGB/6/o1+/
ri1XD7osvEXjOUDQtzQuxTIEECJr8Q8uJy+ZnQvXzdBb3TtHSutdTsEIRI6btSrE0PCcsLwELnzq
lIhYyW1ca/lJ1+OPbA+RxDTFw1sTauFIUyn3kng+hhdONy7GwVs4ft3n81FbVxhQWZrGekxnO7kr
YR1eKJ6hZ2tnBI2Bcknhwcs0h5sHaQmXFJlVpNzVSDheK9oceoO6qxwes2AZwWwTokaT6yR0t107
I2++KsjBaHaBWaq/SI04dCWs5UJpDKq0Ncd2IaPcLTcTzOLgtzvRqOH6TrJrI4cb+bpocdyq9/Fr
R0b+TZULmtNI1HB0TmFKMobQ49NbNWBfOXQ2Y/mjyXwyK4gAqBX6zQtprbcGY5nc+T2oFl5RCaSv
nL24ozLIW9HdTRepR5U/+EX2fvrxG1jx27Yuv1edKtYHSPfQUjf0cnwhaQM5wkHntgMJ01w3WuQQ
BcSDq/3ZDCIbNRyMGYXxDhEu5y3ERCJ9CXD3w/X6VpaN4Py0GlqKnabAj/NAGqx3mjVZPbDg3b+6
uqdz/LPJhgmVOz8oiW927JLA7CYAYgoogYWmvzXPl25qJdfybAFma5I7fc61TdeIaCy86yy503zj
NqwAOpIUecoseOOWlX1yVrJvTWxAZIW3vyZ81v9JCyoIkfKp/VQa6ZlOnkTSDU+hFoOIbaD9JI7x
IJMp6gfDvo1O/nq7syDbtCb6CmBYR8baiLVDX1cOfM732lX6tsY52xwwANMrktLlxSH4hXpQC5kU
wb63sysynyMoeISLmi3S9n1py0Qic8PUtXtXDOAtuROQyXoJ7CSyQTSavNaRXjH7Ao35EGDy9Y7p
N/Vcr7+ZosL72AWgAaM9sivvNnYKo28wPAqH0qxir30gomIJUSv5+AazGzCqqt1CKK3u1ZruSnpN
dYOiJ06coueMQhylFSbzi90ZfeFCgD/YUSf119Ohh0FOlu6t1pEbsmm1miPWIehaN73+jWp62htm
AornldH2iV7zE1LVhCpin6rzOf87oiWxU+U11Qc0y2yY553bQGZPUHrB4kWMvX+uA9d0rO6WBcsd
rNuu1xlbhmjCgT6NHk+B0yhY4VERmdwn3ANuEARNvHwY8NElCgl2unR+uXlBIoKYuG+xx13ZokdN
YeAsnQRDY+QVwGwsmramhVzvovE9Jlwhn+CcZVeD7YrVB0E7rFZ6abd7nDMlLFRwaXRctF+9tJmW
csWUfOGrqxAR2t56MAfE5Fm/uXoL7QJ65rBNwot3JkcGoScd9SpdJcXIqOOM+OuGWpSuxymNPpCY
hHhDh/wyC+XC8Qw95Xl6aLz5TgWJzKYVVk+OwreQ6sPoRJbXqGvxoZQ90bc0RbNdKns0ihy1oSSI
7TD6RFU8su2uMBXtVvV9Vefjy5eEskGDHHxv3sYy/Jn4WvfybSmhMUonzbjYGzFsgGeJBZDL/Gzo
z16YGWNAP0xmG8XHTBiM67qjP9dr5t3gotf+hT9LhL/yuqTNGvf+rcr7GA9Z51fswtkPBYWj6FlU
04HJxlVApRBP25o4WvygHtyvPIui/+sT5YL4Yn6KAAteBekdXEFTqOXkppY/UhaPmhg6KXAojpRE
DKznuw9rPHYCIAsW6tS/irJY6PH53dZ9ssmd/DyiQKC4n/QoEMSmcQDPDR9EzrHvckx1I5p6Dkcf
T0aZyd0PQrIuwUBLxQrKvpufOVm3vWPq5tBPEWyxTw05zuAwVj6Q8tM8wKaVfXEuCkiHEN/OiZSm
AmKfuVmRotNMgg6x5hsPPxkvjZeHS/tV0p6HfpEpMj0MwB+5tNRAdvYo7PCYaOKmMFI1ntoRpaQW
5SQ/ZUx+Lk3wZG/40tSeH542KehoXB2J9jKtgbQeGjOI3O9fi1RMtFkiWDycBW6RKZn7XH6YrO/0
fYFD8/HOw2gOwltqoq2zgVHB5QGIiYASvC2sZ7vtodKCmXVz9MupQtHA8pU4NMMOXnbNhknTFhMr
MUfjhqn7HDTIRleCzlRemWQiJSdo3Bk7zkCM8LoSlUsU6loy1QsdeG+NR/2TFm2ku3HXjiRRtk02
Py2ZVprxLY+ZexUV3/Wa8ZjhOzduut/qJavxWKXr7aTkNoHTyufvfwTEpUyZBVRaItEqYS26RLtN
toAFUcUr9p+6Q+w2LYN6pl0MvKzwuI2V9h6RK8eS0NpruzSxtoUjDefSZnup6PSjYUyko7vFAfHC
+OB2gpLlxaMkvAx1XZ7GOO6GgfxqO0mrpaCi+9L0lBTPY+gzwNhgvW5H7c6jFCFaLIm9YR2WpKSE
zqXNnS+DAfCFlqM3j5v8CVVFxGkDqXyiwiG37bkMTwx1WlOUIvSYjdd1y3xDMPfK9VRb6/lufv4H
kbV4aGSXMn1kgXcb34P4jioRHcWSGC8+lCAQK1jKic1aX66QAGC9eHiuXQwYSHt8Ic6hdGVPSSC3
nXvk8ZnJmJvdvwLp6rCDZUwtltuh7QGiXxt2B6lQwEuY5qhfOZ6DYqmHDua4fU7FFnGz1o+48Eh2
XvgTgNAba9k5kW0W4F6AWMQTeQ2yZL7/hbUtnnD1B7ow0J4wUP3qLVyu22Oz7s2IN9PNy0sBaHXF
3h/c37R4tVUJuhKUxKkASTWDeowGZIwjwQoTe01i+jTMRzL6uJclHhRmS7Rlm9E4svpeCZSC64+y
L3ujplc3EE6lgX+LIst+pOclucN14wpQxMiz/zkzm4NZwdp+XhhJ5P+EIoSM1fPyPoVI0xE6YX5O
sOa0wjKOqYnLnH4iDiM4dymFVJYHgRDa2WVVT6Ozj5rtMDbCvCItkXliGfTMrIMWHPdh3JgDw1lJ
Aiv64ccDfZ3zXksiJ4bzdClTGhGFWDXS3hAiV8FAbjL0k4uKJARi3xxdYZobmmHnmP3ss71+9y0y
giA9xseyGVuSgELWa+9PiZSMnC/0PzMBHZ2EQuljnsAkQStVtJFIX9sbRvE+zDceBGE3Iq5iSNGV
VFZSMA2eo8ajCGD7WDCh+ro6oLRxYqbuMeVY2dDprCxoHswoNj4zkgTfOAmVDdQHri7R2CBQMQ4+
dwbCQ20UUVdPlK0p0lP9ldhO05LhH8mD75zUSZh6Mtqq2D0JDMi02rj8qPggp2Qaj/TONBxqzAfN
NV6ikNA7xk2vytDUMfWj1+GILm1d1TMovFeSGBbKCdX1hARTZ6voagLyO2kemzN2GdLqgkmxIjj9
nMShyNi9zjKWVfm/9edLwKkETCNGYp6Fw1XGNX86my6/ZqrsnGSAEAWROhoNyAKQm69EZUkeLAuA
vvhpE0w634w02m6kBx44zTAdmQ1fgxNMHCz9yA0PRgiYQORmSnabvbh4at6vfu9Den5rIt0Y95hz
vdgyPTWXOcrpKiieM62BO5KGj3Xj91CEuRleF5uorVMLv7BQeR6xNkf8c3ltFoCGLsto/XZByCns
krgmVRRa/vmDtCH4C9FjLOTR+T0c2kkN6ERnneR4b11O2wl5eKSAiKQcTob/6Oq4WEcbZMEqkkoW
5VLcTDovyQyi2YV4bjj4Chrjfl1TxWvdKAyzID9+3YEw71dzPybxockaG+BQU/umWM4lhp59gy8R
GeqI716/1LVJIMcKiLJUNiSCJKXcpBfkaSWSqHQQJWHH5P9c2jfH9exBRwYRLLmy7ssSIX1eezxp
o60Ekw7tSV475mHDa2Z6X9o03PiArKyYog+OWPfW6roHWdwMPCG2XKAuTejXktrOjJZ3p1rYPsg5
nogRBSQSGaEwEkh0Cg0iKaleWOujizbqJBNH9NqGiNH3Or3cPlgPluEP5exZBKsqzBtJSZBga4wF
zCRUjgfNi0Tv0j8V3/3aPNAw4wzUNsFsBkEPpoZ3Ih046PaUYXh8C160EN9eukKhokAqHJ6WemUl
hlJDfE7nQqs25KHSfx4+4aotVJXbSCV6ffvZxjmHB/P0cOwBJPhMeB5LlsrGuschKI3OjEo/QRa1
2dd6w1PJu6b6Xs5i6YY6c0xG2FuyqyD/axPTo4KCJHFYzCM7oL5CIqOSNisw8T6UmCogAmYLihqt
8nzI3qji0dqQtNmka2fMaYg53oSWHqjeo1/BpUMyWSiIZDYtly1GVHh+l+d4hxaFtfRVlbhGe9wS
PB7TKKkZOP90kQp2Ut65K7Ni16uAIaii141Wd85xNkUNqYQi824WJJqh1uBwyFq2n/JpN4teSmeT
HNF1csQvP50MunqjKtjoQSg1exI33ka2WfeCF9t9pOESbWY8oBpfYIWyg7GIQk1gnCXaaOBh3Wl4
4lzxNPUdoMxiEILTpG1SlVWu7cKFpFhb/YNuTkmX954SNa6C92+aa74EpnsuMwp43QGZpsHZ+bD1
JaMYn54+3AED1A/LSlgnWWIgiVoik3dMEQuRLK1oUReLDhnqL2qW4lFF4AgTs4iLutoyKy/hAh57
pJH2bXrjV5TAz707scDzjVjvByWUqUYXi/5VjfsR5qSYySCDVMsspH5VZpkCk8RVhpzkfpp4UFIa
tZOsYZJZYWuEP7Sc+dfaGWHvRkRIXbOsf4u5Iho3Yv5fwP4wbqrvVq7WMVpzgcWoWjTgKb9SAC0O
b4a7d0sDqYKsNNyRFHo9E6Dg+zRg2Nns7bZvtFXDj9zTyhvjaVJzdY6BenzR3am4/mjj6EtrY4rM
KHAr03b9vcSy9Ac10IgJkNEEKZh3dVZ4FrA21xSpI8EASx0D+jR0/AG183zDAOv82gAMMvwgeLoF
Li1i5aQ52yBq35sgyj8xBHledzkG4Wx2TIPbpeJQjZOrXEZSgtguVmGvA5gfkCD/mAfi5RSQTKmY
8PWUmPz3lZV+PQ9lh7Mm1wNZHYSMY8paGgBsozCoWtzHWPLAcz10+leorXWdDQzRV3rylc0tN0jt
lKDf+aAN5I7eWDRHLQSJkwCP0qA8N96dPpdkpthJIEDmZ8rKh0ag+GQTpG7kmkhpLnVPNCZI5m0B
sv0NTWoE0UcHGWijR44SoncXGpzT9LN9GrE71Rel4+PzhJB5J3KTzBuwIjq906cKN/Wh/l8Dunic
zwwrEIxjViA6mzhryIOTaUpwMKX4KFLZCmig5TIOn/L2sVFs7+CSRy8rWoRJTvdVDoqlqYkJR9bR
10Coy1fLEOKfC4RHCzIj6Mk3V68tHoNcklThBPOGNS5roMvSy57mmOGDlPE1/Uh9OGNM224nGlYb
4c/tjgoALTvLZzDp0mTtyF6DurJbUD0zUJly7OPkxQD+Xv+H/RgfEvQbO/7tKKI8WI669zlRhOrU
j0DipnxG9bdiHfha+NaSzeKM1DFwBVc4TFV0Qigxw7cwbIZChtuL7IW5Du8yaFYLXAE4Ubm1JIRN
qYm39X8+IS4Z9GhbsL2ZiPi3+1Wdp/tQ7s5Y8Xgm3GFTv7YrmKg8B3yipKPDohQJkPSN1hKHTec4
62+DKeTag9LT70Z9wXEUfTMGX2XqJYw6DahYtICUfkyol1qCmGb1cBh8DSC4eSOxmfUrWbsVTHG6
P6WIkynT+UV+V69NbX9o/cvUq84B0kec5nk7oil11917Rhwtv9bZkF8i1NSZmIHuI7gZCr5y2sZw
DMqRDDqvKao3TTxndGcydRD/WrORp8XP3ijXWDzOSRJiX5fHr90uE1hHiOA8YysFR21jE2j3B2re
kNrukA2IvOtY7gJn57qQW4O9lRNzwFrtIMsARlD2EEO/4JRUR9oh9CdtDZZEpT6LSMybi5hNXjiN
BOw+hOiGa6xCo4BGqhLLKwlSxQN6PSZKdYpryctPDUFfPhSki4pCsj3eHuXuBmNI0pqhpkXrNGAQ
nOveUd65FAznbpxRRW0btDdZ9T4hDu1be2C+/R+0Ul1GdJjymYJ3LTqZUI1ytu5YTaGkBaZMykoN
E2gCRcWgWeTgy6B6Y0WPt4wODp4r0mVhgaAV977hp+/jQgRbVgYXZogSYPy37g5AE3uS4UqyvmEg
CWWtEALKNO5R1oqF1auNAsilguOSIOb3gHJYT4UDd6tC5IagRZzQFZZp4f8rg0cVagKKYn6mOCS9
Bey7GbuvuFuZBK0OtoadZkhh9sbq+5gJbiEr86h59ke+PtE3Jt8v0Z26affpOoY1oRpEe+P/+FYf
gVgmbRDoWfyhoyCj1133st38mwoeuDVkolDgKukatTQ0PdgdllXJLMP4KBaEiCatM3OJcEVYVP5y
WDtK5YmSY5k1Tf3aYNmE3r1pzzvBEUIyEmKF45BVESmGkVuZ530P9bgOkMzcZwJqFysKjlc+YtM2
6qncsYW6Smmoel6c/9ysUe9wYskPxyAeG8KsEEu6VoW2VWjkepCpSkm3ow+tOtZB9faMf2Lv5D58
zjQLIr6PCnxsABr/gMkuQWOeUttH9IY70xhok5sA+kSFFxGvMRrvX2PTtLpq0hiWEY6FhagdJeFa
AFkN260sJOMDLnVF9Flv2+wByheb3B09rjWEbYHxGWn5cMhjlQzI53JOgfXOwaTpT/7U0sMXK/OT
hrKBAJdYDB4WrQXy+FDyHnPY4vz1jIGjn26NfJqqen/iixJEu8HhWDbHIZfa2ZsxjGojQxTBLQ+c
veeLDdKbY388m8a4VVf+E7ZIO7kc3Rg2Vd8jBEtlpr52CQaUS6EsMKOxDczIyhFHe5hq+quSX3QQ
2utq+O7Zx6M8KTt14Z1Wj5B8WidNI8Vyo40bg/vSeyVE+iFfWWEoAjKcr52RKZcFhonZJtRwRtTh
0fhu/wsrRDvV7gYTn06nYQNoO0ae2qpMHoM/8w/bMH08r3DFul4WT1LT4UTo4vIvKKCOgRTQBCOy
2hmHb0/AGqHxX8lqJgUaLpreWVwqeUxztqjQ9P/kQU1BdIkHsdyoQmkBGkPpB7d03opPxlVZWN3Z
q07jajc00x4G/UboYe99FVPpZ/zUxmx0GnO7QaDH7IAbwH4kMzGMjcX4MkEvFlcu0UlZl0dCwYzg
/63kihu3aUB+75vjhqlZBkz0Z4rd/bA1l4xN2JZ8PKkmUHPgVzn/b0JuYInq4JpXjwBur1sr7uyz
iSI6d9DmWBmvW7MDHi/nT9bvq6rEpHoy4DdcTtj9cBbRb1eW6aJAQqAVeq1ejnH7fq9RUyVlG3Zk
lugWEFhzsHCe5udszF3d244oACCF1RmG9Oh0ASD+38Md0r1RQmgUZbeegA26XRef3p72lKdn3VLG
F3XzelGHi6wHSrM6uAv4hSyVDNa+vTV1WBGQ+ufewIq1APwNKwFCTjuQCNzYRX9r8OURT9gq7Xh2
x2dFuMqrUnoDVMuWbMxUyhhIRCMQvA/jtmQYa6NaTrf0mj+Y43RySi0ZYgNOHMITu9LqjEXD9Vb0
2kqIfF+Xr550mtIF9xRYueqJ759cUFdbTUD/3dLXTujJS3N/heC7HKDQu9tL545AnSMEf+zi1geX
BLiVZ+Du84VnJBOqTT8bRteOK2DSRENVk6c8EJDbB0OswLPsZUU0XBkYu8kBH1Q+fhatqwOqEhlH
Sx/m6AYk8tw73aK4ekBPm3ElwqImAUeKa2jgtVJYlGS50Rxqgn4D2nCIXO+nqNUkq4HkFqlmwE6g
aO2ii/YsAs8isXzWI3BNjBMEzBE7yD3PB+RsuyQG4IYBQVZ80cOGhEIFRfBubTYwKcrktEhjW/bR
df1j0qmzx1uWzup9pSoQWmH+1sgA2pVBVUt0Rcie2A625GAuXF7Zf9psV/qj6jscYGDH0M7UuYx7
+3Pt/BemCWhNWHus/4u8UJESiAxxTNOfhAhNYzaV655s8U54W4DujWWT8guaI6UOUIkANH5gN/Nh
m8AZNrvyVU5KmIRe10DTv2N0WaM6nZAfbOSEcGu+fID7MV4Ro2mBDT9ICPqpug0jc5Zt9EZEwliM
pdzF/V4XHdSECppYOUS8bfJlnfLPUfCUs1iuI13z2hJ+1+eG9tnCEU8Bxtd+VF/hubbnXnPdMWYb
OLkslfP4VvttF9FgLkrOC899IJGT5MAL5+sOJalbs2aX9IbMPmEPAUYktWwINjxVEUBmZ1Rn2yTg
bh373fQoMlw9PyofLL3EZl6flyBKfvwjkkqmu0fxiTqH8MU4KAHKvlFYLRAf2nmvh1UTbUk7Ldea
7LtxvYbvKrtZBzafyBJfXeFSQrQT+FOONoHF7NuQ9kyOgSfiJZpb422fzbi320K5qfm4PeQYiRY7
zHgFFaL20vhSf/K+BoYUmqc+ImAzr+/tfP7KEqcx/ZKCwbC0tgzSbLCkewsMTMPsEIrDTMFV1rJj
SclhwCPQTC15jKQ/Oj8ZZzNK6NhDRJy6WWYyNuyVTZxglQDiDcWzcU4LS14GkqBLkERZ3RYvixSj
zAxODskZC1JVKS933so7MfIEeVGB48tNwgtxVT88oZIvM9Q1ATUVoCeSQ0DL5QkSMIcCK2R/Z+BK
e6/n1hSvx/7fi4kyMy1eWtoAQYRWaicrsJ2mOqvbrprls9M876Rqd5cn6bt/bQU6jwxMZBfYo+ky
XKtA8yqC34cMejZc80seMEtky5hKb/iPLkMx6H8+ZCotbAYkbj0f495rDQwTH5k40u8IyY0XdFLw
sL+b13ZmxBKFkKCWy4PjvlQdJ5Za6BYWpAZfDZWV2uYoA1w1bmZ55wgopkgfBdiCSIaV+clEu8ft
aqQ0qN/8Z7ndAVemL+SimLy5T13x2cl/b8HzmHEPM06XjfSWx+7mXng1JxTKdzcw5yqvxBXuNqOs
WjPX8TF7Uq3m96KhVnWo/CwAEoqqzndICFtuctvKPqC4Ll+3mm6ifH86cQraaTVmBd5pNACbsgwO
YrwcMeD9XaVVTAEB1NtCVDgMvSIFWjVUh/gZAL/1GKcxxH/e3U9RbGHfY2sT2pEFZ0eatLARjLJz
5fo2YA80mqX0SggNYClTfIqv50XOlNUri7TOLTn/yYAXOpVAd73N8q6HoW1grMwzgkWJqbaHmVTw
/FAmyzgJwlecA9JUs3s2tkByZsmbDcB7AAdsgBJ0o4UQFqSXQym6AJjdtEtkxRtPu0nmJhWrkSMh
iUmA0T5Zn8GZxC13cFe0KOtMLodjU3Lnne2r9qgd4bTO7pXYH/ig19Uq8Qwv/osAabb9edGF7tSH
hemvu7a/mS2CzrmVaT7gZSAHW7MGAxMZQAh7QPw3G/45OXAw9ucMsiZ8zX4KrkPeCPpbTXUpvNAT
QcaimdeyjLDHr9GBqlTDDOoQ7dDJY9wwLDOmoQy95x38Slshl1lFbJZqoTFBeNN0oMgPIsN9wfMh
pnbXV/hDPqbf3ssPJv7OcDl7ozcwmgwH76SyAoyoxD4Jqt4N2tMGUCs18/rCtlYcT5ILLScxJ8bW
ERha0f//M5SjyR+J2AqLCaJMVXujwMzg2lGzNofy7QwSYuqdN19YUKAffBDnJ0TYm0RmfAvxaXsm
2+ZvhAg94U+flppxWzudNLtdM0rCUxJXGkucQWAganGEFIXeoKGZYtfyvaIZ5u/dxDk77YsWBMCn
3AN68FPK77+rrx6hOWOjZEPJ+8xDzpTEOdO/gZzR2O2m7wPlt4XTNKDWpp+7JHVR5BNWRy5SXrq1
ZXsQ5X7EJzLusMfrKqFNIX5BgOtRNBIYh/TC/f3y307ihZUHNZ0pk0ft9juAk47TMdDuT6cPzacb
HTzGCwJaT5XkTqp7jOgF6/yoASQsSCRRGLIHKL1iUNh6h36nIo9cBikiJqhHIeJaLT/26R3HQg6N
+7gpu6Wxs8JJu2OC0iMlJSeNqiVQpPm/JcnrC1TBt1Hnqp158UBzKUIRJcKOd4KmJgq7wqLt58Iw
Nk1QqCzjCD7GUslmqISwTl60XG0RcogMK3uYFEpasE/My60NJIODA/83ro6mvaYC0dFgv+j3DzHT
83p51lmFU205o36pbm4x0Enl6Asr9xoVr6Lm0SzTI+A8g+0oAqYShPjtO7/icqNBYzMnhD1QvJ6W
WeO0xue7jTsq0tAm1FvwDeKYPCpzcLPYsxGgQCffqTrm+Fhhqd1KP3vj53Gwjp7qgS/beO7S4gwM
UoZnY9IZvp//2Jc7BIUg2Pfr1K2GPv7ACGb4vHyv1YOS0FVpQhNvEBzugvDK472lR3s+kA/lXRj5
bIyLbW2RHc6kOymEL5sGH+SuD9ybkOlrb27euUC26v7R0zkX6z4WHXzWkuRGvLdO7Yew5b9VcX/I
eZ+EuzoGIz81eo4X1VMmXTnIKXkFvy7D63KXrJGBFNAu5aOl6WjNThv/eFU+t6UgzeuiFTHK44Wm
dCDace8ZIl9zb/nIt40mLInKLn1QOREU0XV4qNds2+mZcNhOF0MpYxViweo/fJ4mvtoyOqt0PqJU
cxSzXJXvSJS9o1Lzd7UYwSwPVCH+nWZXaDROrgbDs+MELBcdIhdFYMU9+d7H9/X0SVUL40YlIkTL
DqDVopbhUhsTze3Qp9ZZJj1KTpO8sQTouyQ9ZdIey3zdiAbXxyJhkZiTJKSoFlJrqp4C0lnvUgKv
nSDZSLYZoFBdb7ImbbpWMy+f4ruqWAAYuOspWl7oTZ2Yz4KougHoxCfJ/7MgdMp00Fcf0dHlV5s6
zV9avSNDRpy4jDzeaUB4xz5MVbXGFxdd5LO1JyA8xHwEaIXRE6qebL5yXB2qWGV0+rD1gOdpYqa2
BtQWuRwCKkLsm6Xo3ckxZ98R8XE01PUBYf44VpyfzhXNkY1mCFViOIkz1V0HhcgjMFeM2DdyQ405
3iDVlxZE0dPC//ilv75zVukcubE0rDrqLJeEMQCy4raaxq199MCQKziFP9yKGPKT25exemM6N99G
/AVPv6OsuJQx/b8jPFruH2jcm/CVUfliSATCeHONcZJmFp2gNpx2xRYR7UPSZzlVaBtO21/biuv3
6Sg8OYvNB24ClaXI00yAwO85M3+Ku56JDoEENLStTEHPWirkVv+VOe0q4U1A+OjjhJcTewCS0hay
kD9l7U1jd6OmG5RIF2FDRBDk7aCkl4dZ2TiBRLifzNjQRPXprWqlBjGe0qi57hBB710S2xV3N5Bi
gf+CyOble52QL+22bdLCBiAYcdfrt2wG/Rpqtj0z8d8Jn3CqabaKRzskubb5/nrYXXhBVVX8eceM
MvmDqY1gStiKsgEjmS9uJu3uHomTl8LVAPx3KIXClaig9TFtDtJO0gs5VBVtm61tcmP3fsKAttkp
oZjdtT/gwUWu1kKinWdCzfWxSkH0G7fqIUMQQY0s1FWyM/gAf1a3CGh+MNdqMkhlWmavrcu4K7r3
nPPShecp/H70+zR7A4CM9ly4RRvjEXJvlqzM9Vwtq23Hw6UUTBwyJDEXd8nnV1pQ4rpagwl4pLI5
DbYQ5QpAE2x/KszPdM7FwQXNE/3e32AmqmEgjMFCQgFUvqn6Na6Hp5WeSwKKGRG3GwkwX/ersQd6
7xsPjaxfE6YggxQjlf3udqRYQ9w/QHcovu/RfZetKc1dZaB1+izkxBJN/x6CuPMbYFG2BNGphmOq
S548uG8TuThfSlms5Bex7uyUIMERBIhLM3x0/X7XJzJnMTMxbx707CvxdsRfg0T3BKAxnQmHnZkl
38Az5OB+4sfHsTosA2EhjjXdxFop9of90DScq0xMeDGQxwa7snEP99xe2U1Qumo+kx9jH2c7LKuB
TV+hYtfVca7Rof6wWfutxCmxon12bBiget5QnsaI2J9X6nD/zJWrshyitlyRGhD4IkkUitEmll8m
F2ISpJL1FHXjSonbM3NBkFf9oPTw/nrSA1orMQT7KxJOSWwEdNUS2F6kAhhL/gmk4M7P4LjAsRYB
d3Fcir4xiT/ak+0OSnDLpoAycKq2kco+FKTg+piWKiwUVF/cJzbRtoDGZfEFgXpTTDZObHCjBOwl
tGhhgZweWiF84LR8Tv+sjrSONvQcBYHei5FRbGvpBUwfyYsGUqqxNkdI25b4bzyRdkbRAJfZcZLj
4wLojO+gMiJiQCLdERS/YfPNWKUeST+TfbZGUiY2Ee5BbWjaF7eMdUGf+aWtQWSmQLICLwk5760C
cInq1SgtAV5+VxUE/mc/1PKTHwRxLaKqto2nUSpL/FpUqcmmAWo/q6FxVBlsbALJTRTS9eQYeuNz
kTpcLZIFi3Vt3meuwZ+VPnfRQwDCT8tjnwp2Q3qIb8gzUd4ibO+X6WfIvN3M8zK1BoQ8Yt79ThN4
Z5fM2oidSUIQ5TrOuWz2pwZH1QVvYVyCdgozonvguDwJsiMjOwKRBGIOYkRidcu5X0iYq+okBPCj
loipeDBrnhIInOrHQyzViF/+SYSzLvrp8uCnTOb5LwZCbwuEkZRiHf5GRuj+ZdD4EpemIMLQtOdI
sBYk/1Bw8HEnKVpdJZanzhWvM0FZEd+U4WWnWfjgTLiMoc3ntEOdZUiGE1qCXuvLw80puTWZeVjb
LwpADOyOJtYvKoHJH/cD1IPgGtGTjT/vYBkD9u3q6XxS6ropn9L/INYAxczNPMUyYM3d+E8rREXV
9bJoOnKy/OBsLGQkBv632AysRt0a6ue0uISpEgKNaBTCg3MfB03pPEkkipfxslvYb/iXA5/U5tVN
xNhUFA7RJJaszMgCrG451D/DsWnfZvBX/M5sYYjpjDHzTOFOfAYZsHjodyojLlEQn0y4hypdxEcI
WIBDJNIKvbwxiapNfnL6xxlnuH1uXet9U4ErXZ7+WT0JrZloFx2LLTYBPpFilugIzCWAnxwp3XU0
4tpKVWY81fGG8Qzr2zE8m532ze0xOzgsiVHlGJ51HRu2rWSqKGyvRhAYQSnXrc6wNRDKBhJjJMfI
azVKhnQKAwOYb4crvMgWNSpFy9nE5pAa56BSHraAcK41NCNORliJzql96p2K0TvwJePidRpKh5aK
0s0ltItU0rQGtc4Dirg1P1odAz0yN9/rKGO+1g14x5Q9KNlV/jJtn9zWRhCrwLaquDHetpaGVxWy
Q+YMcJPR1fuz6Zy3LBC033mKXsH5cyOJ5oNwNhunYrpQ7N92C3YAO3au4AV5iPTvvRHLnN8XWQkq
jTUujcgYl1Rv0HEEgcSDyUB+gPZ3wk9IY63LZfM3fGD3GPhCoMqD2WTCVM3IWljOAPkT5YGiYRNK
PJRxJs9N9OQluys1bQDRVsC4mytrZslL4jL0MiJLUvxuyUWOcMEGwqvTQ4Pd/GvFDBqdF9w7SXoC
AyTLpadyaoUNpwNwjwpvHnxZpXfWiyL3WelnWNYiXGx7RZFUlsxHWlLLqMRpXNNKnhwDPFdhbAoa
4XSfVHTBVtfqdgewiDHR6ivlY8AMvXDVoWD1LNIDOkXdIuFiamLe0NBhtfaIOAcOT0SDZONqKj3X
c1XdQGclUpnPrelzIpyzyibxh1gyGV6yXrl2gUdxX3wU3SnzvCpLu/m9KtDyjFuQFMs6aA8Fr4Lm
XPty62gvYYMlPL2bxnoLidctJIs2k8AWdkbNwlWYSP2p4WoepOrIzfhVS+iwuNpEIMP5nOt/1lq+
44HDeLYGnU7jQB8XBlPjQCtYdZNZQ3KLRJrSICgUck/1ZpRdj+uF5H78H+9PZgxkGFLJ8tlrqBF3
jJjv0Nhpdahs4mJ/vzk1I7K2lHJe0t1v7sqCV4h11dmo9Xp3o3Cw7dIfnbg5usSm8lGZjQvWCtya
opEbkeXO8jQ82FYAQFEB11uGtZk8SGXfLjqoKwT9mPXJWYJgbuUDkPWm/6OTuApKdcvR9LFvd+SU
ySzo5vLnUHO48rtnCmaIKppWFonAC1Zfi1T1T9jABWr7h9u7S2RIwcnL0jaFeTbkZxO5Pm3xsNDe
eMSWvKmsNJAtsXGm50tSHZXAIuQ4EXNjLphz0n/3i9cRH6wH6+K21faUE2SFiqElzpRzWs/Z5Rlm
+TRFGWZqzPA1CnnudNJL/qORQfJhXGRmTGlvzrEwfgblBsMNOcdDDBYO+5mWtulyEi9fXXXVzCAY
0ctNgQ0AqjW+dE1q6tKZbu9HF2ZZs5UkAA2VNjlh5NObNEfVcI188B+tG8d2eYSFC3+uAV4kqyx7
pVfF4ATzcHYG3/LBgvP87VHCwL81YGFXbLr7Vaq55IiuGaFHEy2ABU2ngLop8XzGBhqtOchWmrjV
Xl2FEjpV8lhZVvv8O5ganTOFez+8P7zHdoCmq3ZWcHLzn7Ze4bWKYDO+t5S+x24dK56fmu9KluRi
Oi163TIFcFrY/tSNN0rc5s7r/uXy4gAMwnVka98l3lI4S8rcfzQX3NmDPadXaf4OP0qGZ++oB+pf
GB24dROyO7W4bUBRjg4G0HLtC7lBjaMqWFZZoGh8fzAD5NnYNy5P9WqyQzASDvA4oMNDK7DlrbfR
XmNEFV5xbLOAi7W2lfSwm0XUuLlKvu/gcByO6jeGgtdFpTGUV4l4mC4Ts4og9cBJcZoAqB9Agn5x
0/aK7cC15/yHEeShzGiXgEbE9D1fcB+6dNcpeA6ahJzNIscElMqBLyM42jqUbXhX4loqBv/G8mQC
mpbX3OyvQSS7QOlAl0uRJzR+xoEnabmyGNajey8PhcsykNZziWPuNJ/HG0ht77DgcAEjwBBn2HD9
0XqYQPuZBURNlmNL9V8flqR2pVQvggGStqLxZj6BtJE18qtQq4AhXYrnAHvQtQ2kdL9yIIRIJNc5
CY7MSWAZO4qV3C7o4QK2gaeeIa2ma+2aybh/mwlEuOffD+s7MV6tIcXg9oMdO/4i3T0+XYabrXAT
p2CrVhLV7Bxy2W8jGgDgbZy+gWY6+60xoSkX0AibIsg4Xvq4BljErsTehWZRv9Jz79tTiH9ZlYFV
kDuqwTNgBui+4cKmC2fwALQ6X1bdZsb8+vlOazgTz5EI/put/yY71tw381B43FFTqnT3qSTevOj4
XpI21c3bHxD5feRGZvoQmdlVQ/SwNSoj0TKDCgPp6OM1uD0ftUOTNQUsLZdZkaOUie/6eWNmqeGu
+zV0fFvzXz6dxpD/vPFhzvmmuzyvmFSds+pYAB5sRdUo55T8fWNt4swbml+SQSBRFqHzhHcuOVN2
vJ3ggUHIBRXSeDEsgnZFELbtsawU9uugeG4vPXMwWB3LJapsSk+GxDNIFZ2Vi4VcP6zJWMrt08wA
qf3UNBD04BC8juMWEMzTiDHGT6DXdXAlmoazfrZ58OZX2i9vorsf1uSgp0W8PjtXBq/axtjUO7L3
o8pehtW4dDHwGD08If99ntUKZmr2njqTMYLp7dR8otP0TVHPw5h/qMgiVFSGgcTmVjdbQ5baZLZE
okHoD4EDZ5hn0AFKy+S6Db1/wkkTIf/rKTd+HhoLZeVFvu8e9Y2h3BNBBYhSBFa0mr3kAkkwIDlG
V4Jst63JkGXKgbWz4SV6cqCcna1DUmzWNC66esvRKE6kRFP32z7HS1npcbfbt0swy9HlP7qdr4MP
KLdctWPomCYgNtdu5Zq6Paezy7Du/R7+iPN7golhRZKmzilylxrqvWVvpwfqD1tjwEEjX1+VtDsZ
pJJ31oMcqhha/Zlo3NBEyBiorivMPzUk/8uUjGCh9ImJjgq3qkxltQNdHMW2mUy0WyhDuqVs3gST
2sS7CdwvY+oVb61DSOJ8dYhJAePsf6+sj6mZHaRQo5q/4yDATaSfO8iSzlF9RWx9S185wipklsu3
0SMFDXPFMGiUkvU0BoE71sW2U/pfWrjcTsdywQ3hWOX9uAfdPBhkW2HSkwxIpAqUPWayePvK1xI6
AwPC4E5a7NWROxPYHqvVYnjxdUGdP2sHFm66Q9ehid1Og5jZ9KqCKoS+Hn01VETUBy5P1s30/och
sw99kJRzty1mw5c7Pjm8Q7lbyHztp7INOCu6KlmyNA50m60EGwsBaVGFttlgqkZOc0NIdR5cuRR2
9CG1hh0Pu8AKzybK2L+2UlQEAXxcDaHiLB8EmehnbpCisysHSz1NpxybpGuL+j2xHl8CwKezNgPU
4FOVyqgOI3xUD4RbKZNGgEa5e6SGgRSniR1a1Hs2f7ELI+3wdCGPIUNZoBqtqPbjBSKHawdc2yNl
cSpfe4SCN1EF/5PMj5UPRZd6ceqoAqgRb0xia9G2D/XCfZHsp1o5OFGbT4BqE2aoLtWSksprceye
ryp1LK//CsZQ+09VodIlfO3/txeEcXqgZjWWGx79puwXBqv6Zgdud/34un8R3iB8A0XVwrgf/b4/
wkR4/WCPu1l1VMU4L1d/FQNAiAHZ1rL7nnDXI6jt+QmZC8as0g2gJzKmhxwsE0QTGgq/m/djc74+
i+YU2uCWda/fgfUUYLaxNrQjffato8wSWQYdLS9ZmD06xrxmDwmYzBQPH4lItgo6zzCLJQPyY3iM
Tlp0sf0pE1ruNgdQ4s9Ry+LV7oiUU4CYoDnNL1aDCjJTlktILYz9aa+EQ1bWIM+pmidTy7y6hRO7
7N0iscl71SLCoXkUoG/m52cxhvY+lusMKYy4FdXlcJ1BPZvOF6v9BlLr8gCYhzTNrqargq7TWjeC
BCv9eXZyayrQ5gSKBTfVaiQw7z32z3MUwQQrWTl7EOtaNSwCQq4gP5eqQ5i+H7XDAcY7cuzcbz0z
U7t9+89PhIaavu30KGeKc1qYvb/fXCnvxKrexsiFdKjWWRUfcdV/uXS7CGxExxjGf9HzRaomD2+B
GSRvRn46YQQiUPaW14zcUH4QNKJVE4ju/o0NIv+FDOM6M8hV8pEpscglUZIjGu1L4jZlClIAyl5d
rL4d1vSuLIUAuGsG2CLC4o2TDf8PDFgx+aADTc3+VHcInC39POS7tUIGFqkDs4eh8d5ntq7spbpX
1gv5vvSu6F5eGU7SdxI+rUVFwWZNFgChw+kVE674c1W+VDJiYsI8m12Vf8c2dauxhwo8ebZjpHlp
PIX/HEnN16pAIeCAiqqJAfwf1Mv4mxUphgfcxuvO1jUMrDNrfCGxpC2CIg4AGqbIOi8fAVKRtJ+8
d1wf+h6NADvCZnnIb9yL0y4mU4j8uo7itsJoFpgXmey91uOtklU/4TR883Q3bMS4mgLjVcbnGWPH
tgGiE5ZHzGnVn19GmfrFPW1fRPckakiJsNEnaiMg4sOuRNRWZm5N1dTrraaXli1OIU2KKFAuikTn
Yy6nVrdI48K2ESoW7lliX9lNZ5ptez2OwUzm18TkQc3X8eA0wluK/QlVDhq9Fiofo93qAUsA6zYd
AFjgnJH7nPw+Yrgf+vcMmZw5BgNxhz7FjvzHNSnT+LV96dI//viEKQ8V0PuP1s2RVMGtSY3+7kWH
Edl+3b6BmtbMYt4yx13VY0Ad2BLixQci60YadaMheFNRmeouzufCZq8zchA+c2XLWMnFtITm+kUm
rsYIgfcX5nLTeIRP3brlzuhJg8rV9aS0ERPFt/QHO5eDtCf3sWcHwW5Y4+tW3K6eeoS1tX4C+IDt
cEEqFMQyqP9sIj82mNzC0jEpr3cOfFnvzCcbIe6HymlK78nqSaY7zDICYkJjKVbJouIeOScCAey6
CPV6Jwhl2pDxZYMb2cEzUYX9WO40koUp20C0qOImIVXj+jWbsq6iBS3Gn8kSx44gcymf6AF7MCab
HN1Q/32xtiFwSsgcpGOstm1lSNR9z0SdQ++szjWb9aM0bsjtrn2jtzVwoq71Bg9t84r/6EQUvmHh
Mr/8fc2LpuZYUdoyLchB1n+cpFGvJmUw9U284fs68s5CyNlTTj+g9tSvmJn/A0gYNLOpf+FYv70f
axwiUHK+6UnL7qNxJiVPUkz4I1oYSHafEYBqSo3V51XDNlvO3isGFWfehclGCNs4eh/MmA1d4STT
rUaVuMQrq9m8dA7EIuP73FqZA2LZOHibIIkpAxREP8gzgyYrk72wG+yb9TknI6nXIKLH+DgsXBHS
2BATJit0Zm1LUxw6y0poWuSkePtyaIqeKJmOj/2jsY7+q0xpKNEKr0qr31dRFnHDZBq9lEya9PDV
5/+qfTtu7udRduCR8URl5Fy5kS7Zs//2nsR4DkKJ3pUrjf29s3ig7RQmaeLhVNB5cvL2e3t/P6B1
FxFxrIYVa3YgU+UVrtSCscaeZ92H0A5PoAAHfDrKEtcWGZniRarkKwFntzBBXH9DiH83RAr1zDEn
LKQtEfoSACW6HBZg1VLGRDDgsOZvX6Plvvf92IkhFHFbC/a7IV55ErT43Vx51ClUyL9hHDP7IriG
kq0KHIfAGgm4Bi7n1l2gGwZwTgZ5xvT6+Yh1PdHfkuZnBSR26So4v/XosOGFjM7nb+Zovqawtd7F
slmCgywEE2uwJ74YLeoKz0McxAY+uGpJp0ro9hYnj9HruDHJGBrIOsQt8SprhQHu/VQhcxa/iytP
+yuRr6Vnu4/9VlVLmIG4iPkVdBjwprXv5LuwsdYcoGAD5ntVjWRtQ+sAVD2qOzPy5QR3+q64S/Qr
ZLZ3yG/Ia0ca9ZGLJyeZTP4+tO7dm3vEvzuZhkzCx7OdBs74rgtebmA3BpEDyH4mLziMp7AGDNuC
G76Wi3IdbnEaC0ZzfgU6FPsQRrXzkx4GHpIeuEWGFOqcZb2QIydi/i9r70x49+gKAAVIHH+9jN3K
+THDSmmQdtaKYCNWMg9eDUrkGZ7XQGObe3cPrcEMyOZQ/VR5VLiHrMqssGQE3MKrk+ixCC6+YJGi
5J+4c6M8SpEC7rxwYPjE//xqOEl4eKQSfzmErDFV4FOtJI1TDUfYBCkW6VZNBtlNl3X2OdAyVxeI
JlWZFnftSDNgDGJJ7N0g7qMoYtTUXN285tECEkgsBvBXAFcUCnBACbKVdp2tIBZAfeX2uw5rfDLj
OGKDeaH3Pcj+kHinaHDsNqB/Bj0DXA0NSjXX2Nmbt8xYrHDqy/aRadwl7V8utmxDi4fkb+43x35N
xEDxiOpNcdcjBEDG25BsnHdtxcJNc+Vd2qXabmsao/h2isnxj+bpWMqLODlkKpZP6lgqnym1h/vV
cLfgNHYUUqCARGB7U+yOpZxG9fu4qn8o50CosQY1P1pwe3LsMlsVIqnLWwtYwama+GMukenf5aST
NDiftd5me8sK1aYM+JnIEFbXzqQFTRLzdd6kEE2FIX8owGefETXAJKBJvyRYou1nvShMPdcyvIHK
OiZAk0sLqzuGhNfmiVFMz4JHCpftJzWmVDVBh87eh8kq+VgunEh3g2jUW6AvQGuaYkmdNzIMIEAu
fIWoUwbZBYBJN0QNxDRqgJUq/1S62Y6repKXzMYlhg3HXxgUB12xO3h2w0wofF9hs8ppeAAlVQ+W
VRemgXeplwKuXaU3XF57GtjmdXF4XmUwJIRfJN0GyiRqKkVDXvyZ+wlkKRFDlY0qw0h/wcW6VPIu
ybFUIjJxtEXUkb9+NN4LoiYb6VlDeIvNeqZxaK4YJXGBVniurukWccKJpPaATk+mN+svbYJW2dSh
HPIwVBgFDIUhjKIpi48SnEgom6VB99NxpEtwqE0K1SiloDKwGNOG/thX3Nww15vi+ncOy9aDG7CA
ToOiHNmQpb9ltkZBgaBygpn3fEiyfh20pM+MzSwu3OidS7wV1IOQLQJOCRUOjmEsg9thZa4c1WEP
SRo7bfvFddV0xPlaU4x1HxgYaPGfun5vEhRvEpnmj1DCQVS6FdmHb50pYd48DHb7NsLzzA5SA/p2
MC4snUpDJrAJm4OGfArOqQXlJuC6zbeyn10UtWdKRJPLNz/PX0o476VKvAltNwws2DFYc/M8AQ0I
uKWWvoubTiHpDXZ7BVJbAWMJMNdzFzcWIg1JrYO0afqpOO4TNksz8/CP/+jOIUFd+zvuU2fSFY4x
SuRxnmzVW+I3LbN8LAHgpZSCULX4aegUnF4UZpW29j5Y8u/ky+oLHQWJJW0s5rZRLPwKyik9Mm44
znoAYRMsEJ6LR8eqc6IiHcjphaOwM7O7L+aCiuiErxfiAlyitJgVRyXg9AZflAmZbHlzcxjJPT+/
Uxwof20GU6oIDr0arsYUx6LcHJqIWH19+kLW5aLpnsI5eBte8v9PYLy7KyYnVWi7OUtGLD6cENb5
BI3YaFyhAaPOyd0Nrdu99Q9hoEN+RejcFpngacdHtzWYg6VJ6aHU+zQk6zSp5Lpbq2pZ1//FQ3Ui
duBgfx3ks4RhqcFhE5jV2cVy7kgobTMMbQrI6Ftgv+0XAntNLm5388wYTwrPhd0TpgNuqrsYjUmX
cEg6mMy7mdYLYXY0sSQSr3i34TaNp212CCGg8nVXhWiJv8KLxeshJoHUce9RriuQuCI+brtCCf8j
MFkkXOB0I6iyAlv/4R+a7lMLhMWafq1UpEhwv3QYqSuXWuQpWRsW6rqkxGp4t8FUK6DIfFrH5/OA
YvXSw04oIDTAMu/4gaeuLz6QmLzdkPx4NVaavtHcQ0toAAnMLDawJlTG6U5kA0bsrBZlqPDoX79T
TNQIgAHaTEBGervPupzP3acCZiiVu29JgWnUdbJiDCAINQURaU9BjRC+d3UUxggCQ8A5qBOtDXjz
pCF7fg+vUp3gqiObRWC6ukXa6Oauo1/55NrQrQYzYKai385L2e7xj/qQyCOeOXySJSMic4jztJmH
4QCMKVmWNGMtzoaMDjKsP0pV7vT/zfZ1YSRShabpZmhNAzkK6Wy1qohMvr0iYKNBLu2srxXlegGb
riVaWc6mLVFZ8l4UwsJSY3Uy3CJ+BdE4DgJ6FJTjwCT2oOgxMmZNNKsCIRlLRohs6zYAH4dgyCmu
1vaeuVWfCpEjps+8LT2CDHIWBcYIZDXYZR0fYTgjYZXO4cRTFjsNZXp6KMo6dkeaqK5fNWWqJQ6N
KJXzDIqpqM5g4mSEGxATmse0n0JiPKzD0UwOswg0PmXWXiF7lqUiaRN6g6sxWv9Xj7XynRQaPfxi
Ruuqzzwt0cz6kjrtryRBBnn++/9arR9mqtXAK2q6r2uo3iF+MbbEPuqRi8AOmz8D+11qWOF9eapz
bL7om79BBBY0FLRVaLBN2JnIUDbPwQVJtOudhWWJv78s9kX9RWeTN0zciILONlR2EhWg+viftgau
5vN4TVNxeFn3oyhWluPQFAZmbhfu+Hq3WHMe6vkzkCD4j5Nir2qTc6pLaDF8GLShd1Suz/jZ+ye0
DwQnMQOkdYvSYDjrmWjGCHMWHbVQFUS1ViXzIUMrgxaa1t1YhpV05G8iPsUy3Mtv42Da7Cv+oCto
BUT2bRcL4J/bEAYhOFW+i43vCNYYIzBkg3275KDai2Fc5ffpniRQMMcmUnNsEjRifCln3tXpil5K
r35Sl9F8lCjS6ATkPX+MMmE83SZXrgaNodjtALUplEP4jvSe4tkoXgl6i6Li0oUvyWklNc1dJS4y
yyiqKe6P9gNFKcy6FY13iDGUJUkVxAIusA5X0PSDTGQ0S9gwA+b8hZP6JQmU7gTavlj6/o4FeMkn
6kaNGnmBxcf9cIoEy+4Qlxtz3rmxrBK/8s13wfCdjsGgixRmlFYhMziBt44l3h9pqRZa+bgDDimj
zUHvSYW0VW017yPRjudSgDTf2TJaz9wzb17ud8Uft82yJ7JQtRtxfvjnrJ2NbUtOTDrEfT4mTMC6
So6UcUeNwgYgjcD9hw0jfaBahLO43edLhKO02+JiIxJSx3D93qaF6qM4SEFiCz1M7EGJMqcgS7pn
RHBeUPKe2Zznxwrx76daumBNbIs/5vzaHaw2E2Vea7BXqFEcOarVlf6WUCTRCmO5wVetND94VWRm
QXw8EQbiOswbTLS8HbLZUq8Zw4+pPfDbBHTBComDmc1+zHUuChlu2ki/0ntcFXXXu3i2nPJSSfmt
q7ALfm3drl2E9MXAvsO7/A1ID6XOFF0rVZR69cufzGAfWcwXWXt0GapswdR1z+9g+nZkay5pzAX5
HI/6gQyeMycQvEsZVw/BRwb/lp4vBciyddPg9GHDYI4H4j6FnuDcijuXQWk/ku0YTwUhZKDG1L3V
Jcg6Z9xrtNcLgfhPVOJTrUgEUThu1idZ8YI+VZCyU1wyMxGneYf0nQAQOAm+SuoNxKD93DWCv2NL
vhmYuxOe3Wzulb96wUpCrK89HVZO0WY1qxaQlChwnNJbqkMbeYsnKihiwOV1HI2bf+bDXKWWcYo+
syKb0jAffw8hNgUiGkQ4JNq/lmBcFyqRPvCDMM+4vnhZXsfeIDSCcb6jrtHN1lQ6VbFjARpGCSVv
CPUJT+mWkjet2Y4sRAC8V4bqjKuXdbf59pEnNDx8f6AXMyi8tn0AnGNChrUshvXPf5Lx+FF3id+4
rlFaoZnOjGgtk9YP6oLHDszWl6CQanvCupgNtPLCMtQzK+xpeBEJXKpYKKOIDDy/nnOQH6xwGM9K
yqj1o8fkL43sUn2b7pW+aBoYA68kAv4XDTc5kF7OtrAgisITOHbWeShiFB7AASD3I/zu59qbjIcp
d5XaOhI7ZTtaIg0otZ5vkMHR5hQi6QLqf6jaX1yGRJfRIhyW2AvtqNPOrDpSohqhC3tTNYOQd1wQ
jHLlumneXen1Aq585k3GBONlhOSl2usPJfOM8/2eTL8lwQtCNQ+aA3u2+ShK3vUDun7NlyraEHw9
a6v6oprPXivsOY8O1EwL2jM/AhHwr79DSQ2G1IRYNPmUNBZvY/IFRdHUoxJPNH3+uuIava56c43+
9QzQqJm7w8AkDnCNv9JciTqELX1Kvv+vb+vc520/yzeU9VNSlYgIhHZ9r2FigWkySFaSLJWE50xX
ypNdjCJj6Qjlo/LVbigRC4M3CspSALLm1ZeVwj7nQkN5d537lpxQOnrX368pVSEqvUKZdIGjqgXu
oC8CxQldzkVrwyyUyfJvbdDyuLB74j2jY9M7DPvhxVmNhyUC1UM1y22yLX64E50Elm4ps2htydNa
YO+SnsX+CPCZg6dvuG+ywJ43NcwPPKPlAjxKXdIfeauzJ0Imh3gAX90p1CyKhUUkxrp3xq0Cf9vt
rNgtfw3lnyIVatArxKZnYszaoom4UVqPtnnoCQ5oNBsAMF5xXJsMOyutWTBbTCYKW+9PZHbeIVp5
scP5Jir5nby2vyRh5ky3lt/5wWCe8r62dwKUCU9ZI//sOVRxbLizp69oSVzDWYtypVNLvWFmLdY4
qaxjTDDOiobmU8C6iBtmuKSu6ag+hFye0r95HRtIiO0mJ2XAD7wzMJDtES/9vuNb2US886tKWt2a
A/LoyYvSP7LmSGsccP3d1TT78B+mzOA6RCmLzYth/1szdVUwJI8I0I/tX++9spor/LcQaPSecJKI
pYXElyBx2EfNExfHPa63j35SApjcxwE5SLChNlo5Wrn/MbX7NuYSQUuOXDLbCJQhbbMQsj4v1VA/
jBZo39Zt4Q1oKudWrLj3dQU4d4FjN2IUW3Qcf4tqgK0FjrG27IF2AVqpLADZVQGCY0wZnC989EJi
I3fxsFjEg4uzUcdgd6UnW2XqOMYXubuMT+gqj14SXI0ZqJYgTcKICTeTuSyV+6PWjHkp+VZ2Hp99
rQwbyk6lH7ZcksfUUXvOQqbIZ6I0BvD4zjztqGoVxcyUylkmy00GyGFb5zgDksLWObF5dhblN2+H
d1yBHW6/8fs0rLxHLx/LudS7n5qKmKaKw/I+29eEd87UE1ae7OtUYfBzrKFygF5XwkNek+y5rMYG
TOYG6QUXe3LqZ+oE+ITCNs8qWzMUINkBnRXGwR579/pLGILhmCavcYrce7f33WQ5URF3tODLhdGD
99qMyckbAzxErWYUKbDoQjJgyNGQDgQkOc9dI+bKadIy0A59KZHrDfynSxNs1Z4YrsEUSoFrVu3O
H1fk3AYtAx68Y++nzP70kklRkLOy3SQjFFLjykhXoF/DF2m9baaKo1AoyL4mA7AnSmQ8jF76+MMx
gg4du3tuQNCxH+LOIXxsfzUtA/yBOwj93oTh4/9US+oiEvfjAB1+R/3vfx8E3bhT1syYzXNQCEVK
OiGtN/+ALAMzwg2j5dVpwDw0LxYuPijyPk6rDygxqG1trMGF2wx3Fj463ljKij3wwV3ht+Pn9iow
HhQ8HRChBgxk3nwm71wfNOAnAsr++FBKvjmZ9ZvFDAWfjb6fAE55rqPIUOMMhVPfYo0JU0ObiG5a
ws2Bj/13s15l7joXZw/xYZyJmA2PBiZD7GkexR2Ikc8352EMnlnGBYsrYY6ZFrKsIj7BRn5SAbwx
pCFQrr9kgAHFNq1fWwX4dR4zlG64q84X1VQO3a/upekGJGUCWy/9iZYGieilLu8JqObM7WKHrNoT
LZhXUAAosZ7MhZSHp+vRkji+OthQGzqFR79qx9VbC8TWtHNtziFZ/zZMK+iq/919PIUGACvrA+hj
MBMSdsZAZgGBrJD16fSeUIwCy32PWVXJos9a39hSKs2I6Kkm7bWiCQUZ5LoqRlLITFUZAuReoIK1
95IyDupwx7Ann1Row5eYRJpDMBj6wP0eAssOOiJspR23NaUBoYdyFTBp9DJf0Sah7GR/x8UqiVEs
eaeqP4NW1ZXN5YL7nWk2ZXCKD5gsV5aNsSol1lqAt2z15VIF5bGqUF+46Q4UjHSvdNn7pxvkm9lY
Dk+i8gMvDpuKpXfEMJNva10RsTXHJJdd6Oy7lVfJMy1vJGgjIshDH6cTVHlikweO2oAwQCjf+Ion
hwzyH+OWrVamZJnZEiY0Giq/f3XzYyZDXe6bO+7rzfxhQR2IpipNjuVXIQfFuiKmCH9G3XurQymx
oe6ViKzGxg2WDjd02eUUWwj7DxZT5Uby78kGPLzuwmLoLciIaeOcZ3q1uO3+PQW2OkRtpaHDdNpK
4O3GCn1DyACO9d9dgg5GpQFhQjcma6UXK8Ub22OCLTCXZ1Z+CAcOefynV+8HnmJ+hwRrZb/HVOjS
kML8/nQhQZd+Luu8l9tOQiM3wpwiGmFrxUdauO6TpFNT/YWqAe1YRwM1q69WsE3rjunfocDKICgg
B/4u7ZKNuXnpGvuJhDJTSYIo/gn8vviS6xoEIUA93W5h+8AHLpz0NetyNDvRzQKAIoIb3OxuyB3L
FX0EkOzcuF0gy4MQMke7G40SiXVi3idx4y0w0g88C+ftqGBh2wE7VG7hyVoSAyKDgPOD120Nfnft
KU/dEKyh0XSLSQudWtcIHRAJkZnwvVhzC6MLqtti/rP4xCTjeffbIkq2KRyFuHV/f2HoSjOFNpwX
mJlVmCx1ARjr4uoxyaarRPKn6eXj21xDsyNhAMKZQZG2HixEm6oY8j3GB8UqLQqzz1vTZOcGkRkA
8RwZ/T95aH+P3pZHNW1C7gLPS/lUY0A7HsLyAac1xWjqgj9PI8yqy2sPoQbFg3rsG7M8meBtH2yV
G2r489K3e7Dr6u/0D0gbv3Mb3C1bNODV3dM9Ua4JUXptu7t5t19V9EY7abB1QpJFLevyNRxv6NaF
kIcmggnECq7U1CWI5t/RZQzaczqwf6fpa3+tccBQQFkPKZtJWJkjWVOfAbRwZKEpDttwJMAGDRf7
aE7sW2NrRrezexJXlmYlHfrw6Ge1odu+mMpMGEfgC092SPwtXBeb2rOWRKUVc9nqbtdZVt0Nxq0v
ADijKKonNbUXcXgKd4MLxzkXWswtoVyaaa3AsNwcjDOU2l4q23eycZoOIMhl0SHdgSOCNM7Scxxq
8racq+6xTGnWVx6icBcnCV5TbZPKYaAqwwrYkKw06naCJ1r5fCix4z2uvLd4tEbPNoHNbr2M9O9j
mJ/jUUMlITS2viNJ8J1F9VqVxCymFP5FHy9VEwXkNT3uvrnjy1hAmS3qYtBvtCZ4k+KfgrQqbJ0q
uIg1gFEmttC95oZEUpYwa/CW9QTaUGh1JZPB8qcHnzW3gzH7ugzH9dAQJFt5GsBMUQrAwFKdsap6
7m7P4E74iC1IwMbxyJvebfjJSFT4r3F823likzIqPG6RyvF+wqKyj1445irSEh5rYmUev69hytqR
i7nDuzFJc+UADFny2+XBlgjjSbuATdLUuGagQZmu5dz8Qoq0enbIa7aTSrkoufrQ/Whyq9oLd/Zy
64XcZIspwl7IA4oFEalqkiBjCBT/jZpxUlZMaQN9/ZdCJv1sv5uAtrpj0kUynwFMLTdjhybrWBOF
4zzwlpYSoQsq+0tS4SSZmD4QK0VQf3ZVeXvWM2Fs3ppxCsRnbptpwoxXhcXpBkvIb23NHK/11SgC
t9J8bx8p+P4f2rNJU67Oodb13hrR8CppSRm36T8QD7IW3DBddBU1dN+yowNfj3OJvU0tU/nMsTLS
h3kBquHqUvujXhW50ukrWXH+iJJDFvpe69SNZC1MiJcZW7D8yZTIBx+QMbBBHLyMRIuPxedP2ajz
YrjlVBU6G2whYyD5mE6Kj1xrv8dTychCv9T5arF1ulHV6uz5YNolenncfWF/HbpBe3MpyTMji385
Vqy+UbgWRfA+fVr+KLHKij3EylJmB/pd37IZ/QMvo0GQtu2AyDHZkDtLPrWwMHdXIjrjY2KExq6l
Qz+hp4n4beHGOa5Ny1jfn0oBlP9gg6PTVcPARzbxKQhuz0+ExH6dUE0rHWeUZMji4joKSE+rbjDu
5w6K8GseLrmqzNfC94AZ5ao9s6WnZNk/OcZkmHkHBNdRQjWgvDzt40j+lBniJ0FYjDzN3zBJOHlW
OXdo+eM3edsTt4VEeKqgPzqkd9LAiQr5Hg6Tx4mrQY16aSSCESbfM8GlOmBZ8ltOcuZc8gv40Aen
Uk0BGQvjw3BFZapUb1dgEg60/gzMftmlhYVCyuPdW/TGhiyEJmLCrpWyPXcIEslI4NC45Sv9Sblj
9cbhV1jDUW7/ouswfb1iNr9nnZ4twkjg98OCnxnjX6V7m7MEm7xn2SYd84sJe+DQ7SQGZjZ2WIEX
kNWknad839u48n1pEtSl/WsR8SWKrs6tbmeM6P6cNUoOeDFvmKESL9NFVLfNUZRXR/lIl0M1/TGn
UkqUKRM9mnX/kgOUBnYGmp9c3onr7WDyKIIMOx/PRJ3/mS0U+q3apPjFIN2nMLURdqvt4KdcJmZr
JxBZdu02FT3WTBfpBTkksu8U+iAf4NNmlUlWLpLDtCm/Vuwl16oO6l8xPPJQK0YYwdI8tQbKksAo
nmbfzdlObSs3KWSmPV19zXnbt+9ZaZWCMw9OnkdltUgh0gldZK98MkPlRqiZNSzFVrx53ezSv3zh
Pv+43xtEvr1Em04qQgWvzDD1EhgOr5SXXy7cXfDgvAuvpzmxPY9BsnqNE3nvtgxhVu+f6rFO7lIX
RRNs17lLi1g7dI4gNMFj60ttdztMeBR/H4X9ZXwE8igMaaRhQh4/kuZlkC7Iy1Swfn8229iTO1Yv
+NuqIaSCk5/l5bOIAtyd04k0z8kKx5qKJ/Ko602uBRkg/SKrsSU4hfyIdBq5R40JtW4zmRDjhfRZ
qkoBsftr+flk6M02j0uzgA97vQVWEIDBYTlPKc81JrPCcWCeSbpu+3Ctwyhj+9DGr17+G7R4zXbC
DpV+A0nJTtLg6RgP8UGZb8wtE+z47izuNpm9nds6UhdlSF1OVQ2wGPm6MNslvFvYiu3vluvPw+2M
PkuoFhNyslKs8ae3joR1MQLuDVXxI1B00bbtqSAWiVTHTBNV70yYIT/Uf/QODbIcPSLMtGjjcGkw
PIxHeT9eAj1yofKcxAPF4degM7YIxjDOz4dOWgsXcAMBcQZ4sa7svZiG6w9ld5b5TVp+YllGSVUK
zyhLCYoGWk9c3KE+0ahO0FpClNYAspyOpZ5auE84pR2A/80jvww5x3XWkik//JXgIoKdZlR5W6aO
t0q0ERuAbJLsbW+UrPzKpO+FGmOQ82/ATyeeawqU2zfbXBvpuEa4Kv+mE5XGd59EtL88S4QW0nqf
cISOCu9CSB6TlivwGxjcP5MOaFusauZXEoxyqSW5JZUzuz+mogmA81kJEyMnUTgcmbTLzUoHPO10
cMRDC/CYub70ftzI4qi23xOJ9F+b3Oo321TPyhxeQFtSMdepJYbWybqe+Rq9kZ9QjbTjY/2eMC/S
9SViDF3INCw/gtdxb47RZDmgUG6UeXyXb7D3aFnFfVkQ36/MWR2M+dcLUaJfY8m7Q1HfI1WhDMjR
+ixO7pSNa5HcqCeXKmpzIuS0IY8wGgEv3ZvlhByL3cTHkqXaiwkNC0UE1zgRJ/3kimyV5HKKubPD
gsq4B1P/Qs3mzwHVnQrMajaYtd6Lp9WwS/vbISVl0y6SogmUoHmrtArV26iBptPhmtuObZ9aPv8m
FCP84rLEhQ+1oIw4sUc8cBnx0n1Y5MvuPRsB6u9fojSyUIy20QCjodixq6000nTGbIoW6pnARGgb
ZkGMgRSCgKxIWTw4wTU6KQy+nJqpkh2bToj3FmRkf8NF9LmDgHXclz31KojEQHv3CdP3/ScZvxXn
DjK5Nyu93Rf70TCtHwXkHmN8jKKGa1FoPseRhOJzYFwuZ2HueQ6gRYuCrtnjiBDBhFu0LxvDzCLb
L3BuDOGx9Ox5WOKCjcxlFwGTMfi8kClcrJU6eFvbD/kqMIHonhjULuVAgWZtruCMgFyEXMNIRL/H
VJ43m5AKgmoBdG1pMFzHbBrbLyX/0sbi8+7hMd6pEMNAeE5EDjgQo0bieGYKij4mQu1OCubSSh+I
EiF8QP0ieRMuvGsq8NSRCYsX1KreGrIZo/Ez9b2k5qYLK5SXbwb5cDDIX2k8+ecSFQTsFmlkCSjR
4dH7HmBomHcl4xg74gzI/vAyMoQEN81LXfkep/cTDG9TiPT04qyiZ+axxXlPRK2/n0sJXAQyO9tK
QZ8kq2mr3rsOUIlQCX6zU2jxaY/sef7shH5W4JR9I2r5WJsJhxUj7j2qKZDFZBy7/+g8XsnlY/iI
HhK0PhxVq9uujV/ByZE9QPod7Lkgr7j3dfVMAjPhL0SkfTjZhumEIzknI+vt1+t44o57IcyEAp8d
FPFGhBt42O82nry2ZHHahGy4CPCjAVuIr4mK2uok3M+sjsouS5b3kBhrWubs1r1a+kTuxDKWytsX
Q18or9928A+z1wMnZaX6TXhox7WPCEQ6N/Lg+h/XhfmdpsJWdwDpNdHUSh6K1jaNgdaS5dKiIBkd
pWBehODNX+nXVbmRTJMzAkXmF8CsTh373GHMIQKTEgbcUVxd64eazlLUwLqFyqy+8qSlJId5EKPY
V3ZIUg60rQ69/J7JS+EXVFaz3Cz3TkwB+iT0Ro7qUZXiI24dpX7zcjoXGt4+Iwconf10j8eW2GBb
vTXg8+bF2nqBCe+U4Sv67VRDUT78HB7FltCKl7s7f1mlhmPoNRb3TRWG7IDJToKo96qd5e1klLVq
HrvnRaD7ebA9seINtgquVHjun0WEGrexPLmSml22yP9wezuDxDKwfvpnUhLbeyXTF5RNgzhUmMSn
xnbMsWoBOUMi+lP/vlw3fpZYwWeTFtV7YSXpcPvEMzrb5sazfiNO0f82Z588VLPGzLFy4NRcM0T7
cJjKQc/GRKsL/OrU6p1S0mazTxtldVsmwZ6GTNaFSgY2459Th5JL4I3G8Oz1GN04d3mzZ3jhl7mb
bkaakEGzX+BcL9R6Xw6iPSpXx5bv13GoY/fWpuR+ZbZWC6OWzq0k780pID9xdk9mAnDgpGFBSxra
xsMAW3w0uoxsgV1qqYo8hbv+H8kCMwbPYOfWx8FfmvHTqYyqKmc+KHWKOi6hLGo1gVvu+HrvxmZj
BwLMGyrW3ZXQy2qYRsCKr7wt0ditg0okhpNvXAPdc5Jv87pYxP5WiNg7w8pmA9rNQATdcsRAqvx4
6hMO60IOSfk9hoK0O+wG2gk7T5lomMbe/41VRw50Sb3F8+9wx2kWJirlxboY8v/dMW3ezCuQglx3
YyqthWnTBl6wUaFZZY+bH30f4XSygcVQtmLgs2WUHYfzAkzT1wsHc882m8e87gj2CfTOGOei/SFx
v4MQn7Anx0hslSmC19vm3qiSnwPo167joBhSHjbrmUXRYSDKRAxvnnjpef+1X3mlPrzTogY6v6kB
zOi49SPKHCx+xr9w+ZDwTvFYK8Yc6d3kL/74C0kUHc0uD5owz2MEMeoSPXg5BNTZGFeeWp+0/Wf6
zuRW32EzBe+wdwWQBeIKuXxLtRYaZnvGbVxfZUnadrlcS5S1vfyv2E1OBoPTlOR7QQlEnF7CUb06
45Y9NocB4Yet2KY88Z1ZSMLTCSk7/pczyIz53r+r+/qvI7C8BsTUsV0EKnl6FfEABpX8Hqyx38Xy
8WXXSg3up6deRRm0neLspPx4nvVVwXNBR+1VDufUWY//a9D3EXmjCVPM8whs3dbuQEMVFjLZYxj7
ocf56JeeZ4y5mmIkpniWAO0nUg96H84iAGNM16MDm+/ERoNsrLwPESjVwzlatWppPrBeVLjcPZ8Z
pDtjYlNXtXZdTCQkWgrcsnHFIfrO3yM3b6Eb8GdciWw7H2mpUPJRp647MXQ5v+t1zU4dDC3zdbGW
v3/A0/scbs/qPLaBe9IXOndtVxFVwrTzFI4wiWKaxq746ZUs2GXpQUuqSQhC5b+dfdBwmfqyouJ8
CeVABgw4aHsLgZy6Ldne4+9gIf9KIz0zOtvhmODpQyxdK40RBrLlhFsm49cid1/YbQLLoehnH2E6
deIHHLVWYKJL5yk4Dp59czcwJDAe8XWnhwvclAFaKEUCdHSa7NFiyL6iX7KqPTVVfsbMPQKWcToY
iLE7cWY3saOv55cFdqfdhEA7z5/adIYjqMcv6CaB6SpFoxa7Xi2VZrY/DkEXpmfN5ELFjFrkwtJp
6oGCw49EnQyyfDxiK3ZChGOUvdFaw2jBMr92wzM2VGqYAKCOL2YCxOq1z0Rk/vFJIF/1f2Ote7j2
ZVgypA+vupa6nIVfJ7rEUbqQqxSU+q3ne9T3m0XNk3Ha7UqOzFz9+pLBp9YGstsKjlYVEaFIBoW9
301hb/nAAYww1Of4j97vOq+NfQZNGfOlwb+yIlDNmVnJ2ygPo8lcbeOLktEnjD38zyAIFwvgECNi
RhA2EzeqDDNRkIOKEK93IzhWrRQnx0JyZXa2Ny+rzys7kBzS9ytpB3kcNmZ/UE7BU3chwOM7Aw7O
L0Gfy+e13Ow6kUx5ih0sYq+kno2+fowTKqUUR8dAoCqWzbzpoE1fOBaKmqLSmHzne+ZJNF6O4Oay
R6k4Y/ZhfEwXFSXpdDBIB6YszfVg8+MxuQQTetcin/tFc/+thjApU2SeE4UKCw9BUCkTGxQMrD6o
QGLgdkluclqwMNZaBoJc0LFn/ywBS9CHbTFGe1yG0ZymlJfzIES3+1jvjZNokRn/ACMMQPGPKeLq
zISsnATOPHagIxhaeQN888Do0RaDdNBXwiuLFy8a0gCT1KylF7ELSWmkHNnLKa1GCfxvKQVLdNmH
oreacsubCYyzShePKQm2SImqBRKDWDyxRLgeTPwWfrMOaIXkYrrUvEAka7ve4SM+mj6Rmz+v+zRt
u9ajiUQNpxWFYpMw7eWEKiVESEpfLo/qUksPKdhmdC243gP7OaHeGMKmDRNd3ytAXE73vyoJttPs
KJUNYLSHDaUMcpIzL8qHzb2e45QdiBs0TOP2NzDoKLKCL7KCtibNSI/XgfSv+68lXn/9iQ0yPsTm
RD/rMQ3/545N4Dvl6WpbkINcQq28fgC3EXhYlAIOwvKQafvYz0NZSP7/2LUC5yVqoGutDTiC276x
MGh5ylWSnY9mB3IUO2kwC7iF9Qa8YoNzOplArZNbf91WCTCVGMjpgHP+Dk541SHdSlkoaONHOMbH
vonV+6ALYg4JoiQDYN7uj9s48Dtdlo2mGYY+9IQ9Z+IaaORRFyDbyn+wTQcOJFIMemmk/sEdmtAU
aPWahHjyUFAZDyvaI5zCkKAV1uLSkZc1vex5iV67bG8isGmIuwpudSgW67xkL3X+vGGEJKmQmFCA
9vrkk1uw6f9e7wFHfN+/e+fXKpl9bKW4zIUdnj9ummGbBGraLtzrj9JlcozA7gzYLAHc3Pxoj8sh
+3+gZdlvKM/Qnjx4oeWn286Nu871KJTeKjkgtE9mZQIKut7wr19E33nTKjupWWft0LS50ZUOgyJ0
n373wvAbfAN0L3TBfrqPAy/EErIAuMSfmEbm0rXxqyjoZqjTJmgemv9wQ44l921g27jKanevG8kg
ViQGMYTfoV8TGGETwNbofkcCdIbPHqx6Rea1ldMbfUQGb/QTujMaixao3xRa8+OcnV2aBV470B3x
UgBRy/A2u+9R/oEtOmWVcjbT3bwD6Eia2yjNW5aJ17MiWkwQKUaIeJNXmmCzZt2Yrx5J9pXWqOjx
n0sHMNKcTDnDjBXelJfZFgU4Y+MLjlpDWjeqEZA+HxifWdZtaxH+y0/t2kiQLxrINKJzLHzZn/rt
9sU8FEjKwgvukrjj8QwRza4qB6dWHoDcsqbrCuvd2zX1cbXp/s/3MhBltmeB1wiSe0HzLnol7vJI
TG8qvh7+PhNCTeBWqXgI8OxhHmaWok9uXvKf+D5ENqv63k5SBQ5E0C3W+WSM6F6s0enHCmws+eb2
y+I1TWt3Dz8KMwIWr9e/em/BaRlC/us+JnHx5CLbJE7uT1Kwbsqr6sp3NLNL5E6VsIU+zLdfPhaQ
/vo+3LlQBGmDggA4HVj0BM3yIUsy7fnm2fS2kKnIXzrEjdXicSUUDKvWDKDtTlCY1QbEk46SNwEj
K/9+2XIEv0Hu6gJsCWqhxFnXMwUS6uQoXPmp39g/7rqldhtiv3Mu95SCa1+56T0oS5lMUmIX/c1F
L1FAXt8XtUVGgR9hKkueX8nqKRDSobmSwZZGRHX6N2dXSqsa9DPVNtr+om7UMEh22E0N5E1m0Grm
t8dyxqla3x5lwwtitvjNVQg2w1tt1GCtEt5Di0z002dB7gm41HSEB6u6ZsoCdIXqqgv1czBPqv2L
vNimqNbIiU9oko9Y1axm/L7HsA63LoMxPAS3EkOBKNQpatiBM6NK5/gwEY2FywGR1NVq8IDwQLhP
6eBwCqfE7cWCbuJuN7f45UwTR7YWjyoJRAUGoJ9VjD2MffRedLqnQoNCZ3KnBG/WZUj6Sh20vlG3
bbDegq9xY9/Vui6HUffN0IAZG+O8mOkAs2aWkeblrjoFcTseAQn4k9irisO4vIRvqoeHKS0yEGfG
fHT79BDoK1MplOKRRc2BKRECx93viuvaBKr1t/L3zkcpcUnJ7i+BmipR08x4ypeFrfQ/uLaZOHEd
d2QazWfCjMeIyeDIQrEvFQ7HtRPwzx1+7VejT2fiG2SK8YDx0baH6MXwf+axCQTvVXCyaTajvUyY
U39EShoXerAvSrWJnuLQO/N5HBeJF58iYqYbzPwo78oqg0ACBdRbdAbtQR0IbhOBMOTdkEMNq/PA
LqLGVWABl5nwK29/HAB/5urq8bReuiLySMZL7eCBQTsLXoje6cOPQrYlvI+XwBo8/qPrUxSOXB+X
tPl4IhSgUiD69tNjtOzU8LyFkhZLoakNnYK1H5y5i+5il6jRmj0jJv9GYyI5UP03HDpnXuAB4wKT
cU6mY/O8R7nDGeJ25PMrPv4F2GsiyW23dGp+VhXOAPDJkzyY+CzBVLU3ROPXwhjMGyx3TfoFFcDZ
LajvV6fRcLWt6HNqBc75w0kso687OenYZ2CsWs8wNRslX1dAgLP+tTryoJMefOB9nq9+OzhYcuJY
BvyxSJlXmPnFUgeV+nzcqg4/V014MX9uZfW3Cw/G2HOPzTN2UHb014lb4NIl4rqfJqhFSmEmZaw9
nZcAGPYMPaKhB8WjFbk6sUdT5KarzLehbHIHP0Kv5yvULvCoWWm/mk8oje4eCcNqQB63QjblgLo5
nTf4OzkHM9He0UjyIgcysqZHe1cO8u2tHSlzuQabphPbvgPZesWWn5WFz6MF6tMmnwjqHIXjZmWF
27n0sLrnByrwYPXPCrebzCjQ7ObnoUBOvHcNVpMmeNcEXropGKI8I4O25/tsTohOUlvADef1yGlG
WG5NSCNjz69pPrVXud1AFvFqPXwEh2oiG5EpDns6+vriSIyoq9BJ5i/cfyE64f6PfMY/sbbWONoT
xwbMbWYvcgrbqGUucKaJ3R28iQd6xA/ruXpcii4PuYKt8+fwYL03/NSjTmv0deR5kNuJ5fifCIzj
DrHVTGpkrrBblj1Rxk9pLw+Q5TNywpIvjMFW6Aoi2QK8TKN/a2/K1uDzqXINLxzlx1VPrYseLxXD
C/Az/iprHXpdk3yuLdE7MW2UwdRylqQ1eATeXJ4tjtxaD+jmznhnL5ZwmLrTeQok7fXD1tAS+PJa
lzZ5trOJewbyGPGUX3vykvMUZcg2jRkZ44qBLO+EhdpSQKu5Q/DiiQUe0n6Y3TAtsG/ChxSUSG9M
QUSHWKnncf50/z9ayjd8JlnJzqatZYMxHUaDkXW2XkE9VUCHrD1OxVLDULey20Skg6dpbgpSkB3G
LrcwPKXXvA5jNW0A/y8XZgXoW4Zvud0RcWP7P8jtyZa+khIwGxftqAmxCZQWEh1JoTDUx2YlipO6
g3W5z+ev1kHxk4/YSkdEsgI6WiNizBHZqc80Oo4C4r+oThYBDu7p8zmlgUUQ4YBmIcyufvE7cZ5M
Q7I3wpb91Fb/NorXQJ0oNgB0GQuA53xOzthDv1+hpRgc8pYCNw4DJ26wNjG7T86nS4dKGwMiG+g8
hs/cH286ltocuwCo328+bP3+0d6UD4GOXjk6Jax8T3FH0Ah0Z5kTudDZxzhC67kAg/ybP2qrVUJH
WicWbwE/QLYUdN1V4E9Dtxm0gCef12tGT1SX8hfWi86C0lrV10owoj3qjIzLFCHqwav2JxMdw4xD
fbWesIGRGHlRd1LCM8yKJPLqHvGzDp2VKXMgFIuJQWF2UTr7mX7HRTFZjokau6SCdTaQChyiAHo4
vbnPbym4kbudNi1zDLGv9OXXaZ1Mz3mJc/qCURMI8c02tKUBi5mCX0LyYYBQ+ig0QfT0Bnbl6h0t
6w0wxyNAokNqzuB7/AJQQZQ2xFugPrOdREwzj2HPi7wwHmRAnGnROFifJzdZFFKpl7HuAz0bN4yS
6mFJemmYH81DWECDQ+LxCTY2pNca3WKhpoRM3wqZ4ih6/3jK01NwOEyd44VUq5ivbdKRBaB9IGG0
aB3fLsVdoWJUDJhEwPK6o7DYmZ+2mUf5JI6NIg3QubcGZ2/OJq+8qREsAmsUbHXhV6IFaMpBRRaN
0evEY+NAfnTqDBAzm7mMOII6iGG7r2ivDaQAAS5EF7UA2xk8WHxxNArLqUM67VC8XZTdxEmcSb3W
4ai9QEXkSkrnDC41Pi/hAMR3UxA+ic/PNOsGYRAbIOnbIVFIYkIWQ1AJB4i4V+q8M7BwFriVBYwe
ePODlNNkdGYNUgBnbA417UdPyUuZviPWp4daYI5SvgCOJNHEM7fNp/mab65VL049oeGAMVIFfXBd
A+WKtuHukWNUxKdYXoQatcls2iiep6XUmNALHH3lToFCNTbNNgFd6X9K1QmOYK7prbehqRL+DIsK
+ETtwsRGRDaZa4QL81gqrhjkCsz6Fhz36fvocDqooRL3+2pGZbJSmr1r9JNvYViAPhwLGC0Gvife
9S7DAYRyBTza6ytqUXPCbCqZOjKdSajMn5VL5phJOFlCY6wCTpL8E0S/Tg1nigne9G2Y+uOQfkkW
A8TJV5ZN9LLCgTnl0OjVjcib1yim7fOXdfFTisS+5EsjnlaW+C4BRxhXtOKwC4RVM2uwWk0zcCYM
TgVptXY33F3G0/R9EW/WwhcXgn13gnb+pd+Ep4nFVr5Tb/y2HyYmtqgogdqZj6y0Eo5rXY5Vsf+o
xnE4b/o77GDQtn5DHj3XFd18i2Ndl9Qt5vBTAhLuZ5+6qKWwoxU9AZlNQqbV4KxTsoDMwb+oGnah
3RuY4T6oJ8ZTrq+QckxMBlzlzn9ZhE2R7dRrkIMBvfyOfBjQjvjV/dqpSjHN+IKw7lYGOBeEObtm
npRR/JKbHcPiGWqCuywQzCTr+lifEQEFzq5I4aum0FaD23gKCvHZbFfLWCh9QkrrkYTIkw2qtJh/
HkoXfclDHSIlH0rmcuf3XQ3kpjcReDvve0H/QI/mSZdL903b5UK63+iaG04QIW1amj1UI8OzFero
pHEFDnWjj7Cfad4odP5F9MceFUmEJAXdlW70XrSXBeErB055Csnfn3nFpLTp7GixcnjIYVOzsnAJ
Cp2KJLZPhYDXSxvQ+DVar0OHmtKWbTEdOHEc3fryHRbsQnNISnDEQW7CB5f9ryZCkLqy3WZwb0s9
cQpNo2Ftfa54v0l33403/bPNj9h7UZJvs125RSoKZTW3AsDhkHUWKwKA+qNRcDhEDg0i+Fiv67p/
DQPKUt+Cc81f+Xbq7WhMwN2uQUNhbGJc4nn+vS0DGw+iHdZc7WrkT2tr/lImThDa+wt/IOzzLhyC
KoL4AILD8fyvSe4c4YrNbT1MZKSm3rCldVYQM+mt/LTNQ76ee8M7So4sQio+8misg5BWJzJhGBEM
saXbJ6t1JELoXhdDSrcp6/YQDVt8YkX6UR+3xYLqSINFc3vQN6HlTzYGsORZLTf3gEOMYjRjbwn2
93ryQ8DNmrRnYP9+yhUzLM6nBW+7S9qq6HVZJaeJ/LF2REp2O1DxQoTtHWU6ZPfEeaAxK4TaQ5RR
RBGHha66FCtweycAdI1+HSwJpDKxLaNOM2OiH/jVCdTynz28vPPXg9lJTtRa3AFUNbzAxfigTsT6
2kFnVUAC6O7a8JXYkyH//zzpcTVaJVKi7f1kQhg0sKBY+zZjy0PZmo1rDrD9cVdOvtI/seZs2EI2
uQcckYQNC3+LLqrXhP+8aa8p6clsSYd5fR7i3YyP2iOWXLgvznoLxwemxERbtn151nJyKdqecyPQ
bAG6MtLyeI4D5bysTkKvyrSA7yALHWcytvzwa6zJwUl2Lb31vxDPMN4kQJ422CVC0E0fcO/Ij7a9
SPw2KB2wUnJ48EEKp1/f/bmtHM3EzjFkW2pQYG4pcadWCt+IfuvJV6Jb4Eemc1oT3PqOCvOTLpHh
2y695njfD9n4/deD2tAVwLss3H/dKEgGCJ8fe637cbYnMgU5Lmt2DvM35LuyVBEVK60QHMLmQBTn
yTG7s9s3+CLeGURat7MDNwWcNQrhhNzf7zkgH93BzsVU6DytMal7LzVwVYzmfI0iOjXElgdoGTK1
uHpDT9uG+nMx2LXchvM5PK9D5ikbx16/YtLlJdZX78vH6aZKqcWV7Y4VfhzTbqA3vJHsqDRtyufi
uRluuSjxXRO+3l3wVZoX5AhcQEFznu9J8iTckCbBgsnBlHY1CNekiTfD3oHNA/u/BbzQfTsS8OpE
CpE+CC5BvxRV0e2CxZidEBPwectL/m57vWpIIWM/rQqNZbrzmYEksWEN8eJzQ9dVVVDc0efwPkJt
mtndIq80aY5G1wg+ZWMHYbPFKDwA4MCzksHYgtFz5O6ZwNBcihwpxbSbEvlJXLwvSI/bawE6KYSG
jOYsg71kJN24bB4OAdEeHmz/nYJbMiNIixr+Tav7Rmg++wUbiJPwOVYCVtk6gDmUfo5Ot1nqS3u/
/q17j0wZRYp31anmZB5oBFRdyS/w2xQI/zXOpfmTSiZhhzW3fZSg4of2pl8FqkmNVKkU6nP1azXH
UEy39YWzPHD+7mELsanmArVDQLvWT5uKcnMdDK4I5fvK9kgOv6X7/y6Ys66Tzr+MxhGStOe1RS6C
czJRihJgTzKI83kFKn5PlYYqarY4lsa/mpBYiH0Jxt1LMzbgn4BS/PTgCbotBZXkLZ7HihAfLA8a
TBTq7DQLapBFYb0bHPL9cyJWsIzUZehc014a4UC6vP+3+4PPRMMUch2M6YMFM8l/Z9aVuAyIi52F
kWlwbYYEGQq8+s1nYvxA8yCEF86ewxrN9/8KmC8Ej4PmmUNq1SCpH69PWXQDYkcc3rfBJINhZ2yV
VBWqy5Lt70ZOfBPlEuznqPIIWsgqTvJvAhGSwuyhzudLtQviH+ybwCrZmTRit0Rxx53B8ht2EN75
kBChwhMvdJsr2HFo99QHy+TeZ+lSDrMjP+Hzpc17LnnTc8TT0Ynz79NRjNMJtXwShIJQt1wgk/Ri
iZTEueA86n/FkkGgpGA+9cRoMEJKFxjt5XNRzeWbxTjBKy3xBoB7jJzfoH8rUTogJW37vyBw876/
xBD66eInsF2CWdKWrFwJqObwEGSUaa+dg7yJ5Ye/6buKQlPFv+p04C68X3R76Qxzy3vgBeImJ4Du
rKeJdbYk7le52+KQP71/4LWaaZKF9bJvlieVn+gfMzu6nsFBuF1+YKoj+LrsK3SlIKDuYuD5H8y1
C0ck09OOwfCOmyUx7pzgqrs5RsVF3YrwbJo9pRf/WXBqgWGy69MSwq3kXYwxYPfbaxcJFx+g9ypQ
t+LWNXlZ+7tjKOrk38kNDH31Nqb+JEOIVBFlWIM6bZ+QLAq0amo63JyVFElnCgHgW7ny4Bm8W+4X
5N9BDZSyGPN9G5ACMAhJIJ1mLo4yKHawz6swsQwhdy/rhAZJnAy47xnNS2zqu5DUyJv8ZzuMe9aC
eK5eN0bi1GlbcvxgHLYPwqoPi+iLP2+t24QezFhHVLdGmdHsE+g9Gs0svA9J4HWzAm+EjjbYw/Sg
7vSiQQ8SS1X1QmigIm3wfuby9VxZs9RvieCSDBS7FAMXYam0wSNp43HPyEP75E8c8XfTq2tnpdiv
KqQhS7zQ/NYP3DzgMhSm5eMljuUcc+aj8L34sC4Jdxd0eAGpsO+o6OXJ6cBnqMiEw4AIqeLcYFcz
VLiyEWrDkj44zhKBv+RW4gXhz9V76z9A7unwxq2Hj5RGJkRt9oIaT9U06XIgr2eUpirHhsyNk+uW
j/lU7ReQ3JfQkEsykIxlc5l5YAYkjyRlqtEj1FzvmhoEkqsKS4IG7eC/ZX10aH5itwOpqvcCEaoL
siFRgAcsDiOujbvSehlPb4vPbxJHXYwKjfL8Xg9rBKcqrdYu8WOdsraWhzuQ2ILASTvOOmZpZH5y
m8/K5RRI01Sa7OlvP6B+LxyNmVsdgM3DVsERqf9pkW1lIZCVe0dlHPLFBg86IM05sEwEKHuhgmgv
GmszKGHu+6+FUYlIg3wbuYB8QGvhoPAIP1fAuodEXGD3Tj8Qcn/jsDEQQ0aMYnrIOcpBdBNbwtXN
xU7sTyI3s2bs/LtcrDkESOEbhifRjmibF/9Yxsuyz4EY0aVCq1Alan6/StqQNTzPBZ0Nb/BSQgJ9
vOtR1rJKsKFz4Rl2/jJ9KAqMSS74ixXcUh0L0alsNgPC1hwLTcCMOskhMbOkLapNKrlRiGKFv6GJ
sHwdtwmtbbNj7TsbWfNVY+iw0kZ15i/hK6hKu19FMP68ZWBnNI2DW2tI+fDnGqzK2MaFWGpFJaWx
ck9Eg98KovAREihNsEzJ/+LjFen0jtnduMSci8pmSu/oXgUDtJqJj2niVU8TmSXq9N2eruU7m7uQ
yVdzejyBSPaJ+7kqMmxqoG7oZYo28vrJjTU84SQDB0D5iQLBKMivm5+gZc9/CVLdplmUqwfJoBVt
rPXWAMB7uaFGSq9QksIkaIXAM4NLJGQ9rKZL7kJXm7spHlkG8y9k9qn+pQ8RTf5+gc8Eb0kvGd/9
LdCQQNpfJTAn+qM39wkBD5UOfPfiSIcPMvYJX/rcCZIY60r4ZeAxk0fq+sXT50HU6Soo04NRload
NgVZz3hqtrEfJ/biHh5qxH8L7X3TjRCbQCkfU4tpLn/qVDY1mx3wUQqkccDKwCLcuBJFkRl6loSb
1wNyZNlH+L6IxrZgKfOCALUkIjYp0OH/LRXqm9G6NhbrMqQF+rhXM3AES4V4DCwjLiQvroRtMIUY
vH6cjCK+AceQUBHPUCqF5NkhhzkW33BpZzfG9qYc5oK1R1/IDjtS6ho7LHAdS/9hi4+TEucXpEku
NiCI/cOtzsFtFfJAdOjpvNIKV3Dicqd8aigpK7b/nRtfXKh3ANnAcKp3LB7ipeOZojBNuQRSQei8
G4YnzfUaR3roTIBKWqV2rjR4fTAcs0jmhoFF12DY+nICXi66/mtaNxGLKHVZCONkUZqOVGEHkIal
i4OSHR6w2JsKMht5SxuHxu9P22UuwVGFtClS99kfCOVGqULfEbhi2s+UqK+7yowk6BXgOOvLKQCw
zJRk4IMSUwRGnitQhMVvtZ/BXTUmS9euT3giWE5VNAoqRL6ybpQDcMSLfMzMpphtmC4Rl8XzcJ6y
Y440VzCtARFp5gl6tp8/Mup1GBpMZY98hzSMx3ql49gKdoQaTuLpM9M7LyPIUpJa8RpSvg9MlocH
SvwDCqoXNLrkAhaXRZMjyzNZ/8uv/xjzRBYW78B1aWhhHCBWA5pr96MWSk733+m9KK5wxPS+H6q3
xf+MVdQbvMF2eI/45d6kNf9LajiBnul5Z4KbWT3LKUZ/6BmYa99SJXsMxTLAwTs5Z7djZrGrySEE
CbnfFfboD35x3ol56OdyQLjBc9cM/n0O0JpK2FnjWaGrs1eJ8Jd4VxU0mdM573YYL8vyoCCrry5j
q1Tq4f2ht3g7xnSJWd+2sWSRHXCoqzW6wLzb19A/yPT29WL3Ezn4Z5Zpo07gGK2Jyi8yo2rhfu43
YojC+ovAdXJsw+EOPZdCyvJNyL9Zn7dGqBeUFFtzq6/s7Gh38SixOacn5dk1XjObIIEnxqk8oCCB
N7l7kVwo8GM/XVqAQAEWH1Se/9qmD13hd1RSioob+lAtR6uMj/gtG4RETjfR0e52rXFlizep0xin
q1ZFujwOV8IGaVOgOFr25R4IG8u7HbBrcnCdpUTW5X30xuZa+mPN6t2ECs7enZUk7FpOLRtI5CNG
glTlSoC8oXWnSl4Mf8YGbrIBC6sUsxKXjtS7D0Fux/ZqS5FFkvGu10oHOkXyXUjoHJw1hCQVCY9/
8pjWpsOKCwFQWG/F7WPejQtgOyuvV31oJrA7r8/PyXrbgZkS/TKV4spZoxSyYLHDFgx2dHx2aaA2
acUVXv27y21Cr+kSiliK+0DDyX4CDgrEZgZvsuTS9eZLGpbT2l7c3KmAbZyw/TI1/8OEgl7x+yrU
vJQQ3ZsujTRTezHbchTnlv269p81aQlAu7mMaBZ5MfFdkuJNy7RRE8osj6JZXW9HDdAAuowFhkdu
39icYBgBh8iowIivNbk9ebt+Ko9rNVVMpfju6TUOmfHMP8aFPFfV1vXZEVKV/9fGLto7z9DjtT5w
5ur89Zd0/XZt1WYZZRWUA+B6Qn52JACQxMl3fXzY1Hzp4uXkVL9BeUWLIRcgxhDKy1XDwsN578IC
jT7Lrp9Klc4SEZiRNKWPeVNpftFRRqYxg647hcfI6JnbW6dRVTpocpVYy5KZn/xWmM0poGkS2Wsg
fNifvrVpntz8wgvGgzC+dU8geSLgpuIAkSTS7oX6i/140843x9nFr2vmiJuHfTKlaC1qt62j3iJJ
iff8IzYkVZ/2S2OCI1nh4VnqL6SJZ6vVf4v9YyeXikmOeN+EelCf7VA0I7ookFaJRqN0VuujWCrU
egXnTy8dCx13VbPyawWSwX0HdCuNeoFJJKI62C0F2/FD2fkUpeTJR7GEwdVXK796KEdKrz7YqfJx
+1O9OsRjTAw8xTudn7LxZl6ifNRK09GhE9r5qWNUWbda0N/j+z/b4sEdMehAEmTeCxPw2bN6C5gF
/+PnyvQW63/nG5tqtfh6gzpss+0aH+dCg/7GBDT09lH8SNL0l2vrunZd6oBZRWg6RuGbS2P1lKZB
adc45f5GqGQ/PcKzsOVtUpD0kYYYZizpC2yXXR76GapfbdQSIK2IVXPtnVZtVhVRrUfnh6AcGm8K
TXEcHmLMPz/R0tYOhdCaDs7Ib+0t44damyQhIZQrRW0+Bs3zTBNAllhkzVT6BJDEvKR3mrkEpHWm
G2EjMcuQLF7mEdPJIyZxMPYWfABmAALsPxVmtfcZdLRvfViDoI+F3CQYvcCD6U+i4LvNZhwA7YUt
gIhz6+OFjDrOC7z4qBIy5DcmwjIrHwRqUt18xUMQUGitaE1iaRzeaNa9c0fz6qbcQVIAl2ra6cF0
YHKWXxScqJEgOCHgclsBmX9fDBzYeH/dOgkHgA6Z/NnS9SIdtjCjUeropw1DNT/C2zq+xHuC0HyZ
i6QXAdRahRdGAvcTuTwgKb7tlZM/dWSWjoUOJYVGpbpPsQW0IUbCDK+UoUstB4qbuNaAujJAlSoS
ULe31fLHWfEeerr/+AcwcZSZqYNa5HgwqsqOoWDb4gDhHuDazcs4ubCaUMbGzDd8GjcwPIcsxtV5
aD3E/BOdtndh9LDYjIefqNYGCQcLIOi+N80UY5RIIpMjkB+DXu8w7U40+xrFhkEhsRZvJRB7+Lvk
DBU3g1r8969N4Yn5C994j2E4SBRri/g3efA9YjCtcOZeUN7Han7ujSpG5PGJkOsbqxSEazZXWDwl
6QNpiGh6s2ucpejibWM3hNQhp3UJd1byO5D+CJQ91u9WDfmn9+kw7gWOCyIuzw3j8LMBeKDhbbcw
WRfGo58sfCpVjSQmQH2z17ZN6apVYzDHx5JjnOrV6bgt75AUnOpSr+mohLibZlzW+rHS6jr4xBF/
ku+EMoyAPP9bhjsGAPvi91SagEDTvcm9SonQ8fDZe2wc1DpCmTuSJ0NjL6xZDW+UmPAyY7Gg2eAC
9K2w5NjzUTPLJxKwY68LuT/QgclCvKM02e3LdQhSpp4OQ6fAtFxlACLdDROUtZu/ecUeBckERyi3
tWYWvbdy8zcdB0vj/xqSStuEAGjdUaa6vyv0jEeHpIQ3oFlXythKC/D3pCt/7BMYY6XJUPpfDpS1
H+w3lE6b5NAAxbO8FnqJRyJZEJYHfuK0LYAv9GaTfQ1TbJ4V7UoZzyx7UN8aPlrOFMaiEWZ+cywN
HS5UYSDbdfnwyb3o5nWsud5zqMN+o02rwYoYtimnd/cElvLlXQD32olqJoKt1/HzdLwTGlpaDKf9
Yc/KzkTD6ppoRWq5SqDRszpC/aeCqaT/hEY5pn8jR1Qj6pg1wiUKA4stk/xUDvWL4B9hRUjDDOXp
5vzcouaDB2spl9PamTBHs/nUd9ypIaOQx3TGTIX8d2Y+QWrjrX8OFd0PbxxZEljSvKlpyJgM0MFX
1NhfXD9XOVUivC78tLr24a5KLyQQrtCJTv24udi6Wr4W9GtglL4vw1OQ/SNk64V8dhfA3sG9zDR8
+HRGOZWFoQB8veSEgCHtwo3TLQNm9M4Eb9m6Yp5f7gVOZvKN15wv9/gNjJZsPT+1yxVlAc2Do7dp
ZFxxedNkLRT6mqTtGgC/dKOwfaJITTYfNtHioKUci8QXMvzE4aakebbOkcQPY5TDfwie0zXAe3wB
Tifbmp86nRQVHZSLn3AfNjcgGo64MB4wCM87pybO3LpsvAyKGFftLZSFiy4dTR5wL1QEMdSlPgFB
4ETayrxd/ii6L9D5jpAl8FuU05VzgGd+Okne1rHURJLkSaPsNi1+AMyl6OIO99ckZu4H3ZeMBLAI
xR88XMW58ddOsM76n1GZh1R7VaVnCKhYjktK7g4Rc0yNIx1YUgg6YsffQ9YEyDI71QlxP+5tdsns
5VSfPUrT/NX4Pfl4H/DJR+2nx02baHJb0SOMFXYXdbz6mNEW0eYX456EYC+qP3+k/Cw0jF+WiG+l
gAP2uz3BZtx289v056QCi4zrSosVAccYTUUC7rL9LWJCtsi90b3rsLF+VlaQ3L+ZrIjbySMAuz09
uuWo/Ipsea5oWy3WSYKtDf9E/zvDDH7eofsV8cPj2qPWDL4JnpQAxFn3CFA4WDiryZf5GX17bG4m
N5NB5BI60cqlUDHB5XOPyEJSfOIfR7SRFYrkt0RbJZn9sXNlasUOmXv4EMb2Lia0sjSjO4qFA/N2
eKxLURK9S05tePPWnc+Y2UGPtrwe0mPq7LqybMXM7FejcXvFpe1jwQd/M2ZIpYIlU+kuuBY+GVHU
VIjiwB2JG5IsUqG8kWFMRkfpxd7NxzeteAlQzTT0JUVZGf9e9oe8k9GjeqOFyrHdq2BKsPGvtA49
fu+kg7yf2I+4jmhvCat/nLHt1lkj9G7Pn8WRxvVG6w5SG/vfJmwxH/BzH0VIQNYdMLW8U+0aqVRG
YzZOSnBVv7e+HmUeNTJ5nNDmGg8SxxYqKZR2WXkPqaUNNRl1OGELAHwtHvdBXLhc4S8zzdB+wOY1
FKXySQElsJ3jkqiA/h14k1FVDs7mPqfum+I+dc68J6Sl+P1Ni0KK8F21zn4RBLywxZLEFZxzSSeF
zLoeIgqFITRpBdL84yTJEXm7Xv4mHSRRK06syUmTEXFo4I0khO1+SWMzTEUxT2KaqR+HANYGx+Ox
rTw2kQFpL+Emq9pfYnv6EVIxIjy+oIx0edUM6Hd+YaIW5ZyIaO0XVuPhjlJuaVU4N9/LSH4qCaUP
G5OJmbtrlUDSUAKBxOMYeyedY0N92CMuOv/SZ/eY6X0qFfsQdYUNkWNapitTqN3d7zGYvfijlnmq
w/Sw/ARZg/qAM6BrpeDKWXMhxF4CQuEu3jM+R03epEXxp3WL1C3LTzso2xbRopBZ2Pa6C5wQotqM
3YG7obOtV7u8fLyVMLj9jQFp64UsPECQkk3q4nK6UqvqKqW7+zXzFhHNqGXIRbuAtwEO3pKeuJ65
e8q4AwE9NpMg+uzWKlDhgniOlDS4WBiOguyc3rFxKWNTxgWWlOINHjJ44vaAEZdQly7CA3xkBt1o
PCg2ORS50qcVU25MCAJVnlBIifOrbRQOgPRxeJlK4XUU7L3ss3TbVwCfdaA3YE9/BgKxsUXK0YUm
WknUgXynw+QQXnwIzXQ2H/hUQB+CBp/TaDZPO0O5dD8SBqRsag0ABFMs8bbIjkJ2hOgqr9rLWzYW
RwDfmYFkzwmZcVgcQA8Aki2NxD7zCXCuLfJuW+DViS8Vo9BuvRksiBQt7Io+s/9vIC8HDMSDzFaL
qagg2v00ZaiF/obtW+8FNKTzRlJpTbvbrDr0R8ExQ4sqnB+270w2tnkUdNF7dY0TAx4QcZAouLMz
fyPvBv2Jii0n8bhYdUABieaY8R+Oi7m9YkQccVQ0wq6gj2E+/VMI7JnAxAbSVjv6PkphmYQqLzKE
IegEv99bpm+DslhKyjoUOYxrKm2JdoItk6GpueA8JjkvljDEVZK6Ddsnr3FgJe17NpFICD+gS9aS
fnaw58tFvggafo0kZyla4uQ2G8DA42nVjzJnaXAwj3yhOEQ4gEHWHIGfWeaF7gAYEkZDlUbsZvis
bBA2GF0dHtnUv4vJXLTFwLfGxb7sN6GoyZqfgF+iue2f+Rb4d+EGIdozfKAvMBU+eaa/p/ojOjk2
Yl3pVo3TBBJH/KbTNaQj05KjyFTS3jpO6ta4xsxuCMEgfPEjr8ROicd/ZA4YnycFAIRHmmD0nhD/
pk97jmdImjK7AYmwFqwSmPiyefC87Tka33tsdQ3gc/OQEDs0Thx9fT+tOMVFGnJZcX8Sp1cobk5h
u8kagA+zi/8JEgIP8V/Y1AMzjagpFCzBl9BftsnNPySK7+o84Pps52RY2udGIZOeSS1z4xEWhP2A
U9NYDs2if+zoigCHv91r+LQiwUQO5veJKbjX42vmzkvlw/Lxut4uAFpJunUGE87ufFMuri5EkWoU
x5E7pv/ohzGJc+nwZMkm5xXYX4BH8CXcfG2vvWmvtF0jJ1dlEHD2YH/eIH4uBBJixMe+tunEoQhU
wiMY0zDsqb4R1qa7mmIDpIzRLNeRwkdrTsclXfRacGp0ZoosjX2RcXBNXmxtgo8JDhgEM1Ksz/ZM
J29NEogr08dZMpLAFgGeuN/7+Uol8X2EHiBrbS4tJH0DZhUJPzV5FTYqWYeG9wp0fYbN6e2PvinZ
l9XZBhIb3XXnwSiy6PjREKsI8Nm7Le/06pHhRL7Eb1Sg+uXLNNwRqsq2foq3LPGmEaF9FCpKyGQD
n3exSJAevcuZaVOtxNoCMkH5Ix98DRrXCsHU69kqshaNRz+vk/w5sV2JcgbX2yWD11E/zFVPh2WY
26wgqVaNYoxN+bmioVdjGSG64zs6c1/9bcWwnDaWKHP97ybLtwHo/jhNWD2vyXZylMwzQE14t1L7
IX5dSp1sKra3pRfr38pcmplJQ3bKjyJnhBQk8cP8N+wlaVpO8+O3fTHHfXcBtaCWUsQtNjvQsLe6
WxvVmf364jKcUkyJEex34gMvFUw/PcJFYLK+q2VTXPJUGOXGDzqg/j1MHIW6oh/dBK61rjvT8SRt
iW79clmM2VG6j/UQh2ZhLq6xrKQevhxSOak3d1m6g/GZKxriFLX3IrP0L8ajjRulrg8YiudpFMpj
9uH72SwT6AYLiL3oK1zF/8VjCBQOislQygj3bdvKopcYsNDxRdMTaLhJUKl8gkv1ybQAFW6jCEiI
BY+mytB0R8RDhoNf4b7lxo/XvXdNl17tfQ2+zmUZfNHlc7fLce2gdXMghZb5kKy02SHJ6L1i9pZa
tA7JLRffdJn9kyJxPqG95/CYWgokwcn+jIwk9gkSTNDZ8FYiKYHPL7hjycCs5lVB8qxq+mNEzHUA
kAU8J4bYMHmFnk5JZZAiIWTjXjN2qb3q3bU9u5h9maDH4VQxvQWHlxCap23uxRcoSaQfvOwJQaba
yJFinbZSIfdFrrIgeFaQGBwGHP9K7nzpXy/Gfbt5du7X1c0nafTiMANJ7yb/hr6XZ4RaLxP7jLX7
tIWy7uPL5Chy1u51ELTe4V5rQxsRuiU9W6vB6+wOJgsrAO6CTR4eTwQlFY/iHV2EJStip5wEYy9f
yI1C5I1iYiXQmpRHgVofh+RjE2cONmbwHhTNXQPXnt9wlwCpQGl6WbteRn40b3z1eBGv8SxbPVMO
3PpkuA6eRqC28j0DBmxP2aMKHrQ37E70tICzWLfpBpUVjftJjSSPZQI/AvO0lwPWGrQUnqqBsL9c
w9RNpg06mztFrCAELncIpQZQhv2IEOUq4qdxJimmA9cbrVE0EhkS+q1a7IdqIfaJqjPLkK3Ru16U
1NCXcKUjS1PIp6ZgdTIe38FF+e4DulVyhtSAuLo3t62ajolirbvGmtRwAndX9DBqV55bq0FrWJA7
J2yp35YvCKJB/oOWS2DLLDNnLnNPiH7qCWzRdjJ5hDWilNjDgO5CoP/Da8M54kGMoaOiiUzFA7F+
YEYazHBP8HE/mvecJCITazoOi1r36GWZl2l4aznPNTeUiyj6y1tuSVES3TWdDyvKBPiRq0jmsgLc
8oKtRg4VXJiosigVhbaBekqyrUJUtFFz8FARBlQyVxXytDZCRqcOw1uZp8KfqClDG3y18l7HVa2m
FGnHtsufcmhn814A5SfK8aNfm+/8qGILALvmiuCuuXM1CqiVY/x9d8e9fb8mcxQthyyqzt/IIfZg
/VWKlu+EibUd1nZXMJPxGgKBiUyXkvsi61ZulkNeElR7l5TufUo+dgZxGGVqJRyOqNvr1NEp+hiH
MvxOTG/48tcp31ECgYgoTRslfoI07UGoV0Qg22AbWLE8E8ajTaM0NL/71wMBE8/5BTvW+WCwmL9s
JrtzdylRuHbgBjnKZ6RYdIfPXlGdc7uzolrsdtRXm4VONZWLD+0t5mUHBsBZUNbWfq+25ZFRjdEH
MzIGO29QukmW5WiAF3fKC4OEKxdJGs/ag3V5/b2dF2Mrz28hY4MzIjogcFlo10bTFb6v97BrFMO8
SXK0F2mzSwJUO0Xu1lwbclXL64Rolg6tqrhILgRuAHqDbuo10rPvLQ/lL+gA7nfOH8eD26pI1zVN
pwdn+xbIqUiravbsw3OFzakW6RLHPWZi7aw5nNdtxYxjQ+s3QwOXOkBCjdFZU+fR9WHjn1PiqqIq
zXG31ThQelL64zKxNoiD+k7+lCZ++5Df/J1bBTBc0Mcr+c1alBFIH2r/uDtLgLQOk8KsIl7anGl6
6tjeW2ZsHQ0kTH8+VqWvL0p1dGxkBgoB37w/jdUMj6EVy/YUUbqpwOhHgKMbf/Vr91xm+2Jg5bcH
b2lBfj+Um6EHjHliVTUkolRRs6teBFbNG6XNdpwgqYV0SW+pzx3FjLwe1ZI5gGXMsYvhuHhAaZug
00I7NlOvQB5SaobmXdqWgVB6u/KxY18QrxifQxDSXNWFNdEWVAewJJ/b2ma8oWnRVodKWGJptGa/
imuz/ubaIFIwXoXgULM5BUVtly8ZXI7Q1DUFO0GiziUrvS5wtrCGeCuiW/DH96V4FW6xsMKGIZqO
Y1YaYEE3Vn2vUIafUOKBkZkyO3ybHNYY+7/+yVEhkvJ1HG9HorlQ2aadRchrdbKUaxfjlnQEofOO
IAh0Rn8Cl7pSRucHorCkeNQGLMUO0ux5KJoWCdDwcZgBkirz5/vfp1pGHuqJxA6baQ817OmEvxBH
srcBN6d1WPP464JSBrE57L/b+pQykmmCG7l8EDqcaD8SZc0kQCqk50c9AeG05dLCXvfTEFkkAxzM
42xIKZ8FLJjSSQ+xhXrCebpx4WKKjrTxEOQJApxBsr9kfVk5UD3LVqp2VViqJyVGH6tjMDEXhYzF
WFAs9iyqszEpaZgiBAy/7kkC4NnZ8vauJjc6Wa4d0pqN83fbg7CQFF0Rn3WxiIluzkI/Fh3aEhfW
Ngbh50fdYsvrM0cCNvGLCZ7PpTZkm+LCG9xkPvpy+VuppUZxiyaqWy6DVCtFldyf3sFBAcjS3UTu
RAEarQu2KfN3u3KBEI8bRupRg7urDLAfrpJhWwADyEbZKGtvVFDxzIK8Orqlsn4AS/IFE+OtSHZs
OnFTfeeCDKY+UQm9/6yprQikrjoB+dOWNdhcpRchQ80rYeeS3am4YUrqB1wxH+KsYtl/Bk1nxZdC
gCNSkJCC22IlKW3eGe59r1KPo0B32vxBejufrbFaXAfTbW8rfAjUW7r1IKslFcrXnMw4mutYVD3N
mkEtmeM1WiVd6rNm3aL9SZUnos3Y9DJ90/3vPOWGP9qO1aBrppsQMofdjHrWKv1E81jN32zoAiTQ
3I43w95CRUeECQOwNAJlondlmpDChrs+LUcfKWRqMrQUmTABCJQTovdKAd5hfc1KYkrNTxSJNb58
b05PSWO5Wv7gYRIMG1nRqCZWG+Y/dmbjsLnLhew4mFq03t5x4/6AGMly+TU9hmkR2UxXavgNtpbV
8KbXbqNxWC17AxJchkxZXR+MiuLcrtIL18StdLGHp/p5hN677tFyzG1f6qPpsdc5Eci7rp2C50JX
DxFW3CM4GZR3H/8Gg1ckDwnQwDjnge4bMSvwwpp/MbfYDK6RnqKulY148xCFT+x0rHufYNONyOR6
S4Mp52hSxJ4kO68tHKvmHLvemsdvSVD6cVzyT+IMTzoRIPUge0nYb7hKd/Ayq98Lqj0fyK4USvSI
vXw9qWe2b/uyqfRnFL9eDMJoSw0pYcxMdj8UzZEbQY+STDLKFt6hmNzmttidv4PEEhFum/bisQL8
8LNFcpvxaerze8NlUfnSt96s7XtD6EqB8NUfBILIez+25tl+qRKU82aM/733WFfPyv8W/5JprS88
8XMj6S0W5oB4LZQmWwnBH3JeSnXGXr1LOr9/fxMieGIHblxHyW/bDP691VM5s0RGpMmlBgvERiKE
Xkuh2sRzsvGnXl/LurFARLd8VIW4BFrXCuSH0TvLovuC3bWXdiGKjmmrZf9gtjnJToe/Wt1FrkTL
dvh7Y/etAwGhVhqnN99XkShAmucb5/9NflbtFAB0INeNw/EoCc1W0GAzHvFKR8dhY9/fl/4SWkvJ
zrV0orSdvLqWsyyaq/xBrab4X1jrvs7ZsUXzPulUDk3+DakPMnLytiYvckqLyBz4GK/imgZVhAGF
TslSXCDVuDU2dVK3AsCGKK/dxKNvFIphX6AWLAfzi2D+pFLlPd4u9n5lf/pHtlcSmJWj43osboe2
sCsaEbF+haJ+8HIQiETjMR3RTDp3GZywKbJWb4pLjeSyqNwlCYXy1TuXAQ5U2l19kt4FG4PlSN93
1WRJhekttHHb69UQ9RLf3pFWqBflx5vjh9E6fUsEINWjqHpcuHO1vx+4plCUBoqgjSwtnAecFLeh
2zr7T5bmMn20QscgWhKmV90N5R6g/eEnV+gC9G1xUQF1KgQ/oNimKJNP3IaXBnD2Nh+AiTI+vloC
c3KFn/TZ0kCAhiyxKhK8nx1XAgBtw27nBftlR2jwlLUB6VGxk3E80Xe3WclsAFbif0prG1cgakaU
W4aD8ifj1J1UvQwZUN4DyhjcgtFWCTrR0EzY8KMDuqeXNeHTm6Sc8ND7GlzDICzT+UFTY8PUq/z8
G7Conq7PyuzCZydc/t/OB7j3GT25En7CdhDFT2Fmpfbd6DZvP/lTSXYDXeWEJqkGEtPkSOiaLmjE
r6CdOJjo+Tqc3FBez8ArYQ0RzCDT28shkcxo4kf0ziede7Q74QM//Fxm3ygCdtjo90XcFzI10jp8
jZ9M8h9gyk7OJiFm5VmWBqMSnKWnfhd57tkDJFqHbRC4cFXRfvw8BS/3VKfSKTblVUfHa9Kt9sly
eozFRzXny2esoEW9sGJV4ubPhQSSpeQEC5rrBuhzWZE7CHgguxlVVnZXC47bzFtoTjaB9qWF4lwm
JuwP/johOBXpWAqLiQa+rKD+gfPzB4UJe3g9oo7jvGTr74RSM8rK4RbqcLUOH3UAtOOaSC8twEX6
9m0UMUaMe5KuPPg/h4StPUqjrCwktFF0zvQsbGYWyovz5kY0qiaj1X95PIElhNDi2gMNRzTyv8i5
PpfqSdioQy5Qndr/LX4QGRUtiPWtt4+JXt0ohMm1twsPQrmGK3//JMOh/miaQREJy+iyXFRwEFhE
ooUofGTVlKQZ/EyJUYJ84PhChWWbP0A9fMJtlYCi0UF6PDimAjGxehi70TYfuFbOLBkbsoHegV5N
aZvzp42dmzn088KdC8qusCi3qbXbSOdnldi4KoByA5e8Wi0L/g9U2NPKTuvu8g0RiFRNFw+FZQP7
+jdJAwDdptrL8h+uif04DY5eXXF5oxAs3Zeo4yN5ahNxvka+NsPjvVkMFRozbILl4uadezXK4LSZ
sxaYDh6uDIqdEOg6JO7f4Me1HEeV3OlHtCzsQhWnKnDisQOYKPc7mD1P8Ha9e/Wf+S2cqxyL43tg
KAmgvivq3AXeotMd5sqGSyh2Be+KPQcebLd1Z+hoYadEWm2SxEuAUhVMKZnEhOhBcB0a7lvTgAB6
vrEoj6zFAlwBTpKzUd3QuTOqMZ/FpOSxilZhFIKY+dsc2zfqcygN6pHHfp6SoMCYJRQ6B0BVCmDK
EbgufYiT1vz0k2Mz6YLHEq+wYYUa1hpL5tD89JvO2aDGeIHnh0sUBE73S8m/2RhNVPftkv1Rnxvd
4MWHzv4pne/5BAbONocwCFOK9i547MFTalTePyfX9heDTk/NcdFejLT5UKVVROPUX0Hi2kLLCqvg
6jEZSK9ZVkLGktVu4YnZQjcCWX99oSHIkU4gL5txF9XSgyl4HKBR5Am4WgLPgEoKxfMJxw1LwQ6+
OPeSrEHvL8BTA5UfkFz6x2t2PU1kHv1aAYPZwIC1tC7zV2wF2ZPElFRkVwJvn1m6N9Gif916Ia9Y
93IXL78sXfN0wPw6Mr+s6Eowts82MVJ4l1LbNCtcOc3mE2k5q23h9qGBX72Q3vcLcJK1caDRCtTQ
/fGjoGvaXVDqIgnlgk+Diq3EjfzRt28UWBAQ5ILW/xMnJJ+cxeLAT0bFdIrx81E4XVNJkZwyqfae
7uXKpHa9Ejnl/PWPLRDZN+VgKzEX4KqYMii+pvVo0r21jDw/fn6ng4+eL7szv86sevlqxXWUQSal
3Mf8igxJeeOtSHS34E2XfHzw1umpKn5ACJiIQ369B1yvF5uTzbScrdWID9rJLlqbtKJIJ+YFzqDJ
yW3PdAcJycOmpAmAl4MXZ5hG0fRbTul6WvsM2/UE+zx18BennMDmHaYAYvvV/G/LrlI+HGdq/7LD
zFdSX+wP7iRiw5ljNks4h6TF3BUkLdpvYYg0KfpnBDmDlazXI7GDjFXCx4CUwebz2LecypHdYkR8
BpMl0MPySSCtKRjYR2krIMdaiQcSDWB3B6ukbKY45FKrgiz3kMX0dw6HmnLKZx+FNIQw/lswHbul
7/OOljdK85B+He9Ld0rcSnQfX/e0x/+Ih8kxLRnlS+kqOTRTcywAQbPRpj6xVuKWd26oyxl6Tov9
TNHRxl/AaUg4HfofJUHPCBemOPNtempXpmqnakt4O8R2e4AfB6FjmPIjr53CcMAZB7EX3zbODlNI
8/xft86U40Dx8fYHLLSKLZ/QIGjWDYksTiarKeSV47NLLk0Rg/svWP97+Hh95vgsiDkj6G6rlajl
+5cqyAokL/8dWdyBrJOVdnQw3JLTOd3mDdPgX6L3OTNLyhuNa5jPT8YRbZGqTM415tGbQzX3xT2k
zujP+oFIfqYGYv2E1Qbmt9dOQtzwKsOeCTJYOHru0t4G+GW/r9l+c3tZ2eAYTkMo2PSsKQ3BIKMh
+1rhGcAS41nuOElPUNdv0VkIZ6XFp7jQBpdy4CD2qA5nJ3pmIzkwruRt3bLhcEfdSztzuuHi3FKF
/KT1OXCo7jdCSYEdEqJSD2ejh+qedxas3LNvuafY/4X9po+FqSmQ2gZZMEiu1/rWldvk06jaINCt
LOL43Uhf/C9dV4I2XEreg0QIia5oNiofjNlWZi600qw6F0zBebWph+qITtwtfa5CU60PJ4zY4HZV
frMk7L83+V06Koq/sUD/T0TeHPlkBAYVyv2w385Vd89OKExQDP8oZeWwYoaX8xiB2R29zlpXBHCV
B6vB6QEuucfXd+fe5ok2IV3/eR0IhR2sikZYGmPw90R5LniAymAS+AuxK5CMpbTjYbr3aDaHOEfJ
egeMrt7rMiLnrZubJOIDMXbXKCszb3vB1S1hw1Dn2jKyV/s6JLvnpsJaVigd9yZsyOc2GbK/vc8Z
PZ9hcGLkT35lgS2n6ZXJiHm8YP4rpPBV0HsqkhtgCMwjlcua6i5nhrb/UjToZBGhzrSL/j+A3HLL
tRmIiCDQGmqyA+rFVcbf/6rMxTlAd2oex8surwDajHqoa5fH7yVdf32iAoO7T0uVf/kb+L6kv7Gz
CPe8YxczgPkrBPcDw7IyK0lSOd01wUvMy8sUjlZ4iB3kjnCDlala+Ivft4UmSRzMwwFBIsrs3R25
Rlgj7XV2HA9uFGxXNj7uU1OGCkQ31HV7GepYQhPzFsZ7x7X9oS2ihbQ3hhXgOuGuxLFcCMld6Whj
3Qjsv0dwrTtNmq+Qhz3+0yi96ZGvNDJEI4AQNf6lkFDEI6ZmQYrmBv/bDlBWe8sbzf/6QfNGJaPc
CBZTm9mtFMcwSdnuIhDYjhoI0ECWm08iz+dpGILutIZ71Ua23oKsLYKbD/sSyFUcRPtx1UY8zxop
rWYhv6meunIbBbZXTxV9ysxJ1vKlvNa+/fPKRrgQoF4XhbckHgxrbjXUnVlIbtN+NCrEEAWpuE6t
ITeHdF+Kyc/hmSujWkmkFHY9ZRI9mS0TjIfMgtTqRQW3yXqcEs5bINLlH1eI8LVDWe9kc1ycS8Zq
PyDQMNSsOL9wNJkDTqUQKuxmFgmmJIrL+F5PpKjq5Paf/R5Ak0jWYVwz9ot954+EPAoABd1cUNYl
ug/2DJwVAJ3BdgUuq7q/GAH7hO+V3VDXgpPEAPCg/F3K6CkNB8gLpcu2ExIvMCfU8JjWnBh7+u3j
do/BW4YI2lpj/4fzWt+jAEwD4QVUk9/C2vrtB3h/tjcBFzSVa+0GS+zck/kiBlvSFoHinwoq2+si
o5h4esfrc1/pw/TbT3W4Us19td8jSivCbe7h023c2iG4eR6QC3j0JvXdvoJvhxxy6z4GaW08fHFi
Lzn1mmf3zShwK6B3p1LdUnrQNoxvZXXtjktguGb0GAAXWeUT7+9ekCtyseMdp3F9UeLOudZUCCAz
mbUNWqGvmp1NsoVtOyaT2mxlys7LtuMMaMunga4rrFkQgcwgq3Q12HfQ1vl20mUDavrCcRTuf05v
x95z5e88APELv8x15gGU/vCbA7RYbCsMM/uaepP8+FjHPc/SuQOkOdtr9BrSJjEtn0xncgyR7eSK
+9+Hf0NzhNEchreVyizIPvSbJetruRx/H/0SMymccffJuY3FrYJmdRSDEsSS98y6LnurMX6oDYRy
v4ashO7bK/H2IZAvlWz5WJXKJtoEjO2xYqG6/h3ijm4056MZb47ZgxhBH8sEQjErfMq3d1tt+x1z
ZRd387saMWlJETUlzbdHAXLop4+5uV0npgMM8/rY6mFqDXhJx0ErqDIrJoDTyeThZrCrx1jFdPlx
p6BLjRtaUGQ4QX9gqh9q3i47wviLswHK0wDGzlW7Vst6dNn+EVbCpUHArQwN0lD/fDMJ2jEwFXXf
ORlamPL6Latizu13ZcPTRMZwsNQayBNY4ZwGIP2gnRsRnoEzM2Tc2Mv5ZGaehc3m00ASOTI+3/P+
4f0xuMP7UDctXwwzdwvTVCmk+74wYoYfQX8ToMXscABWz0yPkbHRNEzZilLNB0ekiOlttoTbIAs3
1LZ/CRRY2JB9+pSieGWXlF2qMq3rNoT8lMeFoEyfQGrvuMDA7dQdZ0nicK4lXTOWCIFdUyDNQTsu
iXlldgNkAIrAmfXXKwy+BS3ui2wqPZXORyBrC6TgRSzrH0DJ4e7MIPBdwbkKoGaQN4mua+ID8+s6
eDb3ipDxOqfiG/4CCk2LhcVBvEcfsX1JQjMxiAqlwdYOrWxbRu0c9C/ABknGSYJJ1KLMO32GG9VP
acxaSB5fIMHNDe+oTUOYXOcCK709K4KNwSHx4Zz06Vy+e1OP9EQvIMoAC4rgzdoavAaWPE48oDUS
I++9BRB3ydCohd391CDn3HnXAhsSDvY5lZrqySPeCqcQx1eqxQiJcZbOIqfWoHk4DI+uL3MPnwTJ
qj+eGvvJoXcXqWc0dIK8ZLEpALFxHOL7wuSnAdy8/IlAI3fGl39PJRuHPeiKkLwfjsH6sdVlW7Re
lI7NqXeQGHEPz2sjis6eMv7bFZibK/Oocj2AV5KYTlFoaEfp+dYlsQr+ZPSuf+1WuG3TaqkKGc9D
/9qVSn1w+dgCpXKS2++71G7/MfAuaPYPLFTzr6Xnd12FPY2NWbGQBc6WDiBygYIxA/TMPRRK8wAS
NhzbCfIpyAtv1HFe+eyxO//VwJ2LVtDMlEWyKLpEjmnse5fDQmd1icuGUZYJZd+VJ3UfUgYvlWml
qkKcV/Jbk2vTkFo2+gOVM7+YzAfLMX2anQZ7rJC8pp0o/QlRMNtDL/61B3PHf8In36SeB09lXqKt
t+xBRL65ll4dvuYw+thxncU9UAh5mWCihzlzuII+pfmU+5piIDXDA9TF+WXyZTeSrYCyKI5uhI10
PDnmuMH+cUpPXEiZ2Jt3xfaggL5llY+I7DeDe1FedqRCID8wQLVq8dAUSDCp+fU6ZOYOkLDu3cHb
t8qCCycqgQJxD8jb7h96SZW5fB8ZOemX8J9wTn/9WGNnuZcESvIRgMBdFWUg2o7aUZEAzsL2viYp
/mbupxa6Oq3tfxnntZPdPcKYr7D1FEYs2UkZK7flajeqRs+55GA3eGK4etV1F910LRpZMhcp5x7Y
bbV881X3OdDi3LTnXonw2FkpG/AElKCW50aqSl4IlHbkrWrKhI59CDme3TxlGgrKOAn07wpMO0Uh
/pVKD6hdgUdZjc0WJocRxwkKi6LnJ/MIBOm5++4JZwbYCvvFWPzH9ZMvRRg0wPMoJElBZo1HL1Lx
4X2IgWsCE2+6VKhevo0SB7YGtMt5jngk2S1zbg//9x6FjiiD+eZtcA+8pBnSQmEj/ckUAU+mPa2/
6ee1NUNi8NJ2OD7nB9m15wPyuYpeiPwKo8Pfv/bmK+O6pgi9+W29CoUvRGobUQGLrr+EcYGUh7we
2i7klpPHOiE1yZYvuIHNyZcbrffgukSg9Wp/ZDTQ/R+Beu/eoopdpE7DgNhinf91pumdiA5nJFpV
X8ZuDtK9lcR0yQv1xuYLfVLqhsmbLoXAHGbIhdrjsbHMXMQHtuMb2XGSqdBt7yV9iV0FlLbNSzlL
caqdXsdBDr9s6+ElSmuToqtGeaG89/xOIHtXAavq5fPPt2ZkC/92kSmxMeXlBuMHPHAQLGMzAmej
J+wzauftBSKCBIBtAhqI9tH0WgYn8ZbCwHPh0//bGKrr7lkJegNg4fpnV/RvGPgJJxQB8W/zuW8W
hDDG+TJcvYCu5h300maQffFIZEQW/alyMymqo3f2UdFuOFKGSNMBU99twsaX3q/YukedEsnSCU+w
34lKvkv0NUe9vr0ypE6bMJZ+dMU2T56DdHSn+aA+h5qu3ewpSn+7RQugCAwCYK6p2noznFoauH4m
892qrE5Z3MhYgmXTjudWJA2Jocnb2VcToifZFv4+fh4hNdTQ95sk5BIVABL5Wj1OOY1QLmNu+JD+
vNNA3wzfqeYFe/6/vDYTGdXhwwELTtFJMY0wKqemsDljkNCRliPvBNp9B6WJyREVP1qcKQCP/evh
Dor3+oufOHmZOah6iL5ekOzz+Gd/tTxbfMZ3Z6CRXo2/RXkCg2WH8yYOa5BovLW/VtVrXdmPeV4q
CrF98UAvRkGIPwdk9TyKGyEvUav6Yw/ag7JV3808pgsR9+RwH7bLJcXupYD461RNdik/p00WzIYw
cL8u56Y6p4Nal5vnB7zwQ589KuiD4TN68OqLO2OJnXameSAni/F/joIZhOz8m5Meur866TEhIHkx
dTALRyjXvtGRdpZDzyGsNFzZ8K7XTnPRoH1v4FQDqYg44nVeCnl54WesAXz1JYg3oV57Wyt/fssu
grdbi07QcocEqQ7iOOdnzPx43o0WspzC6mhJeYK4E5xfjEymqbWoO2BUFZ2PQWBEeLLGNkQcyFU8
X0PubY4CM9wG4sWcz3Z/uJQljyhbJKsuv87NJBHlW3sC9gDm6XXeIFXXs/M6KjrC5Zh7lFhRKCO2
o4Q3WpFx6FhrZetO6X/bQvY1umFT1nInjpRVS0wnUcPMJOYUbypZAvHL0+m7dKvSIJe0+xwxYCHc
9cWahsWzKgi+JPExPt4hmWQRfbapZ5EAU+j1Zim65HW5NT8/ZUoyGcBWvZGr/cA3wTbZoIqAC4xa
OjMTmkC9iOiAPe0k/tE2LkFiYn8wAnQSoKplmwixCkODHvEb0td4pPP5hUvxCgZy3YysHYHTIJm4
51qo4uaROot5rQ8F00eIboJ6moHp7xF+ojpyrmJg4hckGRmC4f6Y94HGo7e19FGaXmgFtCOLkmWB
iAfLjAPYURcyqzjkG+9JSJ//PDe23Z+yEJb2nt93ABf97f5LiHyDtjaYHBUS0n3RdhSKd4IQhB4f
ZW5umK0xqSlAlG5D7ABuC++eL9wCHvtEmk6D4Xcfw9drp3bigThC1ut66JCo8Z9nEvSAyzEttEYY
ODj7EbxSTSjWqfr5DKFzrL+6Zr9g+cb8+cCmyInwvzMOhCKAkFe8bR2LyH6fFhF6ZiRYz4Vumsr/
Kl0r7xanCyzIuc0COPvJKwjn8mekkQvz3DJn1Q42nY80aYuz8KbfPOU6xM0oEsgkMElAUnNTjzaM
hh/AlT0TWgqDPYN7QjAJBe99Oc0l1OqKc8F90NbIKetfKbqR+qAN1Pj22Sym8x46qhwC3Hd1e1Kb
PPAaC/P4ubnFypigrHM15kkzixzHBEV4krLSwMXd6SmvlCoVmp7weKi1gJfPSf/XS67/Oyck6GcY
6NN+IcgjxcoVg4hOgM4/zN14aNNLSGv9GK9PXTjBeGZALU+JVkpSmXbAq0vhrJw1foBRVdv2ABmg
Fvk1tg/hUfvGNEDZ45BB9yajtyfRu/vAKHdK2N++XVh+8p2YEiYQAJRDKx7E9kQlpnVVJ2nKCVWl
sO6U5oXObokJCqDwrTotvkO/gaMuIq0gYplAMsrAtuRHh6rojLdLXWmGz9CwXY6jXaRVkgQSzluU
8n/6vgMtffHjJihthY7F9JzaiDz8N4ZlgjDOBEanpEvcvDc2aaoxG+8D5eexUPV+6S1HWqRUI+Ma
3/THTlhbCXcYYpsSpuW6zIw/yjQGZ3IYz3fJnktnQFgoGT7BirH+FHryl5Kr7WdeKUb9JqtaO8e4
8GbOTk7Iz+AZqpIPf+3mtkHRAPiGk+3BrP7MfxZoC8tPtl9dpGMeZPnKf5348MhL1maQ1MuwYPyp
ktZacke5YXdDS7RzvB7mmyxthL4pqpPttE7OdIZmBVbNChuUfGjP15L147EiWQm7AnkLDsIBTpa1
WAPXZLQZ/pGpqYolCChZlIeAaiVG3do6yvI7dgGdPKQDbCj7vTF2LnP074XWLGlLIwOT5bwn7BmS
s8MZbGtl+T+G3Cf7MeEwu5B4U+qoJpPrbxHywKO9lbeJH0SvNLCNmAFuonyzNixdEYSriavNRiWV
8MrG6EfJF3w+1KWaMTg/E/B535Dpy6sm99JnWSBT4T7eCKNBaq6z1ysZ4gZeawDUf8KII4+OVFOw
SMfHB1jT2okT3eeiDlYfeRVhvICmW/ZL+uYw9yGx2BAaBBnNuzObuXKuCyRcq5Z5qvDS2iY6fGJ5
gN+BRhOAKNSN6bukOh2xDjx/YbXWXyp1AG3cG3MDJx8peSSpjaVn63kFQXT0BApgASnXDWKxkvNt
SctHg5O0wGJc9MqYyb7L5HMZzA+qUEP8j9nIxI6csban6x7I970SrLmgapI3pdCv8GBlhnjok98J
6EpuZTiMI0PjJbBCm4huC9ftiXaasymJz1NN2gi5pWuxgxTF0ublElBZLGQot3IKvEZOJrbalBFr
D/koo/GPi4GeD6H6japMYcEqK5wVwqCu4j0AnlanC7fUqjfGupwtgDPuApR9GXxLv7V+j0NzbIRu
wyPNmfr1ZoqGTDRZzSdAsRRtcVuIbUl00L+zK7CBzjPGn8ZeS3+0xgQI8XILRQVq2ODMPdZVqlwa
hcU0mlGGdjTfIZwJJVM8kI/7S+Ijh+VTVvqbpLY55ccaYGODIzwuxSof+vgFrSDd0NCzTwRSFyt9
SDJnm6xgR8eycnOM0s1veSw/JhpXIbCwEe2aJXEtg7yLEX2qFEH5+YmBNqKibRYzaBWvmcepEG7/
ea7YQcSsaOHKlrqka0roaSfcV/FvTtESFFDeHKfFtijnTumSPauLkYxhUBYSArLhntRc6HdNkWF4
tmO8ATVR9wdUuyFoebmQ/lxmAMXcJ2KjFcTHLW4T2CVE4ejix7dTe3xptBI+DpGflatIcebwDKcf
QI6vCi4I9jtAx1HwTgBNa4M3cOFA+S8K9Cqq6aBYfXlpzKvH1XEKCHjSofPgbzxDX2ZjoOagV0lz
2NjRfR3JHDn8WgrdseP/yxMn7i1czAHdmgpnvobWsqeH9XCw/LJ97hNLUzE0vh48eVprUH/m77KR
P6xt+YdaPaNcFX3w639vvLG5tpa768NEBTQcW8i5sn93d/LGrJ6aCkCRZqPisiJwadGr5qkDHEyx
9OSqvGACXbLYUr+7iBcGwOJikQ299ogtFz1xcMlO/43uFPml8y37yApTg3C3uv/I1Z7mbCAsS46x
y+9BLWvABs/nWb2B10tHmUwR/CLpZwUFXVxgmBeHr8X4zbOhHniYdqkpOGCLoYa3Z4/macNt0tUE
QR0pGuULh7mf9bn8wzfeePzm83Hlp0vtO3o/gPj2jESyn5C4PJqaBz1LmSf+ctGho2hlViGVg7V3
o22jebYDX+FLJ/IMwnL5ztRnkqQ2gBnKiyVSyjzIlkulgOMaokQolH737r2G0oh8hWCNRwnRA3fI
z8j9NygC2T3e94Pbq9DKRBFZ/xqnQiKUopcY5Qg0YmbDur4yEvoh9+aiFpnlvN29iHwCcxoxOmQZ
VHzPIa9nnBUALQ0I0o3oFc0FuUIm+BqIpZ6Ug7etRQ1zSaYGjYIRnnBR1KW1pGr3WTUaBhr+MRRg
i2QwrULGmKnTdqdL67tPsXa8nh/f8LGqUaGrnXbFoJUETfgALG+gR+4YIkFo9Cky4Jr78PdvfGP1
tQjQ4fpuqtIjtBosUfyhoA3qaWnjiHDkdEXvYhYLR2PRDfARgNv1F8K05NlCoMzjsbhRGTwp9Iri
zdKkC8vF+YRqulhv92wxMtnx4YE6qUy5tPu2QV2UfhtLiK/sWf5hLGi5CD1qqFHbv4405sW9s65N
WvAWYSnl97CHrK0yLhDh1DJGjZBOA0WHDhMH0OjMB7eeQmUoDfqCWYWlwjhmnnjOiHCHaKjsaGmI
jT6GFvblYwBHFk4op5KRqAtjc9DCHu5Lst+vQupbMbqFRG0pLUqS1100i/H4EGqPN2W6tIi0CAIP
K3+G0LSw9FGlgM0dcOZuTci8me7aWY0x+liVyXTJ+CckrSAR2Zrgy4TjzIj2vNM+by/cdA+OrvOA
OB6fpY+cswmBgkng9NKKGpQyX4nxRR3nTEtIzdB4AqgsFVuedp9cnajeIC5uud6FuHX57ad0k5P9
PFLwHppNkJk/etQpzRc+zAgnlcQNR3xsMNHJshYzpLd5odKQAdQDNlbwKP3/nbmLztKDuVCvZZDa
Ru5AbndOPs9q2hSn/21I7UBAK22PNNW7N3Rg0uCLvuEkky3/5nwgkNT4dQ8O4I37WmtCDtaULxy/
bJN54BnnNQjCI90cFdQxHKa5Vmu7Bh3mucI24kWq2UZqa6rITFAxNc6unqylIfxQHdo4H+8wLnco
TZTfEn/1rjGi7aDaugsq3lnbMfsSK2jAw4ZddXp0GP94TMkh3t/imzPiLb5mzqrRE52GeaMc6l13
pCuvncc0WCzHEG/I2h5r5GBUHQ6ESRYHx16u4W0zV3COzoGenv8J9kF8lJA7QfIYG02xDSaY9L/1
jDnTpLMMnzWhqS+K+TDpsHQam3fnMEVNYfF2CLeA8g3wgVxUKdZumKi1j5TEHPGMhrwod6jDiKWC
0Qba3u3y0xjxmNvCM1NGegQbM+wP8gwOeaFsCTRl4pBiXW66xp2IrkodKdOExSg3uSNihbFVbmLN
XqTp+whFaNsdRF7zHodi+ONFCOWrUH7npm4ysUG8V4MwXtMep7ThPB3eIRrNucA864s8CVHSZH6J
sPN28aR0549siK7tEOK7iUBwNYobhRXaBgqwXbEqIXyCY0jY+dL9qGDNR6XtsIr8hkgS4hMR8mJy
ZfcfGrlkJIAu6TdSvacsbBSYIz9BmYb5cwMGGlHr6Jm60DuZcBMBwCCvJ1XzWYsP5YhRpVFvNhyM
ZlkB6PfLv/46zTC2LvGolytWbJPfxAoLa5MhOjURD2WMYI17YKNwrcLfKrxC5B3N98cldG/WF5/Z
w28xZY2WE6ghtw55QSOk1/uN4u+XEA/ThVn3pr7TzikPM+EREMoHfGFwusldQeyTCorIuEa5v/B5
XEzKrc4BBqtg6OzqN/orPnAti26dJagsf5YXHih67jgs+b13vJi83q9OvZqI546nGFQ4ArTZ019U
NnDYsdkuzQZvOjqo7KYvVyybZl9JDuTSM5urCLy4Xz2hVTQJ2lSN90KZz/uKg653Nd2bmgJVTyCv
7Yj8lvKbI5Javt7VfkM6LsO58QGrSqrMBHQHJ7e+OwtFKS9+Kz5c8JTALR6Un6rtATFZp72eNyql
+oYKF92fbQ/zNAy44MydCYAVH32qFItqaDqz/sP6RCFp+ZvLYuRGi/2qS1UYMTCezl4lYJ1zMNpp
vzAsO05gl9mGKS7XXl+PLEdjECl+z14AOGmnEE5D/ZlGHkQtm0V7fXjm5yiQFmlJgeZ3xLAHpOte
9cewEhoU+h4c9SV1Mat0Wno0kOO/P9yNAFkr0c0o/DC4YUC4/YdqFZH+QIQWQt7pPFw785RsPFIu
ffKHmNBsoG6NM/WNPhkInaty5azmBQbbLeXeZQ5DH4JE7LrhBSn40gNlEOO82vRbtrDf14nXKMb+
nS0n5TzYSk/Y3N32FdH9ZaoqWtppos/DwsbbHNyQqa7N50zUWou0HotETWf+fjCkB6mScKMmsHCS
iwgr9llMlEaxOSlA4rKWvQPh8Z5uDgsgcsq51O1jCJy/Rp3AondLhknTNQLiWmOl+aM3vOC6oj0f
Hz1V1jNDumFtFZOw1pbpApYpDWJhpY+yAomev/4HiOgWm/H8HSqdbSBpi7Ba3yoVItPp6apOJIa0
V01nq9efic9DQHBT3fvzbv+VIPHvJMr7bNOloCFjHa0jDUU/4+Fd9f9wMUnFlonB0crvYwSiDsEL
ZRmbsR6XtubxGP8UoOJxy6w1UyX78tHQJ9zV/AvThDC5Klw2hgSBYRViS8is2JSMbV2JdcpFx6tH
cD3kr1z+6uG/kPlpGfEeR0Gbu78y3ktzoF/zaKX8praLXBv4PvUtLFLFGyS/TJsyExwKYgA9LkwB
u6xmhgfBz3PX2YqnzJJoaf0tHZLtK87vEWwTwy/1/AiX4idzmk1yfhd4KeK938LGZBdcoGrlJQqC
S7OPirxQvAx4sc6unsxo0+67DVHNB9KXmj/fevB+2bCS10JkQ151GCFA7+Y2Sp0j7kfbsojisFSu
d4cE6o9IqRTgZzwaS9aDie0WpfVIxSHZnOtofZv6Ys4ivnCdnd+tFjedKp0tnwrvNmMlbNhLpQxQ
Ka6+JL2NZXJlpFn0QcaX5llfClyTD9YeZLrVgJlOfU+XwXtXtQY2SqwIb+lDqSdLLtXRC4RYF6Em
hKqYlOqVX5986D0/Gwelm1sRy6Bv8UqyjNC3RN2wo4irp4N/Q4dNog+AkM244tiiZ85iTT7sH2FE
5GNoPzdnVTkl+SQR2RSrZH+WgCYQIPheG1+mnip/iYWV5/kLErnon97I5zy6rpMv0VVGckghiVIO
1q72xcXcp0Ydux1BR5d40r48nnnODgRhl+K4v8Kq59RL9Va9q++9aUa4PoYNBNMfnLMyOayz1knu
wRkHeDfAw0XmlxAU0mXIch3d3HUOyT6yVvn1eqhkWSB1VsJQ7CscVgkAEJWFo7bd1QHJa4mk/F0X
jf4onjxg6AL0/HjsWGJBDWv9AkdzaP8uwWh+rsvcA9SRlJKlveSD6/qTjhTPpiutAyy10xvs99pK
4kqjCy7ILK+1b7xxq/dWTztBGwghcc9RE5+IF86p5dqgugPRby1yvBv0rqiZ4POjy5z5kIbn7kiz
7L2wroHgPrGwpC+091XgbbQdE7zTSAESDsE1Pa66LyHvUvkdq2z+XBuc03ceTMqQaYIMksq/MBVM
daMJRJYb+2rmyREO50I2cQ4USOHXAM5KeJHMFAmgcW04ocydTTOBEwcTYT2Ml3elKWpkRmT9pzVj
F6H1JnWrJi1lcRKzhXeEKdpEzw5G+KHeji241W7PNMhvdilNTNvmd0PQFdPWcJTR+VHOe6XRZrP7
utLIPEjMkH6/zOgbs6xPJ7vA9kBvF99hR/l4Ur3gKgCY38ysxtRDf483/G0WcXGrT3jSPaBChpUE
l4d61dDzpg1wdfScGDsW8/m2h+C5FsiDR2OknzLeWexNK3dZoTIUgmX/XjHEvvD3mN+irGSarUxb
4logh5Cg6AX++jcJz5yBfnotFxwjRrYtHrn1QB9ik+kIyNuqtmpbfx70zNJjwErXPS0Z78Rd0hrD
ocMKZsTkZqOzUwaCLee5pejivWgTbj29i2dAVcKYZG9gTzKSC5GGPsvzbqTd7rwQ6fZ0sGTot/pL
5TiywJ9D1R6nwNuuuECdR8FzssvYGkJqiy7IueAOPZylPmcxv2eZr6b6WEuzx408TEwmZBClH9u5
nBPCb7wjSQfi+GXRBGgW4flOJv+rGtFX+ntUQc9WIwy4eTePV60aR/MBTdMlaLAWYPdrNjcYfyGH
l7MBJibHsVpPeWjyszEBAT4ZocCE0yCxItPpmXRKM8FADHS9cotF2lpkVODIhFlCSoAe0JcKiS8Z
K1eEWkqFH/PrEYkgvqNDmylce1Yi84xwN47Qe2xjIirmKkOI0racS6TwaOsfhK4hpTcRJMo3Ypjb
X6m8LyJih/JzHO1sWlzss0uOtW80AFN82FZ5wK2YKqBduv3mM2usTflD8CjS1GSc43zsvUJZ13in
CwjLi8Ye6c7SKOJFurV6wJSwiF6sx0+FmhevY/vq3CMFvCXiiDMSlLwereXZaO+62DPDqSTV5XAU
rUvpNXKnKCFIoMJC/j9UsKinD20hFdXH06rGbeF9G0pgA0KZ/mXqGR/6ovcECGoBbUAMnBbp8N4U
6BBvygXzL8MlO/whb3IfsXan4uvYc5S1evdmx8/AlzgnSGdO+mObERHYV1eFafqX6Hfal1F2ghdt
ABBfDIsp8KR6HLA3BaKSNorS64iaOgy+OnD8G6Q9fh79W5zR2daj1UJq8gK+dObZzbu9yW+FUOKT
DIWlR72AKhujjO2vkREiVw7M7x1aWe9RDj8Gt6lsZw4H5G8xqiiquQ/5Np1orpXRM4vRTkj7dKjI
VQ8cSdxk4REexcynvKmvaIsxm4WwvMmzbWocBIqNDYkGYhbWLQVwK+/UAk9RgDeInl/adGyRJRQo
ics+cpjzZ9IleeSCApso7W5Zk++v00C+m+ssh1wk+RjV6PEeZN8eMvOub3kl0K7ch9BNetnrNUUy
oOtT5fQoLvtGDkGnUCavVCQmLUZ/l1wXwGG/Z0xvXdE/exlMZPIe5Qmvl61RbzY2mnf01b6agzz5
Dglv1VTLySR7h52F7Ml/PnsdGN0Jfg/VHIyf0OANplcKQdjgkDpTLDCeD+CZLN5XdZaGiVmKe84F
crSBwtA8iEHVjJygCi4XFciarwUkXzgfeHYkSqWwJOyJ10MmRku6JTDhEDHplkw4maO8w+fOmkB3
PL4//bVvgo1jl1+7RTSljEAtH+rG2S8/dDEM7ZlxHXrlwtLlSdwWVSLFptVsf8aVSh6GLC8+xYPs
cwTtrr/ituhw2ZpZzVnHKXOMQFgOcLwTVOOUUeJrGhDr4F1c4O+OrcGGAay0AnMzdK4TAlAMYy/X
ct2PNuSLvXUTv2IpgvnYJQc+lL6J4xRgxKn3YximCnjWvDGl0z/YK1G6W0sxQ8ujOCML/lrVkV/s
6XvNZfX/Iu/p47x2oNpXrEdLWYu5GCH0nc/SBhC1dUM9T1x7CUQ1RSjaKVXB0J4EAHeMVTFEnC8w
LB29sVu5Z1bhzSJHCxUznZyrxRqRHdXMNbtghUuOkU8S2ymfDl7O/OplSnLQUZzEszuIPMgMQO48
iVtZoI5AA9WvmnQlvPP5saN8ZhFlyXMb3qM7zwolLDsoHbd044Zh8xOROhJz8a+LQ0DULUFrCZLA
3lXqKHyoAC3l6qocdsFCmNuCkp85TQ0KxPZJEARReDQBbg3ywHQZ3JGkGU4mCa+mMX8aNm18pXIq
hWhT2htF1L2Afd7iiH6OWBnR+uGVa8KgpDjJdqYR8Vt802iMNOMXtg9e/N+85Z4XX5Rr0FoPeg5W
i1WZxWGzPX6M/qJ+x1pM+zHyTuVCx2wI+eBnObFKbBkn72SO7CCFIXlyphbBelY6BUkie3Xh5USw
ztRu/UtikQqvE7SRkXpdgi7t2LBFKufYaREgTsN5/RHmnjit4D0ZDKEkZcPzCLI984VWC43pITuV
qMy/pe7ut9JoTG8qRyPQ0JIZ2DnKIlnjVhdo/TNkMg0jV1ghr9aQeydiSpxS8sGfEUpADQt5ac1B
AuXGFUKnDEELyL9LGy6DluR1jcH53BrOzE9XdRr+F1X2YjJcrNmeN+P4K9jNOYVv0aUnT+lZnHpG
ABC6Xvo+RbgUXonh5YSaXxBFZd9F7VUAdd+ZRt8fIQhSN0vPhiFAoyMKTvvzD+xxVXGb4Xg7hnNL
jqO6MzUjaLjPQ5s+GnjYFGU6aJBD09W3PlZrlgxCCEEtlWjruvs5hdJ2H1dm9M3hN++FlsdtLTVT
0Qx3175fFCEgYivfkz9LKQ0nzWw+UfCVpqlbA0MGxMZGGJUJs4o7KoR8ExH/lRSgR3AtUUmfHvdR
Jur5JKJDZVKPROZiacGlv1QMSgfbNO9qWFNOoHlrzUV2RNfrcwsqR7lttXVzfMppOxivIRvyUOEo
2FbM9zm3AvREt+FeLMPK8Qf0akL58k1Y9H0i0m1tpRKxlj9kFXkX9MxfNPwN6+llqH7IZf1rdmsG
uZniiloxWOjjjiRgDuUvsmeOAjM6ZLmdI4lP1X/TGNjIsIVKkgQ0LBvuS7qPeCyYANqibvibSQwC
EqYoqHlZGlwonEkfpscde8KXJaq2i1tXMJaKiOYJvh6koJMFgw2ETWblHoE5qqpoBZpHSjhasFtB
e1LDx3O5j74BFcOac9zd86c/u7xni116P6w55j6deCLzljHnIYx+0BgZBvzI2Mt69Fi1XP8lcr8G
JGbntpGMYyaeyfQNNnDOOdOQDmyoo9Mp9PZCafiqDyhszuxCtwP0pwNvIDY1guSJfZjgyj1LhBxf
axg5Kbl9JroNnj0+5HDvNg5qTSBEWlQfwAgUHzTqOTG0JJ0P6Pdgv5iSAxt5Rl1F4GipMGJ+ucpN
VIlkvcIo+15Dn2q4Q/saXnYy+qnNyTEyfp7rHU1skP2qS2K3bV5F8sBnULnUyOWVbLOsKYR59nkX
dWK+/jy8+GHpMNn4Lj+k5nfBdHtpo3fNzy/Xfy1nvoWH9uFiED+Fuu5jP8zjG95kDO1YsdEHuktW
RCBlCxHqlEpHXl9ZMADYudJgOUFiDl/eBmNl9o/cf+4f/UJPQrkfYQ1Mk7CnapQ/wY20rXQAdnfO
6NCc7hCJhH/XwUxifofQDE/FHrdB/5Ebogf0PvS2aoxd+cDMr0mLjH4awXuv2KDrNyd8bndh8u5D
4VIBzZIcYJMbbgcb2bXAzraTgGhPGE/oRqALTgsNyfDZHPKRlRj7yDLY1F6p9O1sznj/nkwhkRTe
ordb++XDPj3xxVK3WBoBHNl/VZyZAPTa4+lx+/ALh5mr/xGwtqlVBjMMm4tdtmU+WzPYpltKT7mF
5uDxgF1HlKHBaa5SKKmcvh+tlDZSygRuWCKCOLRAoBgs+vVriVlHLAJ5rADnxcx2kVflTMYk1wMb
cgvtGuvuDn/MwOjyh7jQls6anDQL+7w+rKyahEQ6rc2ZOou0SHoZqqMtFGlB9MsVzn0GcF1Ya6AT
eSH2WWdUAaiCIW6go89XeMjM4ngMWbuIc4wF9R4XIqzQor4eu6YNwcAVShD4Afs4PK24MBnRBkMG
ADwAItDdnlo50I58CUwJLEZ/xUcQ9OQVDtMF/n5o4mgOIb+pcrkLtuO/0pSF5r/kgRoKjJUAqqSI
7AEoayY/04AB6iZnhbY9sAv8U51xNgxAPT2hsldtFmzTQCHWj73YxExhnH32lK5EJXpe56qTZ8Xc
1Tl00ex+N0yW+jPNFjrmnjQmwtDfmSnFswnXkBSzmq2cyKeUp4JajdJrpMJUHpY5eb1HsOllF8tK
0xLzGo5Foe88XskoLVrBR5nn5SzMNVLYqGMnEQWXdQOzRZ0I/RlvTmTV54x8VfaNFskygyprLDle
f5qrFpxo7s14/lESw6xGVzL+4GfQuM6fQlEb6C4+To0cdKfZf6bullcS1QqmwP+0yIuLZWrvGfkC
jX4nwFCj49wgLR2lYsRxeydEv3qVFqvh1NFFYcvgWgXESlWITjUMdHp/gBoc2it5bHhvzVQQlWrg
/bRw7Xb3jjIvisV48sc9lyMCfxNuryBSsr/hq4hMFBznIERQZqv6MZW11JC4eE8Ihwkl5u/Tn+U8
19lSpfaLYjmWV7ETWBXTYRlJ807mMoYsPKe0hoJIYd4kA9aUhSZ/jv9C2nLhP37uZ7tV3MXE+G9W
x9WpWHSob/1KZy30AZrqVrJqxeSWhCuSvbpBBt/woYPAj6veJXmOiq3XbMO3kxO6wV+Pmf6kKRDk
a/Aslurhf4/bGGqPFeTDiu1HUBBnXA08iyN7MknUj8nG7mPzfKQnOn3Fq82elQ2OOdFPKGL0CbtZ
UpokW4w7gO0RobxO+1/2DIhvGN6xfIlv26V8ZMd97TQbh1p5MMmiMb5kFHYg7a5fsh/+ZXA6mvk9
K55MH2xQjLG4kPWTbtoHcIHavK28dvIzoCxZNze6wzJo5dTA9uVeOVE8hEKYdsqNJzFhCDHHwjCf
msus7W72bZEd/QuCfL2l7VrsJ5X3nF+ovqons/kx9ExTdlc+YwGM7jBvIjAoeHa34Zuy11Vk6X8Z
oEduKXByE36WGCCUX5fQDVL/kC+tmFdUAlbwEvLCadyfgUweH0FiOD6McgrZJJ7Xp04XimSVdbw3
qofQ/97clT9e7G6UXqgYlxsqsj+LHk+2wGIJZjr1vYGuddED6NOMcxbL7xOF98PSrE0NZXKIh1P8
tu2xlt1XSejWjFaCkoUwP0zP5IiSqVjmVOQda6VX8V0iLe9pg3jQTBK5f8tuuBeUHtLrsLe4mnrt
l0qXrqDHSje+K23aueepc+x+QILbfOJB/FNSXogtkdn/GqRp25kVkfyKSgSy6ssUS4fJAB/uw71C
/n+V6b884Z6CfGy60t8+asT8ysPGzg3t0ye0HelNxUGfhRRr4BK+KmsZjyM/uJ85SbjkT9OOwCal
j9id4+bNILtPNVIBStsudbHQkhbqAkLRHs0DdHe0tOoZAAUtN4Ut1LKsLFPzKehQyQeySwV8Af8h
Ak6snwi6OsINZ19OovJoB+rKMNrVR2z9hn7MgVndtYTubYpXTUu5zGd+hRNIhfnFXg3YR5Q4Yh7+
ClGySEKQBEwq2E+QhOkcdJ6AXddMDyvuaHtjCoRKMwHmPelnqIXFqOTztZKyfAyWkRZO6T5+h2XA
R2ly+yq6VbTISCEWf07A2nKm0Gz3P9s+zYFA1SFh0kakQEY/SsUU8vz2qAzZhaUDAoTziXIhDMVp
4c/HHomy7+uL8cL6wAJz77AnDg5rHuscYe/s1dZSuK1MULBkFWEu2CwlCXudi++gOtFGOiPCO1oP
Vmuqhpd2voLbY3pwH4lFmUEyli1S96vCHOjImBUt0T4Upt13r/V0S9HEsDbtlmpn+WsnKtQdtZA+
JMJj4YYYhOv864bZDIuUQ8miMvhchFj7QnHWHp/s2GlgJYqtjGQNOSAojHHIcSCbL4usX8Qzf/cE
KqzcKE1o6tzdAIwDhtL01x80txhSzHerexPdelfjQ8rxq30S1hYOXDv8aSNFApLj5jfNIR7sB9Se
drxjT3BZpZDYfjfq4FBqmrWNZxaH9p5FE7x3b7xqB9Kc6CO0c0pqbtoHORDjiKChYmVw5/7DYB98
HqWOBqqqyyFrEmhUmthKyxtRBwNESQIF6Umhav1GTcn0iq2MjtklV/TfrXrGppw/IxH0Y/jUipoY
oPNYXWSh+uRXEQ5TX3h5Lf0kyyvM2D4pbu0SGXwab6o0IecF7iTTKAlw7jHBqZ5lGptC10NIdvJZ
/Y7X7U9Z+tm33NR1/b7x8/KJxKuufHZKUzQo4yo1wd29J29VlpIFIHDvxQ8lpHZmmfekLExeCDoR
ml1H15TokTEba6quon/3laqeD5EJTss0f7PVUGHTm7XQuui5dGL+oMhdbrULz9bCP2lkUxF6Iqsa
Ljid0mdOdbC/ODxed+z6makMQQ/nVjFjlqX5JdFxiZgOhXRrM6Jv/9vPfGgpuUSBJs+1+eOMgQhd
RwpKp9/IAnCBKR0Yt+eqZAT9sX2v/6o/9zQUZZKBouzNirXW4cFD+cqyltembZqzpMD4NTXThiS6
46ZeLthaa6waYrYWH7l6RwRnfOe85/AJ7fXYEr/tjjpBgiOiq6WPKf0iUksVk/9AxIZDxHu6/glb
5iIp/GIkZhtpCPJUEP2Y7h3SZtYjEtJM63U52KO6tI+IRafBLwilLoJD4v3RGYxRJ0oHkp6vum1v
sgLHqQIrR4eSTKsvUOLcgMwd/0vhtNOFi36hrrvbMb6QkwelDQLHfInWjsvgJxMHXB2tVsgzhQ5f
nbXWuge5vqUZGwxDxW+Eo3k/5rdrvlb3vnA9fDBLjR1eR15LU+/cacK9t3aFNHJCbX1GNmz3uk4V
9EIVZLrA4vVkBxmBpSIZ/LWyQDAzPINrloabQrBuMEdEJ62o6TM9f2OMlzy/3R470MXaCRgpAc7Q
JcMp+iicnYLPwThAAvtSrLVYuOh9Elw/6GfUJ9aQlxTJmX8rqBmyP/wGrfYH8pbnsll091Jy2rrL
tCkz7fLzFM4+iJHZgMMcM0QaVSO4SvP1wrBU0NNX6h8HUyPZ+sGJWDYCK46Ue13iJoBmkwYQZFKB
SrghKJzO7f9Mbav+q64BqIo74gAB7n9Ho6yUvZz9hZetnKwPt8EvTPI5sEqsgAAWp1WfuXq83q3O
O1Tx+mau+ewTvYnWn2xE8CqeFrGYF+KWqisomK/ix3AwIJ4tlxhTeUZbPZfgQg96sgk+9j3oiBZe
Z5P1jHsTZ91faVVybgKcaPtTG8gF3/tHD3lJnyADzuW27P2mA6fg6vM/aCbipjJHoXmuycjmTTjF
9xpshycMqE6BdDHkVH2wgjWlMdocMOJ2UAPYm2AbxsgwhKk7wDn6yShod2h04z4qIim4u7tthAq4
i0Yn92A+e759rz4eokfzSR3/jnmnwFrsVYb2rPOYjIGB1OSi5OpbDq+r6jPYlEK8auXHaDyeOPpS
0uGrjwpAP7XwuMBE8bzuuO2wQY2o2KU6i9RMeD6JQbMeRW/QB3yayBtGTVVa5gIU1zwn+KZy+6i/
3enwFiYwxD/Dx9ZY/4oHNb5aCI6XXMr/EEP015ej6ejs5sHokU7XjwNmk/HotRV0Ja426xXaRSRh
t9M7ZdCWFN9Jo1mpE7v6XATjVzPHun7tlAANCL+ITa6XUMobAm30s8rYw6UnwsL0x++c3I8wqU+B
khXrI0X9G8moPLICrIAh9wY0wHCS+MKG10HBdLXT+7j8b+6exjqU4CyX9pSgaNEJOi3HNcB3P5sY
cSyvf1+7GGedh201kOr2LjB9U+t1orbwQc2p4TZ7zRWs4LgCdxu1cjqYCWpP6Ct4nQUp4V6HPcS7
/ptGw5dY0dW6Nv+c4ayl58+PRKyAmWmpBgjhCAxmBuYXnV761pDQX7T1zttTWU8zmZzfYCYRcgOi
ygQ0luoyVURMG8Yu1URkqBe3cBsnz2g8YibeEj04+2je6NRwfyk8Ut2xjLVoYLYS2fNnmr8ba75K
KqgSQW2GA+nrA0pOQa8nJ47GgDQEIXxnauq934pgTdrfXqLDdaOyoOppWnVlZrMHmni1JM8418lb
zFf7YMyByG7wBdSKS9fqe8najE0QPaCqxEHqJyCYgAzklsyrJIHqQjw7popog9PrJL1Tu0PnSqR/
2uNJPpx+DuGqBCjm3g1b/sZUfNrDvOa54s4Nak2jVqXlqlLtDv+b9FgKoN1nPOwc8DdlY86V/mro
LLVMchi8IMjAuA7EWKFYjZQbwmesDQZiXMpNpwmMmYd7bT2rwhpqxcwker2kP7TcIUCvnMgl1T0z
QqUTNxTB+TBqu7pWWUyTD2imAKonvDFdV/m6n6DbQ4QQz96XpAmhVY9V5dtSrR2YwlCBBxVYYhLl
cSiQHdZio9niox7aXlUAAJryJ0prjqF3VYgxphdtn8K6AeTYUbtK8lY4h423VoiFusPHQzdUyz5t
AMVHoIzGZRfWXUrQ/wQhFuIodMWf2W80Rms7NJwMnujiCxTbiGkgz2xNFB+i56OlHlpmZDxDikDQ
YK0v6PUrpoOvPq1Tg+zRA/jMcgkZnUa5s9+q+gTQvAcmCFdw3WGVQ8CeaH5bjmajhksd7DFXAVi2
ffwXujVnVqMYu6OFt4XXXbQFP8bq3yWVH+373KoVaoSoy5WD3NpIeA4PcOSYPIeQ0fKWhTY/4ON5
9NvizsNYoOC1/lBKIWJNwJAYaVfqHbmiUS9tbcT0fNSXRAEvBBZFxtYoBAYK7XfmAlu4M4MxFi74
Xw8hq4YJ7uduLY4IzZajz9FI/nosvSKK+6EDL62sZwgih2Y8HReR/Y6P42RB6/A6MGQdtTpHAFiJ
lj358h5f9+a7XSeppP0JEw/f/Z2zIiBTzxFSkVhrkOZqs3JvXvk7Qhaa7J9N8yCNNzNBI5QWAOmC
UYIFbs6Jps9Y0iQI5sqqW7gJFa+u8i7DOE2XZg95YznybJXSE80rH8i5DxuTGleM+6fZZ+8HVIkT
mxM7o5I0EHQBxx52WdZzTcyzUmZVgeobNgqw0zVclmudaTbm/bTPgVCd23d6jmBVywDKdnh/lLA6
TXNF+FZewT2xLFTHha0S/WUqp1AiTkUgTXM3w7ro1hYZYem8Q1672M8Q9gYnKdOjEI6GGVq5lgq0
LlE1OlhjOfKZ4b5hNABsNmSncq1jX1Z2p8mAOXd19t+vWNV4tJxBvIGcUww6q6xbSPYJm8M5nC7G
FWvGEV/wQziJQ0oOt2qIw0y4jevuSQXaFILvRZcDoRZBz3yEyJ60RYMOvSQ0AiyEPfiIzmN45UNn
eeAgeYv1lQygU19XFvn11FJUnXIWnJxbVO6Pygljuh9s+ULY/RxelwlRbniCcYywAGvazuR+wea4
euNNAi0SXdTjyKKwwxJxfoS4kEi1IJOWi77aQDRJ15NtWFwHY2CGJFg+gOLwUXLZPvdsgXmBuqJD
fIg8Y0tcme5SOxrqzYgSD+y7ra2dokt9/ozqZfeGP1WbN45FSujgO46zQIyF4aFrfl6mRGsH3Gl6
pfy75U/ohfS+QgP8CybGkaBxth93YYAEHwaH9d1mbrXVasljYjKOzQK5bzxmRxfA/0XJh92OrI5H
09e108AwstG8PaqHbr5gBIApj8fZE066fhNpzy96SxWdFGCdSp6xMG0OScEyvDmGnYiD/E+NZiLZ
s6IRsvbSYb2dm7D+lR2O6ySi6Wz54zkQ5Djx6EhbVKX5Ohn5h/XwRvp6SAEObd1K/j9UnQjj0Zmi
tesEO3DY1HkfbOIECgEe9JyWZuzctuI/BiOutR+0xy1wHRwBwjsc7vuByvvK6Yur5PJyDFWDu50T
0LGvBnURrxLbM5Iazlv4EgiBUysCvfBUCtpLtjTAQIOPM0BVDcA+ZEwn0umFtYmqPswDaVjhylVR
PGwE2RXhe7s+YqNTzyRtxr6i5GKV/UVpLoMnDUe4xQGpqnOnc4iPCjYeiooSs61YDNpOfVcn1we+
LHmhPRS0ENwTpCFmN1FUUWFrGkNak4pyKxoPjjTJlq1EQYyTxtWxKFmEp1g46/YT/D8TfU2dj6Qs
HsqeNDtJt8zB7+XBfDHP29lWsmOuEqbCbxkTB/Aep7bz1XL7FVUmWFnjckyD8ZQad1K8tlJYowQQ
e/s8Y1Erru1mIlEDmTTvNF5YDvgPge0VfPPBr3AA72VF/+mbdigcfagQBS/7kzh6WYwjrMC5RxKd
Oe4r0KMW6zdfVYVv8hDoIqI3nM4aorRsfwVPdIPLxTwxRLzm5VmddfAGCZavKLbdrLlIR4+4E7Uq
HY1JuOMrNI4PaU8WrAguLSaEp0JESAdPwizSzuBjqsMVop3x1O6tpCNfzY5tOzJPp6E1rIPPmD3a
3JiJd3Cl8HbVV3nzBiMiS4yS3rSwWvgoaTJSshno88b/HD/6rSKFfIx7nphWTwjG/mEfJVzbJ38M
UoeFUVUOMm13AHHbdsRXx0flt38C3nMCkcnPYktIbVofxKn1lJG7TDK7sSaydIpE5cTX+HirX6e5
sgZMWIkSse7/gc1YhFgz7/o04c4mLyOFJKH30kNzSn/+3TjCF932rzx3dnyGY3PVqjVYLO+yJuvR
AcqGoY+KrIVlVoE3Ywok8t1sXneS7gLkperz5pY+M5OdEa9TROQL8qbCohrJJRGj74qbugrPyKdk
pzGCyFolHt2nckMLmfFPJFcr4sgjKoWrUmHDyHvcuNVQArUD7IVHgkfX6Nvwi6TBUr1Sidw1AzQv
qUy1oTjb8KZ2x6bP0ufdyJSx03Ymzx0/0SVc5L2tsDDZL9+bHqIgZ9Bjv1id42I60kbVg3srPePb
YHdFm7lt9KvNPuT3hsdb7X5N+KGhHz4CT8gIgi8PhGouHJnr6Ep0Y+zfmp1Sjq0o2M1qHAImhYz7
cRuz6uTbWxMsGFwvwPZ/A8NcenY1PJr+YVy8QKk0yXvvlx+tXQ9xuut67xyLKQvjuGPN9ghy5H9L
VDWCkkp5DLVBkI47nAO8t4O5+fcyxfQTcR+tr3N4x91Uwez2MGqNjnH5uGx8kPtkn6VDs1WCm3rT
DdbBtyh/pkG8BfLqY9tIRUdbMZr1jabWxqup9WcJqMd2DRLABzX6ZJZxoof9jXmsUyb5tikrpZqc
t9t48idTWGGmT2MRT8B9wqPv1O+ygAWpVJWBM3ltqeXmIht3mowDVfJMrE0jE2kz/5JKOvPo0Nxa
yh6Zb7J8LaVs6bcmrYjQUef3/88sB872ke48CvSeEFFpvy3BB0N79vcxxvZ0pOlSvEgbp+ESD6vS
V1vioYWLc8I/k+f3T0JOpV9cdTYif/sn8MkMKgSKP9BYLYq4io+3aO9eg7Rj6u8W9CXpyoestMid
Wa6QrHstg6OcRbuIZMVt9X5anTC2H1im4BsFobnplNqcbla5H7jdCWR2dQ89wrttr7Ok39mLIG3i
Hefr3eEj9JFyfH6qq8BAs0L7vgHyid2QIKQhaE8py9JARSVg8ZaZerID8Aty2svusx0OLjGJgQEc
D0PwG/y8K7nLaPpuGJ78IXTbr1Aig24ZiFNkr/pI98OOcdKA1bJdoh86V+hkfyi3rjAg9ljBLDy9
hl+dF0m6KTAl5DJkTsPkYfWL9Etx0kfxh1qL5JMMxEXNpsZVp48JdUAoEZ04HzcXh8IH8In95fpq
YG3w6EHdMGm6Cig0ZOzD9qQzQSzbUtMBvMXtDyI36AgyqmsAdb7c3h7CydWigvQPigvaphQ1ZLaz
EZzpeFYtjLTJ1xwaLUa1eX7GWINTjp+XTlke9CDYhaAiHnx9B81peXZHQSU/NOBnlm0IuROfKxAP
WugLeQODU28JGmNkTxnvndIqh+l7My1tPJn4eMED0v7/+MIvjyHr2u+D1RalNTqTHLOcZr6El59V
k7WFUcEZnchWexWzdMB7cwLlBNhTnVaBhaY87NBm+Zk+Bz2cU7kzzOnmXBDlxUd42JV57g8zI888
X1fbFDvP/zlDceG2c3YHGRK4fnJB/HoZOygTbASPtikN0uVXEYbauToXs8oWHoISAhjuHVxqt6lP
NN7ceLFGLU/zeE7PaTrfC+1t5kzRABIqUY/pUtxUPOWNdxfQYAk5o6sucRh4Zp4H2trJVmTs+oSC
k8hSa2/TggqEE51FKJK1j7qXv/2OQNe+DK+OiyAqJIB5IIOaPszL+/EAN7TTHXPKDx4SV9I4bxtn
WA4zBIntRcVlz1s9gEWUrKf0Vilt7kuMQVLdCl9TvuiP9BJ6ALH2ibsw9s5YmuNoJEES5OJybldM
aK//FNYfhEEhBJX9KdSo1YIrCgiDLeOsYMlV8TNfOZK0/ws+8s7CxfOHBVogszrpuj56NpBgwlet
NrWd5AA/tf41Muss45KOaGvRac5ifNMRB6hOCxf0Eo2MAquyFIijDMpD6V6jseOmPeB2ivO6tslb
clm2fNFs1iVQa3V6idWCQe/V8CvAHwWC3TJoX6aYRVuMlTAbUXZmYQPFSutEKJP2Jc/0xf97jHa2
RPCcT2U2lQB6GmmiFns06YbXtWrMsy3fAa5ZVi0A1xhMLFnzHqAD52Tt2SsgOi3pPWaRNa7R2HYT
2c2FKdFG5NmWB7zP04hQTAgFr+I5KEbu3Tgef4wQOhgraUPPMF+ocDCekbkXmM69BZd2llErwxOX
OPvNgsWJ/RhIV5iZxo5f0JueIVh5wFB+Uo0baZxecU++0tlBxXulCFEPto+x+aSShbCqK4/USO0x
dUvsLvLFhvvQTWc0hcHdYEBf4i1FPJMZXu9mYwhQqO+RNROYGFqPp12LHRPkt3+zMlIFnsQuIiMS
6wuN4oHcTxwuNU4RfopvYsNsDpxW8Nl4pvFVqKNTfFUGeHnCC1kxzOCMdS1P0hQdPmw0TfRqSul9
25G47hv8PJ+AtWTPiQASnok8vzhPaEFWSwtQrajNUTcu7dnTciumDCbmEUme5ZUgWxTBiGlid0qJ
5TNUUdxV1mPHjTLGCO+HJuHRHABLTB2KdiCy3qyA5T6t9QxRVewLNukdYQosc7ZfXVZmLjTlhI7X
1VYaLsmGUAPd7dVZWG+xvw2rhNhzu7G2rtoeho3wBYZBBBnwEBmStpG6uKKK6TihGKeTi8ClnbCF
hz92b8tmlDERtDOvOIHS625mHV3glm4dxcGJ58noajz75gyMz0Z15V0EPPT0bO74pWT9CiHv6Py9
GbO3yQbF8TJ03uDQME6UVjBT84DQNO8IJ7HTIZuzfGe+pPsPMUE133pM7uDteeGbXciyrlm3ilGO
tNEkUXTk6AXRyTeYLw0S2kKwnjkSLkrOjbXSOV7rdZtuz7DxHcr5McCYCfxM1oJZBMfDP3bI/aNW
QJeB4PtC2FP1BdLr5S5inMLmp+8Yh/ZrXDG4Qv8km/2VnoaIf2MV9cY+89WSGYNzqtFrhCJZlLMl
jgUX0ScZf5Mco/aVHAPYPmU7ci+8BWWSD/VJV62YmCyBYKy1PKTWaJwbNV/tFvAxvybavUu223GU
QzcIceZziXijzX5ltN2TzjDvtSbpVNLgewqc7uzNCJgubzue9gr5dwxYu0LFdpzx5VSSR+4q9Fk3
kaCdlfJS9AbUD6LoNDZhUgNhwdIEVVWQ7xYzujiSJIqr+t65DLkG1aNRxwIsZ/1l2utJr9UR8boQ
IBLC4WEOU9zTulCeD5YyBtySbs8APN6pSG+EJTgu+yxw0ORAy2KBPLCcUihWF6zCY8AWGRW6XeFq
nLnKdM3ITZt1FnkSMMLHlcSjZhI4PXvrCQa1lk82aur8QOP+SbDq5Dv3PIerKCAI9ijopA0A0XPU
iUBIrJ5rNQ4lEsMJtH4DvNi5Lo8HactOpSJpr5YKDR1R3JxsSWujCp76wrDaj/bDG3Ab1sbABgKN
0eKFSwT8UXTpa0jmewiwnY0oOX+9GuoPWp2IdmccejCWQ83LEX+4LTX1dTAQwfSDpUFJyuQBXqq6
VZAdHA20lDqj11/V8xq3T2T+ETxOoBTL9oWYJRnTaJ1b/0PtJFTqfFurRAhcaE7Z1sSmlIgrLE99
q0wP8uKfa7kgqM+SrLT27OnCXQyDyHXpA36Q1F+6f/Pn4Z/1C0g12VA588ILz1i+HeoTtMJVRV1n
eFYzIFdbvS9cAIZtPYmFdcCji4X6Hg3stgybx4BdQlprHSESregBo8kJ7iE+ktYbHe6RETHYO1YR
ueINRyWq+De+1PoAVGLQMAy7nh2HJZ9OvoAlta/RjPQ0cm/oPN1kU5KKnP4CeQ7TBRT4YuErz438
LqSSc1pluOeKlKvQ8uP6Y6A2+O9Y0HiJB+1v/qA91+BJ9zyL1zx1HVP7pfz5QTZ1dyPcjsX6jhvQ
9IFBddJTEn5HzydpXWM3FRaglibDk3crJeQmSL3HtmtyRSEa7PgiGCsYb3iGvyHZ7apLVF0X+xk2
gB6rGVW6YRqTJPOjNauIeax8YGnaAlbgGBsJ32OTdfN8LWWfgtUGo/6zD7Yx2NG5Nihbn4Ngq+qg
Kk3p1FzvaTFp78kd+12tQZjWKTPvmgDX2eYa537M03qtyqqZHzfpS/2nlVoQwUXXbin1aKD/ELPe
ynzqhWOGmbU0VwInH619h5mfQxuKtCrxXUwSfSBuj3Vp1VrbEdZEOCRFGQKEtKd6P0SptTctUqpG
ovunHXPWOlE1nkn2We8K3+wrlTzxat0VoDpNQvHjiIvpkcdo3h5p1X0DjDQEj65HPsDsIHOtM1Q7
zhyq2ALS+J3jiabNMqB+XkEYlOw9KqnA03h2zaob+L2AP8nAdN3xV0HAkghDQPeLzkCyaITzve3W
uuKkNjFJ8myOGbrI2UND62F0pqY9wS1MaAaFS5+G3NU2ZzRqXrCWbNthE3eN6d4JLCyB2eYPHNLA
4u3A+thTxZP19ZNax1++v1laDeqNsjt9iMquhifskb2xttpkxKh+VVCwsccfkD3Jh2Y/hSKL1B9U
1fk6GurGWheNBoQTevp3bcVdVOIQszkRJYiYcd8GDH1YfUSquPbVhuZkr6sXjjnfssOFgpvMMwSJ
IyZBtDfEuy4UXAGgIBy+v3no3LzqHdbrfCHB7oD1BmiVURFh/tz5I5TI8euzjZ5WGAncc7heLvgW
B25PGDvauIvbvT5qb0nlp1xNpN7a299j6bfmVWq7wic3VqHcCb5xNEqUuJc9a2u6CnrAmvFQ+d6f
3qf2umQjK+zvI3SaOardd3XxleS9CHWFG9aMmVKcPihC1WIJXdQKRbRXEO1KKc7/aJSJ94KFRjW2
j9qw135gBa2DDq0uca3Zzu8z0vAYNgm0xgnffL6wHjy15c9avsWigcrh2Hi5EboRbtFLnsXb2crY
ghmBLb7K4NKjHcd4o568Mn7Z+V9cSW97dGeO+AmtyoXcMgmf8yyIS/b7uGAeljqDAcYkBcTC0K/V
4Md7R1PAU5y3k6K46ZM/n12XzXPkqaB4ynIw8sFLMR+ddMqDCV5RgiWwnUCzSWAmHtDqBR/f93Rr
t081KtlKMwbx2f6Vf9GGerL643nFzs3w7ukiz0xV/Rxof54thJbLkMLOWfE7yJjo6TFg6C2OhJTd
7gy7Qjoe+Lkk1dvMADqrG4nAvV7xFY23V6bE3h3Qyq/CliV9buTr0HUmZN+ahz0XlLam4a+d8lVW
lsD79JGhNd7h3iDEUDbvLDpMQ4N6nbRUb+ttwZaIp4i/S30CWJI4+XBdcjrWVQssX3C0q7pvTNnT
jCpYNR6Icn6V9Yeir81YQI6tBIWlesg2A2TP2Qlo06++dIudJ+69uvwdW5mwk8Y3wEqzZYRwtdRg
ESXRb9nE4MrFRyXtWeLVp7DjGynrbSO4xgqqFRvWZ+AyOFsQXmpuG33QTvMIDZAAl3xh2Lpfzh1p
+TK+mwOOWJep5DwumkkFIy62mhD3IrGvK5Cr1xR42mdGxEAGREJh7P/zq91eAw6rVEUZb8p7na1t
MNFqmAgm0DQCqOrlsRGXFD2mkNzGNoF+bkISjtwqY8BANXTKIhoM33VplNyYuAxVR5XgNwZXDs2M
1krHs+WP2lY8ImxUIp8IINYoA46tNmV10zscK3IXOPOpeGhFVWaWuZ0abVVq57mYGXVYEo+e42Bl
71deDraV/1Gsc0W+ZoCfpAUT/zH4aVBbp1MIfR/5fTlT7rLSlOicdcTVsM51d8vsXm6ouRzDBFk7
wZhRvFg1DHHiGNYmLf8NxSigTjmeyYfRIKMVsNNCmgQJDXNKgBOIFY9+yHKgP4KC0c/nzFYqrJE1
yXzIqbSzy7Vt7jakkHgYAnQZLGoSihvFPLCtYD1BpZMKMpAlxZQc+9mcx+0i41wmh40ve4exVsiz
BssNt4FetIReEOaoooBSjTCuV5YtKRPFf2QFDVhPqApePaFl3b4gYQXS/JpkIfQIBScfozyIoeD6
yuTH/s0ubj+FTNwwOULvFhDJkXAZPizkq0ZkXTeGo5X4Ca4SSQ8aSwZBFFwicb8/hbr2Tz0rWdu/
GCnJSXJx5by8LTFZ6SCPtB6MDPaE9J0lHe0neekMQcBqy1BAAFRVu0VLGqMiWOEF0gCwWRxuBOxh
L7eUa+wBrpnal2fJuGabv6DK9WSq54OT9fis2DCgIbYd40tBEO95q/F2Pji5JP+QqQeSUN96wtSy
BW94QQZpvvVeZ0a2xUmTm1F3pt3oMLzTjFwDU/r/r8LN99phTyWXCLMSldlyoAAmIqzWZTe3B6RB
Jo/krQKf5jE+0o/A3+lpeLSs090oAtIWvw38e2Y/XJOuw8SNcTDu/Zf+qEmuQrDuWfDlXf4M5mPw
UcMbdAgI1XJ/tmjgCDMMDZzGFrwfa4Tsq+bhh7H/FPBALYSlWWe7PWy6wmn+k8bkf9ZPK2TOETfQ
fk6KFQ4ImjqKO8W+mcrkEpi2irxOsXIEEYknXcc+MPmtPkmAAOHsoexi2fIJHocIugTQMn4WX3/4
vumib4XE8XgRcbpX1Pqq2iogWi1/6jZKYTeE/PMBOtWFMDemFRtRBnI1GeoVcwi4kIxw5HRtMlpF
raDWDtC117c4bliph0E0OjCbpkhCOM1iWXeKkxNjG9RYfGcJTTWuJBPBgja+G8Eoid4M3D8TtMf/
VJ0HQqfD134DbtPXefjZLoJ3xUhOZ4i2NEfeDaXSH7lg2S4tLx++ECREvxI3YnBjcIVkoztuI4bR
8gc2KcF1DeMuionzfsMCh89jLjNYpGiGXbeZBg9MLMr/Z3DE27HsNQ6jYsqcThv561KAFBkMUEHb
Geyl1T9V1NKwX4zi2LWLSEPY1gJkRx0iQdGnWLteUOjLxOyLIQgmqHVSJ5Ofz3x5jeNixWX5MJtl
PpjnMn1PxSFZwhak1KbWJ+rl0D1KDTUEv80FaQmhIQ42yhIvHAQnmgnrYjfyFt0RMUuVR+tlUbRO
lnWkRjDElh88ccox+O1rs5iNCNf78NQK1yEqYyBciNx94i2HmgTIfBohTQcg/thXS409mbs5C8V0
LnovwMzD8ynTtkIb3hKHueg7g7ciy2pb1X4d3/xjbdmgqP2putzbALVppJm5biq0KRwK+2ov/v6z
VAoF12mtAPfUTUPC90J8Q5g7P+LGHxBNMwiBfPgN7aHIPVz6EvAMehGN+jT3731ObpSFx1oLZ7uH
ITyFw13J5BaJR7s8vW42n0hQLHzxSZuoWX9eQu7ltKlV4kZyH8cyAEOAWwL5xJ580a7XPUpmoNPF
3aZRi5YOXTMKZey/ngjRU0WS052dgRFVQQ6j0Bz4HIQ62PKWIPl08I8ZPhEbv3eQ1pkxM/RmvnB2
e6CxdG6hYbGzav0p7fjTAx/Sv3RbxcNncNVTgypb7ztORGKdL8GItmOPajX7WG9Q26M+kTyaFqpx
6uJC5aPiqDLDIdVv6QYSnExi8c67T9bl4TTudk6RVXAqEKcusL1VAYzW+Qg6pqk9oc4CwPx6qypX
8qdSwfmhVu+nDxGgihSkuVpCVYLKinwSO4t+Q91N9JhSvhw/DdNyZ+RBkoIlTchZ0eN/L1R7WLsf
qAtUZFeoPaTnQ3LqGh06M+57jpXj4pz1HTLISLvN1aPAgQqX5qgBHW55zmvM2jYFYg3kLDgLbjrX
UoXTM0zcyK8oT3yIlLrCakJJG0WnaJOjCzlA8WIsP8qoOJUC57008/VWF96GuZpZPbWkqBrFHswi
xwZYjSr8AxofdQ2R0Yk3AUw6ZhjVifNuNXHA45NS4/e40OG5brtDjLDvnvo/hufTbVfbR1Wi3d/z
BvOWTQER5wmUHNmvNRudOUUdOOIOAS89bFqES0E/24URfG3FgBbBA/v1GXCWbb9m6JHD8RAojxW5
FkC2n7iaM0OfmNHaYKi5hZtAHYym5A8VafCdHsxm0VQu5eq2TiWz7nLKBisXrog5urHhEzGMmOwU
iRqPXVLNMff2+Rse9G5Eu3ELpeTodbhWT8OunoKb9CKTjcgaONv1roy+uNAht86+xNk3NNwYjRJg
oY/ztYgplL+5N15/hul2HawtyQhRwmhgRitX3VdfadR9bLWIQ3iY09ctjxX+zZmuU1lOeCQ+ydaS
Cwxf15aJo1pSRC2o0dXGWb7hM9fXeq2vQiP4SbM5hF/OgO9+MmLn6BwmTrb3SsRedOrj+zBZvm1G
ZIPxU3/7yN8pEDR+1w3JpwcXL9lGoCST96qUCKX1CiwbnD10WB3PoWah71fRsQrY6nTIL1rqpUIP
RBe4aUrlhd15mQ+1I1O4fYaWtMp6FunGZkHrP1yIewR2LetX9oaxUdLg6Ls50Y8Fx4/osHBL5amQ
8vQux+9tmvwB4Sfv1VZsv5+yonlxbv1ZnDMdu2iHO55mjFHXCcXWc32dpdtqjG1ZiTMWUzLXsVgI
Ds3g8ZxmS2bW5La0a8wEyIzIoUtjm/stWZE1Zc+5qbzPhKOXV5FKpE/fAVuw+H5c37pl9UlSpFNi
6Z5rp/swNqcx06sMwM93qUC87wDXtb1uISU5J79X5JUA5KJ0rk07GiPDekzgrNlEanB1+qNhbtZq
R7H+Kyrxjm32o4KNdqfvR/T5vOh0bBSOcGCwzdVTILAQ3s6Xh/GyPmqDTKSADNKBG42Fg45izbl2
QzPgNwZ6j/ysbWHsKpYwGzPNMKQZXNGiN3kYTjGbrhW7zDMleYXvS9Q0g3G1ihlf8hywtj3axYN9
I5CZ90a8vmfP+eXI5BbGDKrrHxNI4wv9xqNwYBBg3CZx2ct/948lqLkI7lAnbTzVts938rZ6aSbH
L+ULn5r2JNBXn+YxV9Eqe6lYw9I5bL9xRAVyhN8q6HNnEonh/d8JWzK9UUSafFm9Lb06j7GeP7bT
Bax1Y1K2v6zhf0SZExKUpbOPG7Gox/rzJ8/FJgEJrtA83urntXCgIAmjWAoQ7zi5nNuw9WvrCFB7
0c+JFLhgWqMkijF82KhuZWK7IRpJ4EPJSYIf1H3tzCqqUuuCO3yqSS1aXqNK88k0Z0Rj/Gi/8XFM
D6GG/AqMgB2pBT711iw7dwVgc6KCvV1y2oTyiZ1o2RB2SLCU1p9gkkk839fFhgPGgK0gpx4fGn0Y
xbplb0564grkknIVUTG10HOPEEV7mk/lceskvyCTWsB/EUr1BZqIwmV9+VyY9ZZsbrObMe3KQKuD
VrZp202F52cbZ06uu9Tao1eq7djrrVxJxUDSPZ7bDZi5Acs+a+q5NglhRqkfzSVSNAxyrOBO8eX5
VpzDMVEGO0I3aBRpFXe5EuhyxmBWL3cTWkEQyLgFjw/uPQrKscYlu7oz6Yi35vekzvaK7l//QgfV
jOK7soQ3WxtVqn8CikcYJvUwQnfDIx/RR56ZGDRFdv2pH0pCObWe6k62s5rL/XhnR5KJ395Y89Gu
dOlPl/eylWiWB+q/Fg5JRCeheZn7SXtAb9qHrsyY8AQKer0nfV7+qkvgdqW5RUEHtSJD51nubN0O
6S5enCEzSYL1vyzYif5Iwy6mMp8BlGUfUVwxFO1T7HdTH358Jpw/oMbDg+SoO1jSZswuYL2HcYEe
PZR9Ujiau6p6nTxoVsmgoDrhRetyEUSDfM+acVo5lgAY6IDHE6evbOFZJmEUP8Z+RndKmaaHDMSl
uFTBR0h1QZ/AV2TVf4+W3aHx5be9l7Hq2R3I1aqINGkSiouH+s2+ZgkxDnqkxJv6h2wnRuumb3w2
YfnwJMPy50JGc63XCL+tZE0Qe0QWteNtSPP7V2fKrw6xMDf4VWJTko0hMTnvA5eOJX3N1xnhs2i0
JjIhf1cDataUhBx6cfeQebIFLif79co124RYGPeiCQr+Y2pYxsLJhtO4HontKSJ/IpeQh9NKOQiv
FhwywUsBhFXp/6Tqbf8456kiV86Tt5xBv+divn0x59gazgGzclnIh9DNFHjxaKzLSSd1sIQ2mTC9
4hqu1EUpYWT9nD5TmzQEoap57TGhjCvdWYK+lmWcDk8FY1CFOm82wRZmOdZ25VMpJTNX9yRVJ+As
grJvSv9LZV+yFoKFKC/qBH28/6YCEhKUz/6uk0/JwTw3hJ9NbZ7Yfxul9OVj4vv8/nCTCfLXK5jp
1B36neA/obgEFya8H/L6F7MMcjNYYEvPFWt0O+6Odrd0bN7DnliJmWEtHqW2oT9MwEz0zglbNbkn
MRxpeAa0nQ/oBkPs7GxNzfYDYfLpjLOB+ViJ0de7BENm2o2Z6aDOHbYl0fe5LZvwjH8BM6Ikqjsr
1rQw9pAxVOVopPr6tUs05Bu2J0BLXVWeeKHPngi6nPZwIW/k/kx0xy3fpQY1tPPQASw9mgIRJNRw
bN15EwquQ3vC3NXQe7yuLQH49P9OXOVza8l4iUTdGJEO7OMbulup5EAzkz/o9Jr6qhOmoe9LiM3c
xlvY971Qab+NLSJN1p/jqUfd4J7Yoi3QHojzfeb6HvSKkx132MmyANizysJtP0yvUUzjzXeA7fy/
leGzbGPy8/AJcnCvLtt1otTy192Z9H81lB4Xwoy5E2Crt69ANVC56qvvB5tAlF6rW5xWbkorMO9j
kI5mOpjXM5DzRybru1CAubdrneAUYhWuiZbkX4ThDcczadUYJSzJqt8jVy3egvjUS46nQQIyQpkl
nsEkV81Nq/CYsNXhdK6LC87cN9su68Z7j/9vG6zIuYVC/QgTmSjydfdrhZHQ0nonGwzNwzaSNm5+
DVEXDw9GfIWCyHHHfL2g6OqOjthaeA0B5ge9CPJcKpGyVttzegcwNmztHPnVR4ApNfPxkjAZ/5vm
x5UxBcHAWigqvijHY8aePLAVmMVOVXl6hKy0/FPMv5alWpTNGAaldBPDA7ehvZdwh2v7KmToZ9+h
1TX7aaR9bZd6RIKkIg6qd8XJQGhyuHemyfYsSJsncBSamaqEvZaml+uYKSP415yf2ZIy1dhW6Bf+
KBe81G/W03SbQklbL98rn4v1e9N8mVuNH5XZmY/sgN8bSgoJ9dvmEsq3GhZbG5bDj1Fp5hkL3XZK
dA91TO/P+5WjJG+bXuNlejQ2pk4kccrg5QS85238AKDfW0gIh5MmAde7hdnYuH/CnKLj5ZWu8sbx
ZO/wh+iCLHNPA0qu//so0hmsiSiMUuJYa3h2m2Gv4mts4nRkD8C5Cfpr9pDqC+k+ceQt0+hODZ8s
4O56cTTSPAHgQBWNYKjF6GotypJh54tBrf2krDiYiutYLQ1Ksd0dLaxogczOa1Nf+NkpgoKW9EsL
PVhP43Sc0zmYY1fZdHceGvTXwwU/CeCyI99Xrfbny+QSpGJ/1RxHzT0sKEkrz98+wMmYbAQav60P
zh/BT8ZAS1g2zujbOgc7huegRaEVbce3QONLiS80DhdpWPATWB6y+/Ui3WwaNIzw4PALwVcxkDH9
fQ6HnSlg3oJPT0TTcI72cYoM97PYmzQbQaDH91h000Cd/XGC3lEDHX5ufpTPgOq//O6y5LMuK9FG
EpOouxTrpftGGopJm43ZKQSD/f3+J6r4C1oAn2n+uCjUuxNgObjkHZyRxbuJyDzICon//5izVE6O
XCDSppUjz0CnwkSn+5mCocY2y/mz+wGgC5X1a8dYwyJo69kRryeJpFuG+MxEHUhG1u+aA5nqKXOi
KlkxTVUjacSI91zxX7hM5RU7SwX41DOsc9PyRcKh2LBejS5QsYDtguSgEnElQSOtydbu3bn/DlY6
Ly0hEhX0AB0rFCbvDilov9bOGjIAOIsRVJB5SBDpXTo81fMgGUkN7L4vpr0Rxfi8tvUQHzmBGAHT
MYQc4sOOC6tTYmKxChNn6iuLCCDdgSh4BlwsGEl7MzH7Qpmq+gxRS7y0nKZ182x67hlNrM7h1CG/
9wSrII1T/2+7cYmHTtfUVSPApY3DVQse8kXElUpozXdIR1A9bXQeqNE4IkSJuGobB/+1cJonTCA+
q9gZI/O4LmWTJSBqQG4z13rLcnfXpK+3OUA5/DlE4FG3rOAoluhhX79BESSkiFz3AgrRh7XXU8XW
VzuIYrC8aKu+u/YHrt8zLXhGW7NsB8ZnDFJ6g3TQAyoRE7/r+PxMSkCvRnn3KlFTcP39kHeN06QV
xMPW1O5yXxN063EEJsfl/AShnniGmomG9+aRF2kDRDj5iBP+e3onN2jnrBuBmuWFjA3tsWTx+h3G
eHoQCbHUa8f00slsm0pBVDuo3KOeBXDJvnEK0VLgpaVPVcTgLJIWlWiYDM6IspHDEezuRikibNS1
QzN+5k3T1tHwOwtCb3xpCt/MBfkQvk+Ie2Nn9xiK7L5JDtNzORQ2tcWX71oR0Uqx+jK6Gjq7T6Wd
5JQ0Kcvb81JE/9D2XPZFkrlKAKWBPV8EXoGAaWbL2JnOYBBqJZEKTvQxTGGFYkMDVdRdYMQeXUW9
cixRkFP8FqRzfqF8Pcc8EPO5ZoYSOmJgZCW77y/8KozBNtgKsDuL2QvXMAJRpJTZD2duFftPl1RD
7GdMOe4AkHSCuti190x/fNTVGKi1vVVupInGQeXuy2LLV0NX9VTBUAEja7rQqKI2JmNPqgTG4QoL
2p8rqC7uEsZ1pK1w3EstKKwL+jvFJIemLW6FfS2fGI2wP9uCwmdfPg4HxOYkwTNiOsaBE1qSrAWo
wl01kwu9RlTVF0b0Idcvut7dKUUqV61mAEVXBdGFHpz1RQ0HZbFW9DyCu0JM7jRiY133Fq4wsZ7w
B95QpVMBW/6QhaklMN9ujGmaHVF9nYxltR73Q4vE+cT9btDkuqBseWLKyIZdDJKBO+Uyecs3+QLH
pRrbEtODcVQpvyquljjeg2k6CJBUQ7ygCC8DQHf3EDm3LmrRwXFJoKyuPD6AWrxDbG5yWrpR+DxG
h0rt4MeWShYk6wgHsjgDUBaNwuPiw3gmu75snTprNgaVIOXzwRZfMfK9/IoGYz/TJpzN8HmpP7jl
bB5MZWlvuA6Qeza+LIGCWXyTBG2u9HmW6ufBsOcp0V2jCF+sFTg3nOsBtjH+/HgQnnu6h9FkPqjg
5A0keEziJDPXTj6v7bUkhS4pMaM3Wzz5YsArnVekpR6QsmWiYE4fTs8euWQ2Chog8/K2ZTvNW+YZ
WGPBzAn/LQzyPS1DNyKj2wPhrMhYaYnvjjHEVivjPXFtfrVC0NEQFNcxL5BZMoRxIptu2wymNrZa
qyYLXMyN7IyBM2hAYh9sWBzcoUW0rmnLGF1mVDCQ/35PlMIe3f2CNLdYriHXsg27KL/PhbSgJjBv
NTNbMvSJE1MsdXpiq/qWbQLIDr6gewopUIP+bReCzBEk0wN/VDXo+5RQ5sS2UoVArZZGAbGYsKcp
ZEkYbTePhYHtgtPhaiq6fnNKT+6pE+CMMy76OcU9a4qifrF1/NALuu5OutvBPsMeaOI6tPgYd0bL
ctdtheHpunTS26psEoaK2lIB1D2DQ9bXZVR0rIykH7DpPxaQ17kFwrHupkRkXcOPCizJhAz3Tr+T
202UoOheydn+okDmldjN5fSyemPs5vxxZkFCw2EubQHjfWSrbimtx+9KDIDjjLQRe9cFX+ZId3Oo
95iMpzR0UrZRB+ycWz1sKoPtt5r5NhjN0fLueCYj2O0uhGsUoOD/5XhK98+4U8UAHZ1Wgx6tQNaK
gRlrNsZR04akgfDQglzZzmMAEpBY9t+8UHXy4bMtnngNdnJuXixPdLEiQ/8TmcbCqarJvXdTqzum
/yMD8vy3LSasPNDpFAKZ43Gnx8+v6Nd/gsfYoTPgTxaVLIPAcFDPsduZKgNnxCufDuc6i4suM0Eg
pynjG0nswcLDeX3ihwf1gpiCH90byJbHcjINwu2KD00S1LS4/x14mnEwy2ae7OnLTxZdrsvIlk6c
xsIucnW5s6MFvYcaeYkAP/WvKFNYFDGlJqbk2loLAi+CB2bxNiFJdXIulU5CfQ1x+PmpmeJbvTPX
EtZ6oC2E7IZl6kUKBauLI6PupEu4wkR0lVJgKRNI3DFsNyzSlAtBj671k3gG8OBpxbHv5nb/Bc4b
x5vA6K0qn+0p3SgGyFIy0c4G1CY/giadzfMgj63MRxIUKSbWaBeleKMmFez8gOJZT/kquH/L9nqY
ii9yHpiazItzUzA07kleE29xm2xZUWYuI5Cd8UDya6MsyYwBOw0zy9m6MzkPYKw16VNxAi2Nl8Dk
qBAJk+FnScKKLyWCJ9ageG4o/OfQOZm8AqdmCaUX+8bGQzwAgsjPDpRT5JmHuxuA7/fxR7K6vLaB
ES4U3+Br1HXl3K5pJGzOBacvo59r3L5yDjuRDig01DyjavM8x9oAYXVAC/KKz7CBCFT2Pmxib9Zn
XiLm8VrFNOBibDchs+Mx9Q1bv8Wh70zNqAJBB0SoMUR5GcUvlhRicyfmUjZLiUSh6eLb7nM/uTZW
J+BgXjb3B/mEx5o6dt1sXBeWlemGtGxykJ4s7MJQ7hQ0lr7z409ilPtUTUEs/09PY3lAJbA9sQgk
MyP4gnNqt/kiQqclxG9uNeeGoLulO59+RpjsEIxdFQgqOWa+xzWK/L7qu2znvmZUstqpgYWj2ib4
zQi3Jw16HEriWpFLp+R4MUTp4RXvmh7g/7SQYWpDkyxTmwkPQPewEFMhVoqiPbU2RFJ51vbI0uQE
BRBW+1kf4Qoq3Zw2pkWVPpDB0VSGw09wP8xYNBJaj43OgwPgZSbvvRl7RE2Zn0guqtKlA6lanUCZ
NEnYHalejgzu6O6qniThTIWO6n4ho4+szEu4d41LZkNnDkDRi9DWcek+8a7NdJR++qb/S7xgjNdo
sTpiItCG/TySkbbnrZi+m25WpRaEJiDf1elChsrOZl2COkd1rKq0FuRUF1FRMCLLYxYGAxBOyVl6
ZgloK6VTivm7WIph+V6SqUArQxqLY9Dou3My8SuS+DuDH7TxZA78p8DBpCZDilg7CZrrgxEIyfv5
gE0Ue/kFG04fAZPssjt/AINULsd3OhLo76w3FTDNmOPdEqLCao1vulCijgrqfJt4J8zeclU5t2Qk
SeIuw0sG7mjRiWWz3ce4U+h/H2gVl0NUo3RNojOMMzc9Y0Bk0u4ntWG/Zv8MNL2GpImPdX+kaMzC
y3wUa+SClnng2SwY4YAmlh/LLAXi3NNYhfgiGnyXUcJpGNPDBXi+RG801V7fj6euAt9HU0Ul/9S+
+zaZ/svYbn/idPNpvI/D9w0i9fo+M2+eqnOcvZUSlzN0DxrpLV3RCORlyeRE+1BW1EsAl5uaAz0r
ng14U3WAtF5YVOdit8v7wzeGkcNSHbLhZQ73g6Z3rWx47/7BNKwhLQOaMyzEdUk5FOBnHm//AC65
6mNABlX2nF7IbhWw6OC+k2MdPatNvbGYW80Co581GEQ4AOJ5Fp8bmwnwqzGq2xBA/ngztwHviXk6
WCd9og0ioNnDdDI2OH0zcXRgl6g1uoKFDQr7lDcX8pyBc642733F0evvapodqZCzxgO28XWic3CE
MahjSdIdIpsxF6s2ocs69HhIEF2eXe4f6Cc7YXKjNRXY1K70m1JlxR2bpuco1YejWrbvq7f/Ritx
tW0YTHbaiJALXM31S1gQ07OGN+qAZbJs7Q770N52REFpYqel68uwYd86MuRoeChmlnOFm8Rwgr6i
hUE8y9zOgZOVt1H8mUt7qiX8FJpIOKBn0Xk7XjuJrP5cyHNNeVQKZHfGRmWkR9xhEWy86sBpYCsl
P1I8zeGBA3skVknux1WQGR3C8AKsbAVzPHQ4bLd/egJiTlDrX47CRI4Qzw3PLXJHRon92QuofmmR
nx5jb5glm/gekX4XMdCSpZqttXDAk3QoTWHPMd2ENbjMwmI0Oh8O0jTfPQibwHCVqwQaCx65VYmU
q6trct0RAkdsczxbb7684ZW0O4keyoqQpVWYgwWHRov1RWNerga+4LdlvgpBAJ4qCzJMrb1QhrrH
wQpIJBGNT/WJ9QGFD/4AfHE5BUsZvwKEoub24dezbqFxTqyBy8tq+wsFVWO3SrdLjVmWiO+v/qRP
yoef7cdnOeD1E54UcYTleZOH2obA3m+94i5pSiGyT9tpgoi3F1zbyHYzDKJGHqgkP7U2BK+NEjs1
HxQW/m6UJfb0RKVyhSVRJbxuESyqrG+Uy5VwH/wy4w5SfbAxs+YhJ552OcVP1A4FCZnGNEia4hLA
nm/gCerluJPZ30/Vj2JTdvwSZsmKqwp8UkZ27qT4sDO6WjgfmtI09Gfy/CcPhEtA9obXgb9iOl0+
VhzKd1LUktndaRXOi4Box1puQjpkfH3w7xeZgkG9J2XN/KmQq6r87+1giQYSXVzn5RTZmzANQIqt
xZzrI/PaWBgLvVqSHXhCsF/hDDXrXJwqyjg9eDoLfjLOvPs4Z2uOxdMYXmM+c6ys3VDZilDzUyk+
QEPI4ZNDZjy/sOUebBXgv5N/UCve++ZzOkjTCTQ/jj3pABiZ4TGa2GTYzCxYqG/WTspA9OZKy2Bk
dW6SEZonY3DS2QnihZehoU9qCTpwQIDC9iDPN8AREtGyUs0kQwHWNSTh0dBn0bUvH2waDXpFGPxH
GPgEPYWVbdwA1CETdBoVyvqpynjeBGdsjVB2jIr5Pe+ZLe3g0ibcoWfBLQysxWd5FEldEkjQdNsV
lAP7LB28E7KmhXCmnElOZT48qy8yQ4eC8xwdzoBVZOJWuqbZTS+zNaiQbJ2mpkATxnuwKylRWtmd
TR4dPjN/g02iiDYPTa3jWe3i+7sarQKU8gFiMAoIi5DLbkGTO3BC5M2pYTdCvaankP3WAcYqu4jq
Ed2g7fAxXhSKX3lDqtoipYsR7KYPBULGctjruAUk6gGNOvjYHNYtQprfOjA5bhFYj6wXGLuW9VZ7
k+8VkjgE9xRO4GZ36e67xgKGG75znvnjYXBOdKQYUKwiF/69Wvv6CwiE6WuRfHQvMb4VGLleAIeI
kcCuVxl2nWt7d28iCvBJbdA+O93B0zUcaKco2sYhiumllluc8O1uoQlOOJ1kC/JfQ8zmpDS+i8Iu
41DcpAd8hjqSyKIIULKVnTtjBzGVK5rLF6lmfkAJV1neTAU4zxr7XQa1sloQB0QuF1pF/MD8UffI
33bzRs0DqlDuoCZDaZPgOuFMP0ZvN3azzsAkP11mDwAEzJ6nAfSRJysO5F3aBr8qKTLmgvZYpGzy
flQqkviJmwup+0g+emPZHq685sKdWVErR0+wFODWCJHWuWnYqwK8JdLiLtqoBA7JjJQaQivXmBIE
HBfBs0iu/mm/6/zQMxO89gCTmvh26EhstBfEwjgMwcWe2gwCdwFMTgoUPx1uJY7sZNs3IS6z+jHZ
fMWZqTZtmxPFrmOt8Y8S4CMXvA2SF6Kj3txHtoW8smqs3gUX3m8BtVoyA21Xmy9vuiiftXjtCD8W
jWIJ+rovcB/BRGj9KACWXoBMrDkNlJWHace3v25BERSuy8hfao0cWOvpIZ2rFOOotPNK4hp6FNY7
9OyvHqkg4IXhCx+7b3ufPiCAhbgigz+eKlR+YgyRA9tGnM6i3mXcmnieVZwapE/Yijp2fLq01O7a
mPtrEsqyY3M8Wt7g2dIMWebQxQ+bUd7vOpDPpOvE+C5ScAQdzx8RUIUHt2A99D0hVqqMfrdXppqi
wtK5JCN06nNsULV3AAh6EAjPkn8qbZeR7zKbDSv0hGwdqlcfcQLNV/XLmtjjWtAgNGExB61pZR09
+P1mnYlv0YJ8didI35tGbRs6jYCayIHK23cl4LKtc3+FGY9hC8ORCns9XGo4TXAkWMwNEnbQh6wo
0s7OnIv9ISJgAGKcTdW+F+NJ2IBnaPuCbomzaB1gYA5Wq3oJp7GvemINGTzQzaJTXRZXF3ajOts6
Dm75ozX5gQs/l2gRlqEze4iZIiCVoQfy8CWL2yZly+4gxUZczj55JoE5Rc4rhIHPhMox+M9No4Zg
HGyX5HT+anDDvAGceuyV76FyqL7Xci5qD4gunEao+iHYbx5wl21pwBaQgt6vuoXoOu71SJgtxnp0
cXXlusHp1Kg28gSPwzbrD/b8CajhVivnQUbl/b3LJKZjOPNvbVKaVjhHJtysCXC3rg/IJUA1pw6z
298pcK3+9eR+p9Hw75Lp34GyNdC/1lDs4/J4EZlRP/YAknoQdDEOnnBKSkCB5PStxwwzabSSKIrE
bepPkvQvl2WfSv2TrvNEdGfGad0KfRGEN63JosXsEEfqJ+Jw/sDxirlApRM8Em09hmdPUWL8xsTH
ZaGVFHlMY1qgn1naJ+QUb8Y6AEU6ArGhC8xbJIOhiwA47D4X0CLz5nzjEcWzIx33TDEy+Kms8NAA
NC4mUEhvtoXCJ3P5ksXdloUcX9lHeRIsIB6jkeQiV9rwtj8g/RlIOCoRL3IMeSigo2g0AsTadzvV
G8Gf+n37NQseYoFcmmZ4uvSAI44+6Yw5Kzp6Ba+dY4gyOpz1/oqFxZ3GKQU3SSngWJjl0H9xpluJ
CjlCVot1xMyBoEyfMPbiRl4P4ez+eytmERCuyITecZ+j0WHwFmC1C4xYVsOaujbLpcHR2I5OGuqF
SOitK+TBZLYb9wJAcQCIkPj07H/406FAx0ZFyQWhbKUCJe/tpSbPxcLdwhU+zr47qQ+1NMum5ryV
GiRBKqa4dPkINjPxwjDCS3PfZyxQ8qJb0mrMtTtN3jItFvhspcSvvsCZHRNIpNiWrHq4ALSU8O5I
IllQJLHqtXaXdA0yrUQtYSxIZldH1iIVN11mQuB85jcTPQMj8diRJHiLWPLb3Wo8QqoHr9f1qeHV
fsj8ynfteW/2J49fhA8DH3wpLx6pdH+YtyGu8FqEOXfqrHC7riupCvRFVSuamU/uQOCbP3TmvRLL
EBVb6ioAkE1CG/ZiGHWR0KXzb+KQomFwmLV8DU5yhqtRefdOWxlZuyErfG/Z2o330dSQd5Y/Avsv
6QwsK3iD5b1H+mEM5CocoPXjPy3SsW/yHxij9vrqu9saKqrDdrY1fWLufsTHo9bvWox37RmAMBa6
Rjh06Z3xr3l1pUUEcfFvNBkXMhmie8oG8Zv/GHujzds1tF/s6xD5tMCgR0Wbof+soMhGAu/ZeXDq
5UtUxdIVmCGvtdk3TN101nbxgfc5VN0xU9KEV2lYPJehoDHruFPLOLJYrLmFfI3uzLDwP7voyNT9
CfLUJ6dyzDS52XFuflM5WHrnN0vkZQPr6Ep5ZEf3lIHWFhUt6FHSi1TmSwsO+kH3+YTndrk+YTQP
vzEbVORWSjfHkH1d3HvmDpyrYEgTByAJOAPbEitXjtZqbgqsd0tp/fXpcoDSRdrolQfJ3u3P0Cmr
Y55NzUDruV4sghup0FPvZ58QJjNcoR1VgU//ClgA7lXZHW10i0AfGtC0MxFKAHGkfs0JvmA7ZWBl
T2qMQ6RXGRa9nOcJiNS678+Ykhp0pJE22baxSLdc8Py52he8gXcMCgNrZ2/xrLwiXJcdbYnM790e
Q7alP65nR1THl39xTJizgCkOSxKZHWhYtv78cHK61GoLR0xpTRefDtEkj8o+5SAPT7LnHFevBQNT
6DMubykKjfU5CRagvSW7hVhnbVGk5npF1GhTNcMOfcKUkgdMqDRT2OsbCTUjf4IUULrZdkM0VUfm
MFcHg1WNHehEUjL1c8hHy6Dm5AIqc/mRCYc1YIUvHWYZ8lpki+nT6zPWfc48SZ7o6iOo4IPmtL8H
m1RHhdzi5lQQFxGzGSU0zoMFxfcr4xMmjpwWGHoWzCzpYV9m+GxMGjmAUKp14ySNR5NvPcvk7PRb
q/bWd1rsWDwt5QWF3+ORu6XVNd99If8oaaAsCkd5yjMyKm+k/zHPl4PaV+DZqt7LoR9tIdqfA0vn
ViPkptOgM09MLFYPms7uTrhqfIH1m1kjW0XXKFgB5LBTmYrDjhPapvqWexcY9YiW0DYRq9ku3RpO
9upKMyPW9sLVZoDirU1v2lBKVUeF2YvMCy8gQcHv23i4PFplpZyjF2V9MsqtyqtgMKIYrTDwxOtu
/BYL90BeK2COpOFuqPN7aMS6oovQBPleKRjcsa4+nThy229Y2ggaBDW07MZa0+03gmUwc4x18v6b
Fgpja9aVnT1/w5ZAl+DxSusENX/5zEq2wGjOiZX3wsStLxPg8fSWJz+sy0ddEbnYHsIx6jh7XP8h
0Ws4eCSIKV9lv6PYoKqb6LrTBXidaIEkiU/DSTlUtAzfZcQ+/Ch4XfVoGRSh58yNJhy8xm16atXy
Vc0Gbm2Sij18siCLyHypWKb46aDCzG0JeDbuX0bTI+0sZZCZoxXhGO5Tv67aQ7pSQ8GoiRoNVPN9
NcVVV6fUK4uxENHJnEC5kHXrah44H/pMsDGQQGsaonRA+BTOj+Wewtsqq8qBYpnGnIEhui/kvTHF
tOcjUiPZBvpy4W5gtNpMEFgox9b2BE/1icxuas2TzdgAaOOxE7t7QPmi6zBDPv4zkksnJy3PhGlQ
p5ngKtC7MZm/hbtieyhSqFZ6BIyHHnsq4oKpzoEIGIbjn74QfZhPhQvgdiF4MUUMbqXVEw8h4+DY
x5Bw7jB+87kdxLqfKAELBgiAJAkE2fB1GeS8CeuO28GcLyRtaeMWbKngvkOGUGEHWwkjJo4jynLj
qcP7g7hIIQei/iEVUY9dswxAuvl3RuaFysVaBKaIV8cIa3EOW0fCVXI51OMQg4ftKPtEjgKO+1FN
o19LlwOBH9n9tLRK23RpvXG88G9rKGuqLVeaNvCMkN7X1OTPfGVmS/LD6xYG6rv9tkZru2tcHO57
GzUSQxrDKmTTyAF4ufp0lIMUkgOwH+Z37tzRzKftzC1Mf8J84hhIkPc2B+iWOa55OY961BMVTWRw
kUj/P6erS2ciGPneGDdOk3S+UbI6X6qZyZ5mLLb/Ie0SniSRsXLGJhwmE2p1wprpZ383MuYN3oWc
XvshR9UklSmQ6KFxRh8NAoU6/sahbPgE4C7SYSIEqfLqrPXEWhBuKYhg6euK60rHat5gR+Trb50l
owOLB9JOrt31ltxxU/5rG24YCfJLOl7S192AMK2OTe4UIWg+xsM40DRJytwzGpDmyvt0oEpNuNH5
1SfUszH3t6kMOYjPRRhQLv5i/H9HUfImY52C+25tYxHA5fyzS2rctUkyeBi8fujPRmPee+NXuQCZ
fbw+ZWIV/a2pX4Hf+Ibk1+MNQghwqMNiMHdzwAptZLlPOfAlsgcZjysC0/bymGJ2JM3/hE5fbUqY
Ha4eWe4v9ydIsV1Fqs0YxjYDh528IHm2036NY7hj2BQSHY2l9rAPKMS4/BxChCN8AQcecBTn6oB0
abDpBmQWs2Wj+C5qzskSw8GyxwCA2yDCMSzZSfp3ohiDEnwZmLrEulDEcLnyLuUw+ACMJ373zPjs
LQqt8wqBOp2zjb9mirl13JDqGWpybEzsYIaNyv+gOEq67RqtlrAuu49EolF/idbjLq3rdHWV7MyC
97SIo69Oo/zm9TB7BrKMN24fm7uM8DlD9n5Qez96w8L38Y0SyrEg3/Jx4444X1X1Er5sV3X9NP31
QVB+nAc1Rl2M73HBtCBPxfCdiz4PcA+zgLF+Vr1Z6nZxTo7pKtZA+e6VF2lPbOYgMU9ivCVYDZiG
n65claCzKBAu0SqVXRPT4yYEso0pFqi6npI8NdpR0a1PHTTXGv0W61rM8B1vUc1rAyCe5UoIjksL
zWpBSLmmly32zVrholRGsqzGijPz+4oBz2inP7gyRHnZ2w90f745hH6r8TdB3gm7PkWtBih1PpVa
T7CaeWYAzyIfTvcAxks+pSP2ahaKULVp2OA92I5PctHl0Xih/E8sjouWtZPmuy3emgPwzseixWuC
EYrb4b6Yre+eiXEotKUn3X9hjByxo1prbLvc5FTatiYGlaCAybO8lUmVfoICCJ9qPP1raki0yKQM
2bVGj8hzmxcc4Xi2Z42CVgqgAPKgIHlPQlJHUJuHF5XmO1IULnD01cli9yZaMbAJ9C5GWGF9RMN5
xIvwOjVDb94nmwA7c3AO1lZ+0yIXguWSmL4cnGBT5/+xe1ZuDka7hYbmvKvUChB+sP+4vxiU7zaU
WkNkCOzZD8tcevrt3poDdpZT7DYC03zuUArKkCz5iOFuxXeEFQsrzC/AmeWrYVcM63p/9pAs5gyZ
+bDoSua/q49VcmGtIalZjMonhapDJJvJBMGnDdvvwxVvEV634QeDyznjVN5TqH9Xf4Ov95sUH3mD
gzlaJ5ycPrUEZTqgtHnxR8R4s9rwRHwcdWHtHStiWxFadMoYsdVqVDvXmw6Vv+TDujIQ7GH1RME9
M3dTzTHJ6PI97FfGVpHiIBit6v7hUpN53i7JKzO7OTImoMRghf2SEYxC5B/MdMFeKCAMvGr23Yqy
/SYMX6/7ViXdhANB9o9NOxgChZgGgWayxJaQRaP9UPyCJsHZ/ZtE+9fktX3iu40zmsCQJBKoJcSN
KvobKWkin41DsukLezLnLMtbvXtLXeMSi0zvH9DqRnlAgkWoWQOGCTSmlodToTaEhEO2Ukxbb8lP
jOA3R4m6DEyKhdme8PnRQbiaYwSpBB3376cYQz6/ag5Pl4hRE4Ha4Ac2tJN/3VCzygFx9bynPTdE
FaVoqsbsjoGFn+EJ54lLfqRJmiTwfoTdNd4HiOvO6qdGNTRX7G4uxch8SJRKgIukDilAQdF7B6PS
eEcsnkbCh8DRfzyhmx0Wc16hhFhc1c26aI0fbTtXvAEFrr1RxIRVZmuJq+eIts9lFxpwQoRTCg/Z
dnMNUjk64z5wvg8pvW9gzmZHuIuKPPoSU/BDfuNeWyiGSF9UjqfCZEWS/gNX4Zb06K3FDbKCOVQW
n57JyFhpZh5KvloI+LIHpNw6xclaFIfAfQc1878KX+We7kboii2bv6Anc1lxHHd+Fqy4MaSnZfd2
ks21zOaHzYbVgQdbbe9pywFfFwxTi0ldH0LWz8vqt098Tx95r2g3V2wDe5fQtvSVh9nmTZx0Yzt2
r/A2GerlZx8EGmaHGSmqH6kGHdWuwZpd0jZuQWRSTw9A2w/4q1NCm/CWim/YkxyXQi863NlTy/q0
QbugGJ7MCqOcylKZTiryWQn473Bp2VLzoAx/MuYYlgHuzi0k6GeDb5cNcsAJmdt4IHIhfOwLA7u1
0BPY1nqdKUDwZ0KgtTr7NwE3hW78JUQxKYFYQURDlXaz5mBCSxvCHabvciFkJ9umtSYZ/dEktGNo
eL1Eqr+2qWO5Hv9L2bZTEEspNJIJRrj8MY6yZmzCQbaZGeO/9J9WYoCdeES/bgJyizqalqxRUUOj
8spHd9UaRaIYq3sbMoC+PUI6KVNKH544yRgZ0T60YVLGScRy05AfPFvM976D640NmuV+Ua68PGT7
v3NZtojKiPdv1H3mmrvEoEMBvYI2xct7oLviuezx4hjfz24KOYwIIsatPw5V79zLHoUxsY6hnrBt
k2+TIOEcU1QeUgfGrdXlOlt54W9W5NSw9ITcC2UZV2sw/ApGc62f4A+StQr2BTLrpllEGKFPvpzi
rN9fJQlwDgvAELQ+wBqz4dCu/uJGk15Wf64UUCPAYFVkEAFfxhUjAKzXyQCS2OF6BwnQuCXuJ3be
k1uvaVsHTJ5UMz2Re3fpzuufyh8C+NanUjSNq6hiWiOTQnNjXJ9SzSNZWpTOilPwO1jNDAfe5JGv
HgysVv5hkyGiXriW8ngUua9ZwxESze/cW0CLgc/5OoLcqXjK2We7KqEVIbpcGdTVSY+OGOKpuUE0
+LyFwffYLOXyIDyXaJl6tvl/HtxqDEQwT7t4e2k9pm2mz/xip0MAKT1xX4Pl+3EHRsPrLl72mfAf
aS2vnz26fivU6umC8PHaZD/thHXvbQA60ZWXXZbOUqaIGLSDkoSVmzJCaKNyBVTMlMpRPPPjmcu1
LUh+dvFBse0/g/W/Fd6JzfQVYgvBl2HhchT1yE5uryERkctqClHNmPlaMaglmfxzgPzo53rxcOVL
Y18bH70rxfeyoW4rEhQJhVY+11XVpO+ysdRQZt9Hc3qMrjn2IS834UdmgkAXGLwjTqe2BRztp8HL
2JFRkktUsibBe7uTc/A+74ESFjCU9SwVN5xNfnipN27gwBE/FI7y5ELFmlqB79vx+yfilnH0wYaI
vvK7+jm1Wm/kR0BW0qFimHpW7PJUlr2hr/TaGWDxsmL4kldfGaRlVMAqCetkeqeuDCsQCiY0wuxU
PNWnG+zKnujCDVp1LAUMWCeTFWNdXnlEAqWpgCp8A6mOE0M9XBEov2PV9yhi4JAdH3eNtt7TLjPI
uTCKpXfYryVzX83i87X+c9IEd5Pe1muqYj5SXHk390RYJaLLqD3bRc9EoBNgoe/xJ36sr8xqME3m
l+51ihlY5ysRZnGRBlqCTsQnnMm4PgILrd8VtzkFUjFOCKmsZE7Uo4hWXIxPsVbPmJdfXZhQ3zIl
eqLST9U0Q11hlQuP0R9UqrrinS7KU1TzMZ/x/8aaB+vsc5CXpNFP9zq5ClHNG1Cs0+C5sdxYRqPq
FDvW/RGSziP6eMN9shtGCTbhA51ueri8Lp0S2JtPNZ/zga6WIy3DwAvKgneUJnuw8BQJZHrAJFni
8LmCO0yvK6sqt7Nr9tQA8VW+QI2ZPA3QqH7FXvuazQMpzfXCF014tCaBIaccz6Bn2fJrMNnJSAs8
l6+V/qExNAiOH5HhPjFjkQeZzfvI9v42sHINWVR4GYu3B92j++91ziYD85wCI7SRm+vGz6WMosxE
riCO1r+LJqlQDecH7Ir8UUYakGS4J0u23RgSbeX2MRhKwXLERR7Udyej598wfEwrZ7n4kXaKO4lU
UxzPn+XLyRrnrpiaQFMSxv09EbRx0pE4KdaczY1jknwJ+efpIL4MF/pzj+istp0cT3uu6Ou3qaTA
avrVXhk9K6vgjGA2lJ48/Ni0pLJIelyHP1rPrWKowW86AfdpaE0N/jEJyKQOgg2G/RN4gFmNOSBX
/qQ2cbTaX9ihbRqsBWUk12WTYMacNvZ2lmMU0RdHRb3SGUQziftCurrUhboSZhcrLqaQ2NyQDe47
MwmhfFtjxUxY4H0LrCPkznq1kPj4HEN8Nu5cM1a4f93IRlhNtY3WtUXy3sMhNfJGHOMILnxkbk/b
n8dqQGL2QSh1yJLAd5Zkx7H5cDgyuGUJ2C8tOQkhi8JDWikX7m6rVbI4R+RRw9IDIFwW+hd7VEWA
PpJ0f6/Wfv4UJSZidiF37MAOxDf68UhmQn8Qh4LxMgdgULagd+ioqWwECM7A5W/WltSfP28hdi6S
nTyZixnpAJT1kHyng0Xe0nMRJdOBGnwAiCCo8Hv9ARk+TyE01HjGD/yoeao6CBVv0XgbbbuuGj69
Ha7NhQF8DbGXCxRKhZeT/oeOnH3ZncuoVq+H5FQw0DQD4wHWWKCdHTySV99sbCSjYguDWt5HP5Fj
oNMvA5apA0dtIzCG9iH/+wbAIc87Tz2m9tkqiG4xL5NQQqRRAMfRYXmivA8kwBaNQtJKkTc6NHBs
nkRNJ1U/4KPkLhFcfeHbB2LvywArx4krSULH69ik6EzEDNurRqrR0wB/6oNsf7OonOTysDWvxKYV
ko8nu+vXMas7Ba0W5eAYnNHtjFn9Zn5H13Z5FIaX9tYdCZImb18etz476oqhBq3XMtDTu0DN9uRZ
Ck9Ou0xBed7X7M50CbwO0Xn6ZU7lMHaZ++dOC9MoA+4g2+9FP9kRWqilvPKCnbVDAwlSekiG/omT
qbBv+yKOzaJU8w7piegOC3Wl29eOq20qGOgratFMAjK6yRO8+nz/yRgmkDDaelShtKfgdDrSGO8n
xaQVpXuZ4utudKfqdH7ifhxcNTenMg8MKvZonG+uyRR2aH2q8ezuQuM3OMFUFGWemIpcOKLp0Sch
vp7Q/8/NiGMWFheuKhEZvJpBvYn0XaGq+khR+nHrdtOVlhfuQDZMuopkSWJkI7gBUFc/9ekPiBZo
QlFcgHmK6ub72ypMgFGbwBqWt08CwInBL3WtI+TqlWHA6J83fby61Xv3I5Z8BGO2ApwsLddtDdT0
JZZmLeIpXUdDdb+wnnOZPfF0KDmB8ALSNIQEaeZoBlLwceocWe3AactFuL/7pu/SAp+yUYI2UtTp
QkuFGxlIhy+Z02MTnWehX3oA3oDelpMe5AQb4YQlIIhCGz5o/+Z+T8nWfBRcm1Ozti0Re/fOoRrI
FgwgZHRReXDMXyaWtShca7NCINS+QU6rVLV+puzbyMJVJdZPdorcC6NbbysH0HVXx9wo04K7fhj5
fWyWOdvGXVLKXjPEkCqQDZhxmGqINKtU9alIfnHyYuk5yirA8bNu9rysxj6qiqMV3GMXGWaU5jYo
iW6lsx8exvcXBfyhXMDgXX8pErFSncMrZ+L3y3eUIPnMs+3U6oMLNg7f9c3v/98QHqeqiuy6/8An
5D1NkwWNbQTjnO4cN29sIevN+7dVamQw6V5bmcc11b41NKYNc3Z3nA5tPIHb2EoaVh90uoMpj+KG
um7rWuOtvPEP6oY+NfC7/AoAmlUR5GbmooVhGAuF+ligzkAxN/18vAfdtx+8Qe4pqLktjEBH3uVU
dCb66Q7rcJBSLogvC4Z9v0iAZbRdcA6WOqNPkFc4pWURktGvXT8iXGIVRgjsZdtp16FCPQgRIqlw
nTDatLqrjsmsoDpOa0RMhNbmBF4Fau0PwLf8cDKaDWOBs10UK8mSdmZqXp+atkrw7Dy1XcMj95AM
ujJu4I+ZymkY4j/g6SnZvma32ZNw7kChnoTSVZYEnQ/hoTXe8MJjIHVm8tY1NImvUEu9b6Tzqi0e
OQkVpJUEYeob3UlK7WchwGOKPvBE9jDtCu0gBilPlQMF3TLT4TBWL9YaBdzPy0fnSHgaxeNrK5XX
CqTYDYEl2+xlecPO7/Za5x7Sq6FeBHSwG2O1CCtnity+4TztKRcpgtEeUt4Ns2o6BPxPYmasnm8e
tmL6PBi7+Yzp8FQsvAsPx4ZzCgdP/Aom5Tjb85SIkDN0CT9fxTEhU1WfApsX1pEdbautdcmvmjHO
4zj19c/XWfkhGxNpUde53g8Z1frtVqby5+z6CVFKJJKyQY3mIDwdgg3amburKer+7gO+KyWTr3D1
7padV5rkwNKh7qYLRx1e6JokbV9QcDUg7VMjtDW48eS42N594cEP8SZ8cFEZJoLFPSc4/50dVmJT
BmYRdVcZ5TPOYph02AtRcC7t+6JxZIQ7zbHIpTUdDaPFsJ5nfX9ily3r/9JvojXOKapXkMuxcGUL
+ZKOdXen3ftprnkOB7MKyQ8/f6nI3Qfn1Bi0iLYI8cggd0nk19TbcP2ulZCd74cgnubQhlV1ikcj
XOy876LZ/XJ6qcG+z29bPbhgD3yvyIn5DCbcOXSBJU02BOnmRN38HnybI4qVDaSYek6VYtKFM/aA
Dgi0yc++pWVnOw8wquzM0r1xpV/Fawh7yvt/jRFVXf42cmbMx7FFAHfenopNTDz7idXPFrQjPp53
k2aT6+UV2R8ZHrdl5dtz269CdoiB1YKQO5gY3pc2PIZZVHXFC3ezIwaEytBhcTMF3yPkxEOXzBTj
RtJjX1tp1hmWtSAlsb+i3PlZOHRvXVLQDISkdiV++w2R0qV6qnVjX2nWilWtjSGCU3KgQ+eqR7ji
VigRHgOL6H1R/92K20fncUP9o5P8qofxY+/hwGYjQTD4+azGgV2b89M8QxqCLZjz5UxO/91CrvAF
fwcZFhvizjqAt5AYd10UsBowTZhHBQhqLI02y6zGVpMEMawSxqapAmhumE/OQvhdTmcRJrlR/eio
uxHRHeseNB7qjEShQatqT4p2/ZpG4lwCehUXh2t5ELnGATQprbOAF4iWKKfqsCgbVMUDiWy9xF2F
BoEC6RoMJYPEzT/2sdF9ZKnCvLRkVG8fUTzYIojx603d0OFdY0bYcU2+bGfn+ShHwUKQEe2+bfeu
ij86JpOMcdgDnFLkoC6birV+y1Ko74cKaqJ6fQKhrmzysLzexShFqeM7io8m5FV0LfLk4NFb15f8
xVSwVkO9MPuGLCSkorMdQpUn5K/9FII+2cSdZeurKuokQSyN9ibLvjoZ6mYHjexAzKnZ3KQrZD0c
uEG/9DkJ7EwHH8hMianHAi9qe5pSlzOYY9D+cNm7Bx0+Kv8TMglc8s68jmIZt9dT8IL4U5V8IQvC
in+qfCIxq/p4SxEPm+9nhqDO3PbT8FxfKlm/959hF/9omxRT6JJSx32mn6VZ9y9WGZMEmNWQYXxX
DCr8dg71r7dTTPSVa60q7muiUNLaTCuCXFxv7bNgzQkmkJfaguK2W3Xwlh38A4hdyvQPeNT7LTay
f/nWjytEhpuCIr4vyIqaOg+WQH9tSjxNjUbfK+OZafbRnmVdsU66Zovx9r3fjOpbrm+SAVLXzTVK
31jzEGhfYQYFxMhnzhOS4Amni2KNJSEWDh0FYhjl9re9PwwuMdMi7xAX0JOtYLtZh8x4hY04YYzW
VEIEr6q2NgLnNefg2jZvFMvGv2MK0YbPqIraMtbIyumtSaR3hcQorW86wk3jAjIFBCb8M0spRcUG
OzS87k/AgTHLz47KONPOgfzt8LS1eZ+tU3Nr0QysunOxLHCC+OL4P15w3aGZqCpny4kd6R2p611M
xAXF0WQXyP8g2cMS+cF7Zm6g6IBMwwDPIyHxHaOYtwbXMtuYuxuZsw3mLYKOKncakwD1Snz5UvN2
d4BW2NDr1rFApql1hmI4qRY0If2y1ErTazhz2DVduN8NetJHbnbcBNYcWVkd/dl7cg02CAmJC4/C
sz7nw21PMJNNz2pfM8CtS7tyM/n+fUKPoNF42Teu29Im+8f7jJOLNXVMs4NXJUJC2r/MvrwnnWVE
4hvWOiQaXQJQ1+LYCYIGTV2cDyPQKz5h8sJ1hXbF+0vATlvqEHmfIl980NqwqQwRGSZMCAdg4Hnc
flEBakVTTR7GJGoif9qez9R/J54UxzG5g4Xd/rBTcdnOF7fYlvaoWgmlSrPta/H8nBKw3GKBJ7Pu
EjuNog7Mw6SuMRtS3H9SoIKQhq5CWwecq9RPZnm9nJlYK4GtxNBukXh8e2cIUYqHbe8BVDx8T+gV
FdSzYJpxj4dMy/wCS8kPl/00ODxSnRQUBzziej7KiN2hoqGGeG/GKzPRPGCpP8NZ3521rqGQ9MO3
nii/uvejk7yOIdbaDYA77ev0wqiNlDz3e6NKten+AiuPjAqBIadm8Xub+bd9K7Y9vPZaTk4oeE1N
FB2qZumg5FEgrnonB5T0QiH6VvQ/5HP8TSF0zorbWj8iHRYxz+R41z5L2lIdVi7bwUS/oXgSwQ9/
dbcHjDzKjmWqRb1lQ0Kzd1vwwQGKSK8cSOfIQo/ooux2KIwC7cyreh0GJ9CWFvyuaxwnOXXiWTaM
fuqWgwGZiYfFFm7f2GTxEeY3md2dx2NQDJMyJjuk65cIyXABYEZs6CjcCpNJ9hM2+hIC51IzfThV
wGwRSD/4knnSSVG7bE9LxweAFlPcS4ojGqLwAfyLxQNelPehv5k2oZGRqnQPOzDlfDrqNqtZwKgc
Mxd84253f11QTJofvIIkEhnQQgu0wJ0DOSI0UQXOXteg18Ha7zfpJ9h+0ahBrwWE0T6Tlz/CzcuG
lM7qawd3B4SunHgPcBa/wuUQ43CyF3MHuojuIhGlIljDmD+hEcaQ93Sg9V6Ui0ddvgfLuXAXarIC
DoK9rQylLKl5UiNZIiv9ksYjlicxeZkBDon4AzReQWBDXSF+D+AfywPc28F1HM3Qp0imgvd4wmmO
1kHjdg0//zFtEaLVogj+JXxgXNeKTE1A184cbDsyyBdZmqvOg5KehStVbhPqXGIA3IY4jJur0pNZ
Cc7Ejyb6TcCGrVSVW+HgQbOFDQavdoAvjCM8DuBvZj92lOFUB+J8Rg6wJQb+0ILQ8xtOvn3u49tV
kGESpdL1hSyeYUIj5kREuGGiFW/HwJ6tpEaLIkFCpEaQ2Ck8oHYTzKns17WlqXmF2BL4h73UY2Iv
PIWDdgSt+SG8oqYEvUaL/Csxe1dP/b6fRRDNT7CFZec4dfe1IGXtB2fVz+wpAllLwWI/HVnb1Gzz
ZPpffGgaimKqOnqddW4bo5abulAAGhiYNEATOW9O9+xhmQGZEkWAME7avLQxwkhqlqBngnwiNI3l
UWD8CwKLyrdZiovAIDScb+Jw0pGpUC8Qv+OB5vVqGVva28u6Cq3Mr164WFaUukvRDqH9FLbhTbog
YfOj/Ko1tnxT19CyVXhJOCiLRsZSB5wE79pqOfSHQrQCshKwQ3FpM0BbISwZsfgcSso2s8SiI2dG
pYqkUxBVxpgqwM75jfRPaAYMkbGv0l4kyolXZYu6TxfibbAQ8hNA6AIF+BnWCN6somA6fhlnaye0
zTefSR3ArADqBi5AG4KtzG1Vz3IlORpWef/HDxad5FtCCHJiVIKwlybSumvZPOx1Ro8AmRohF2ZE
03CfS2Mo6xPyHrXuIH2fZ+HpX4UTEV3JpKaVr2ZHimI5mWhN9Lvv0ZKUtH6Q58OlbzukW3anBbd3
Zkg/VUoN0KGtr38Jn7O/4/v/X4eJ7kIUXvaLhmd8wW5DihQuMUN3OluwazhIA5PqBrQoW5zbg62C
MS1ndbz+UjzTncLNJVHbveLsMvqjHyRjK8m7U3roag7IyoiNSW48ZcZ/tw3/U2x/2f2whQ98VcAR
SgW2vn6Ux6sOPZYriUL9CfaIjkR9zvnaBMED6nHScmyGzmxRhdmqchN/5G7K9OWig+sKGZ6CFaMq
Gee8BuPQQNSR2OAKPPxH04iurvu64BJ/wUgkDlF5/+3gi3q91jrvLQAgXncqQ2jhhna2S1E9zi4v
b88bbikX1GpCqTRQcQOD3tKX1QrLJt1dkMHjW1NC+w85sOg/5B/1iKh+oZBGP6+AWThKGa7vgbcw
4cNOt2BvF5AmJEXdCSB5cC/7/Xw+58YpDvrcm3sn9bDfOZduJ2cVrTt2zLFC68S82rY/LGAaTq3O
QhOtN1YFPwnwg73UV+DLw2QJJm8Diu82UElH/b7OronjmOp8HKT6cG8+HcMwRBC1OooEOOJdBcAy
jKtaJg0mYY3R+ThtIKbzhyQZiaVGevsJ2EH9lO8HJP+mMXUexMh3Pkk6AajGOubovsigLEaba0ly
bEfxeNce/W9L0rw3u5BP/to4pDMj4zpvvhBGI/LujxzULEibK6VRKmsobt7yBjcsI6RRc+1biwej
sig7M72KHYwfYxj2tJjIYsV4ISt3dcvjPgnsnBhOL0z4wOlkCBYc/djjICOE8h+dWnZgE9xERA4I
NgVt72mrCINSOcPvlihzyGlqy4PyFu6E+JXbXma+ALf67sT75SuZBr9OI8v67A8RJgW475uJRgAB
8jY5Umk84ZuLfxgU46EkbcVOGIuD+Er1eg8J5VnQG5/jdlVlcEkIOYVyK4nGV22LJ7uGBA40wbre
Pckt9LtEhSVTu0Fq77htmQ2pM+JiESkIzrfSuMCJ+ehA/ZUa60fsmpSbQU9VmCB8K8wAI0G3XZWn
r3LibpZFraT6hINHE8GpQImbsGz66T+5pT7/TVFh0Qq1nC8nR3uokU8cXPwNJ3P6+XQCAwG5+NQe
ANiDc31OF1NpmqdWWZbcjkZyuneViK8EEQcUMDYgdT3MI5nxtDIKhjA4o29cDBL9C98cmlVf/JWj
dIAtiVdOGzUmtQ4uKUroyPFQjL73D6c14CbCHyRqiJJcDCf5xBb+qdMEL9GANPjMfQGyeIFbVT0/
tKSecqgoln9cJVSfVBZiw5ZJZWnfc26ejHKMoWf3US1wkBKrZBEPoRsxSiYJ9FLmubj+XtaPAXrU
IuaWonPC+BHOOujiehLnhzt8QvnOIWdsrHE8OxzFiJPbNqwG4JHOiA7XiPph3qPtl0d0XBdHlt8K
v7//fyosmHwa73OO/Kxi+Fu3RgVfWMyLrCYrL2aJeRURVC22dz16seXxIYStucbNbmCF0q6Ig9Of
kEnIIhIV/6+XqISqTPwDxbXtlPtRRb84ITuCEFLKci2xGs0F/TJG5qlYQRP/Dg+Ff4r84M34Lemg
9loTRM1/Je0qegubmX8G2Q2iLgNycIxKbIG6qMwUCEd9y78zlGtof9qxfX45utNVT5WpGQDUhqtV
ViUPJpRYK2YJV57OGNY50k+Qd43bYkoEwJRYIH4EmEvLJifTzi5LdMxpXUBFRT1wnI7aIp1G8FnA
fzHZPACYVNw8bQ93X9551VzvL0UL+acG1XquZYwrXuCXBWPg8zEKzIradvTbXdQN2eDnxwCNTZjs
rsE6nSGbWrrNkWlIAi/aSUYMiMVgykzytK1rAQfLOz8ve4j8v2b+rMhUMU5NVkNjK9M2ucFmRqck
LD2xt1vko3B1VKAWcNCIfOBCXtpcAvH5mHTd9SGIg4RrkTX7ZndUrLzaRFVMWm2UNkC9vIyBZ4gY
1Kuxtnv2VQmfFYI44/ll8iSvaDeYCuhL2uuUctqtD8VKyq/YqGhsfrF3yGDDu/YzxWvwn5d4qV84
VoK2I0W1hzabLCC2q2qIsib4o1ohb67kbOeXW6mNLBqY+59Ceta025aT3SGCznc6PgG8bNQPkIRr
R02hlpofmySG2+dWS3ylksC2mtREyXPo/ZJ5JN/2ylYwJm9AYJwvAph98nfLJfNW+8m2IXG7rl7H
oxDjPvAGaykYqg4xzY2nlmpve+9zQAa5OnTe7Uu4mItIid4L5wcMRY3lbOhg67s+OnX6Ko/w99m7
yw/aRAieWSEt8QYQOA1IVeB9qdPSVvxmFAR9XJIBBmxRUVLUxpLe8V00yJChPISRxQ0gZQ4w+4Ld
jtjf/lnutgHJrUaS9VxdSXv/qTFZQDNf9bwHfGvobpNAInZr31IN+u6U57AGTajGZjww2RKLkqBD
GH7uMH0dhLSdyOdcnHXA2nJklN6hc3iMSdKCjWNgjTI8rWzj1twvL9bQr8CGIB8tDDGux88LOG5Q
G+/L+emknTIkI0m6DnX5bi9kMKZg2DPe5AnKF9uwWCSpOkxFF0c8RVIntYSs16fSAXKyZ67adwnN
BSfXUhdut1/VAfk+w1ed6kLXO9sWa+D2eTJAHocUaPOJJjvV6ktZe4afvelvk020EUlwmzjIoC7m
Iy63vBu9+wTqXca0GzBhkGPOODJJoZZ9Mz+UqEc/AdXT132fYypKnQmp0IzGVsSaz2n7Dq5pt6Eo
kKA3sUh6FvcE2y6X0+/HCpB06ua0NAVQ/OoF05olB8V18VLSdX/J8+k80Sj7dwyQNP5NN7yl/BB1
XWIyqbTsZI9ocg/3AfUNQqBr4fOFEExckCUHPHN18S5T3K5mCjWdLsdzM9PA6wYaUVNTkqzEl0XJ
4zM0ZtOYFHjp1kjC7yvk4iTKJOnT4E3sRq2+feF8Ia2IYOlM+K+cyoEctsFOyGGMK4pYL3VeJMIi
VmhQsgD2K9ahK1AVbKk9++AIlIqF58Evp1NvbYZTfF1fT38Om7FQcO3Wa9jIi34Ozezeyw5tRJo3
EjD9TJClM/TpXkgAtTLjzH1B8ZvRfYFbdsjYSN6HaPl5mSrkGPD+XaPq3S47fwCIef6ASocQIVV5
sm1eLwddgOjxQg7M39UK2bLhpIcDfCsOI6xQLb4Ae/5j2GBoqE5ui6iQqyEfieG0uDGj58PZdCv6
UqZpi7XHg/HEaq6TWAfE5PE+bnbqIckdiJmRb92JsU7+nBuAObR90hB6nEdoQa+NDACKc/wJJKZ/
1PGyknl0w9M1ONufx7OnZj3SOdbiXuV6UR40GOmOCqOTrrYypimcj5bqOkdHwRcIaCV64D6VaAaY
iljauf9+rKxy9RpQPfahJHj7NzNjQ/VaEZ3bMuGnhNHhXbfCLLBxzHw+3Ie4znYosLlmU+3jIPK0
B6LEzSMP19xCt9tztOGNKa7gGSqv3Oq5Re8Iqrwq3b5polzRTOPfHyGL9O66MNAtizQEWyhs8AEq
96S5dQw6DYUU4Pnz2iAcLGXBKCerHQvVYjgZfCnXB4wxM/g3PtAD+6wNUjDGB9kFxguKONQWtjz+
VrNJb5EQLH5jnhfuwpus5yxJmQzJCSugKDfLMDbA1X1S8RnYV4ykfL9zvjid6Ah1SiyAU5phY3rK
R7NVWo0zjYK9sLA75ElKLvIAdPolqmJkNXXS/ADb/dkK/N2fUvywPN2bpdzPvrnhQsDe4pPKgO+e
7uG7UjpJkyzP6XFqU6TLhr2KWhnhgQOY4tF2ItudoiGRctNWo/AluVggKOMuQFAFVyn77iaEo8DQ
AS9O5Ef+1SunAj95PGXZGAyfrTqxcK/tck2x9s9GhfUgYLGjs7mGCbqscYkJVCN3ccnfA2TPRV8f
fzwrhhQfQIBE2Cdt4Ar9j5LTaQzfNma4dvmt9fxIb5Um4iYX7kvlZQn8+8DYCCHtc2WcsNalGIz5
/2uQD8pHWRNKwc3jq2i1iFWpyXiRHDwPLJciHFqgx7FJI/3OYywg/tHfJ4hjGGw5Y4ESnWnBZMWQ
sMQqwP8TbjWM27RmtK2/uD+wrnx+O4SGonWWjsKIhkPev18cvzXYQL0Rlne/Hjf9n7J1KSc3pmYe
haLaytCGghqQSxX/me1SjV0cs0tsolBcO+4sM6Zap9Ej3Dmi8ceO71UyagSy0HF1LAIv44piTy1Q
lRf7ED4nC+YS4E9+tjrfHyTQNQMpDX7gf8iBY3K4IYM1sh65aBsR+8Zs9BJn6SPlTlYW+Z9YvFrm
YeDdfmYXjDPAbzPJElMU5RT5z5VI9mFK7+Cyd0vfpdrorjPM4rt4f6Wlq9WQIWhX4UP4abrNfwQk
CkGTAoBZdsq/bbVNWQBLKLUKasglnMF2NLDgKJ73F0r7NfM1Ms3U1985SGsdirYc2V/1PYIAeIqH
f6MHCL71ErF7WPhATfCxR2P4DFIFPeqSQgFAyGHWmVL0KT1MjPFRbdVUec/rcNryn0Ogn9vI0vMP
l+4jbanNt5O6bY/SyA8vtL1xjveA2i52LRc05/Pxt01Ti6VZzkNa2nxUbPaT4pVxsbx9NLMZk9zJ
Wv480/p+2ewMVLLnagCuHzKAtCmD9kr476O92KjU7ZMSlhzi7hNJ/j+boPuMfqx3+xgbNVn3d95A
CZT06wUWuoAAvHFJqLKwBWgshy1Oa/koJQ/2ohqDQ2GNyP5Zk6jzuCTz0by2rwmIcOLTRbUb5Kjv
gRqWT0zpSsaJ6SBp2couJNquBIABDm9buSJzhPT8Z5di4zf9KI0rBMW4aotGFpOtFf4FvUu5o/PX
Ux87jJBtWRwkgFG+zrn5DVrQz9ANDoTfJB55T5E0NW8TTMS2C5eUfwp/SCy+RUz5cKCtFz+rbLp0
h+WY1sAh7vwz7l32e5952P4f7dbipMv1PCVj1mcL0gt4nnMlxqK2dBG67nkGrRtjqyf5jBe/C17D
EIEcQh1I3M7lusQcKLlO83lSRGhHZN1D09IkAZ7YPSlqmgufbKibYWClLTyvgmjiPkEwbDqod/3X
1T5Q4Ipq1uwOyqAo8yPf/rScmzuDFwNWFn42mYApYkM+54P1M8P6bUZW4TkEOFpOMYqq2Ty0SD4w
T4AFrbr1+6BmzCG/QK/mPyT0oGMrD1sezcAM1AKQES/VJsSWQwScOsJV0U79LEbi4XJnXpft+xeC
WCElO3p3FZnv3emLWZg3jyzcSZaQUTHTaHwLkGXg+yWzsnf13/rnjfogSEqrXlgLggdxxKYJxX/O
Fu+vHU9RZ8UDNlJMZH46gIeGFE3SF5C+/+4y70YFngeEB3Qgl4DbrFEJV8jVd89hW0XpAZ45IhUm
KDRsH58H64wOjo+y/MFngTuNQvr6bMdT9ZeSoNe4FuqZhZ7cFn1hPikm7cUiQPT9EKXl/FewvDaX
QJrSgJ7qZaJy4LqelmSv0cqy4CIbqylqT1DW0E5G2ZUX8WIRp1eHEBSE2wOVGCYEi/95rKDaLQR1
hPMK83OxtmGgJo7i2y7KtTRafTD9LKSIjgc5JAKzKhF8b3T0fRXGrvdqX7oo6kZBiZA7VRC24Hhn
dq9mRPnp4+L8jFe7q3vfqX22HyevKPjw/xxhxo4h87Z8iv7L2e9d5PVe1I4AMgOrKyRav6f2zn6a
KayxBoLIYA+2jMJZRaxDDAGw3x9/B+M6eoUQsrrztmCFHnE+ukyZe3tNCMSccMfoE4zzIssBCfkZ
+oVEeUNsut0R0ZyiQawtU2WQs2S1KziYuHewMgxyLBpyha1668gLVSU4GrRx1Hv4weIELFRB3YJx
WWkzRx7GTcvZuLJLWWL9zmyMfKA0cnkfgJoO03ahmJP8MuWYhORkx6kuJkZ8gf/v2a488hbo+1K9
uWcC3koPJtMfUBXzLRxdJcOOUOefXyiesslsS8VqltQMrHEhXJ+abx5h3qZzIUIrdPcXSqzk2oRu
OzjfvLRDpfKPeRzbzfOolEkrLLxDSWYfxtX50I39KbnrNqUXyso5bkzKjp1EObTtaoORENzl/phN
zHeaEYvcTQ98Utygywu7CsjQhu9ku1YwEcJPhHRvKCy+XGF7GaFObCO0LuEq13w2hg+rZiZqCIsK
iDxLPICK9g+JpSkI7LlVy6Dgn5xjsQRBrBMtZ28Tf93jIAzhV8xDAX0ly/CeswsQWdMhddKSJTH6
JxBcaTG/AEtZedHg5LQ8B3NOIXvhijiyLdwR/EjHCaGHUtRZRVKAiCZSu0MI0MraQt1K5GY3RZSz
WW0db61eGTK1k1JmBxMDlq2sDSQHTkAtIjFZ3B+TgO8HTuvJjwv9ADpt8ac8MtHMbgduYiGSAXHp
DTJ5y6XldTx34YkkaAXx2qOougVxJDhbLAqX7TKadvS22hxklTj9tU0ypEv9N5iTtPKld+NIdXNK
dl19O17PoYYorVKkvsg8zbsQFH4rIpvWVawt1MQTtq4Ac6ft8OU6OZYMxQt9onpsJtlomYGhgZPY
vXHLCoHZp8ReIBQ8ERVd6q8CyqxuG0Vhku3hyc8CwYO3/qJUKdrvTkqUJdqYr5gdvfborFA9lzzU
b4e7MBRn7yzhR7vpzLYf1444lY0aPl1p6fEJbSTNSdcI67/oH1Z/80kVbHQl3o8BJrKnLj86//bi
pq3J1o55pREbBvXPcZbJG77zFA0AWW98QmX3WBTWDGHDjQz1rOx8SA4PvCKbiv26e534+Qr2UKZ1
4r1WyNHP96g9Gj7aammAbVujqueMBUuPHjR3lB4tmqQ6XLqXgSAI8iDtdIhQqSM8bb370eseZhNF
eh8niSwXXmJ4d6keyqJjNpsVaYfjjWL8pO0hHCCOxLhABaI0dDRObmrv/3+Bqs19UBEM9jRZ4kds
pS6Fhue3wsbbu+v+PDGEqv8LFK8ARByR+rc4HVaoUCQZTsmiEBzJ85QCjBn87OGXYmkhgGxbDw+Z
foOPJKESIb4fP6kwGPkU84VaRLl6yS/shsSDXrQhEtVqggtAVgJIfbFEd5ftSAvTA9Ti7eZ4VvVe
BNOOvekaZvOnYvAzRpVERgScM2AmXbBBVAv107ZjzHPPLgVBmM2lMvLsM6IZlQoSSwXxY73h95AU
cPYV4EXbmzjSI2CWsbfBL0jHbb0muJcuSZZ7R0cUTkXBFxXQNZ9S81Ro93imJccUaeBLcRnJo+Df
CyoRlaVP5m+R3V2PXug4xnTRy9Y34Q6hjRE5Wd4gZuBLHHqVVBGZBQcH3nVXjw8uIkEK6QhPrm+l
MXDsTOgD1xmWazxOCUCURSMgCFQ0lRHfxoc5gbciWM/1HxM6qsg/XRwYCMZX8BZjbIgq/igrvKOg
tI3o4mVBAMOKQisyGTWXqR8SE1Pr9C65r5Z/NU10C+R7McGDdDauSmuVszhdcTMv4N9SBwxLTNxQ
TijnzFSL+X44xWBIhcy9Ex/UwscH3WJkpugH9MB977JSxq8PHi7VzxhJBg6Dlnk3zPhhrYjh4+ww
FxhEjuv31P2dXmyjaE0m29WK5+Y7BcFpgcl9oEZDVLPuNIU7tlwUZO47uq6uw9Uy5xkG+vlIcUM6
9YGByFnPejRDa9MTuZWmR4LYFfLUjONKHERsakrNEdX+kjBumwxwbokEFSw4lU2JaK54YxOjMgDY
RE/kA3vo4pwX+Ssak8PopzjoV8IIwOBXBZEtJ//fnzRij02rOJWwYuZnXeLOOs/LvJ/jzgV+BLpb
8Q0SgIRtJVeRyLclix+cV8ZOCsTeozcelSt5CDSsNgFWM09tcubqxdM/ZQixzu6i3bwIvH6R3+1W
eZZUoEuHzz3Q63qQyREOrwEELQJ+Hp8UAIFaTJB3ggDNC822IgWclu+tYhs1ysLWiaoGo/xKPKJs
WJmonjF5I1Tf96MsFxZ7LJavU3AZxYBzcyYndmB+NTYnIY1NTp6gNVjUFE+V/zqX62JJAOvk1svC
PA0/6AErySE2N2q4/s271etcesHz2teRfJRGgzxKY10DH9sLJpISESBRYK4RSlIjHpDjlk6hn4e6
GYmrWHpklSg2aPYwoZcXgENddMeVUVpud6TN3QqUVq3/sOieNmYllQoI/4lLb24/bv3LD1XnWRUx
cn+r0ktoflLyEecYgDpUwGVaGvLSw7AhOzewEJBMFPIieQIg5mH6rOusVuEmxvuMvbMk0wGMRUYp
bO6M0Q1lST8iUDYGM4WQOkBZFIXYbfpMStHQu39/GrKVE9c5mubjTSiiw7ysVwW997qQRvPOfKoI
pSYg0pttyRSoKPfroloA+25idy2RuvT2AzF5Pifvyc2jDRS55pKaDaPGdk8QrOuJSS860BHfnfKt
Ab6x3sGH1xr9yuQH2ZSvEtXf6ldRM4h+fdVsANgObT3rN+0y8NgN8Ri10YzKToF2y6KJbZ9Eli8w
2kVDMJqSdzFuWsipoSijkEWrcL/o+6aLzBMq4whiDu34VPupZZowsXvusapPZKg27/oW8hPVN9Pg
JcicONIeuvgZo6ArxVX1XB+5llnzNivsDLDbBE/9axoeo124+6WEsHz9rK2LJ/XEVZBb56Z6FMC4
X92Ed7EKhX6veReFGwEM83Zdlif6+Zy70mcthGf9bC0U5A2Gay1n+hpHUmQBAxwCqFurBsrvC2XX
iytDb47Vla+TkjOoR4KVIU2hMAxHu+vt7bOxU9HC3caF3L/EgRJpUUVnwLeChJX0fUrQJN9gNGD0
kvmqrFv/Vy8ZGGLy8eOaWK1x4WXrwLep4rP8U69tcVQZK5GjxT4ELu+uBm7SdmlXXpuRJEocmujt
Yiw+WTdVsxyNiHk+0+2J8++aHp3Z6bPECro1uYErGFKazhS5x7sIvjlWBWu+tnGEbff1trVG/BEP
E+GdSIzcNr6/vxseF7sIpJWwfcqERazrP1EnKwz4L6LXglQX3EwT7vLABxEI3fXeWVCZdbvVjS+Y
LdxUjuo35GkiDk5QHZCCfrrmjCKirQOPYQ1OPY3aLi47jfmeDgnax8fcAowIgrqqGPC2e1q2v4gB
9JCNOAZB88Ralnbz0fvB9iKN0B+I/GxHdMddlKSdjO02sce6w3Pb8e+TSAHWSf9qMksPd+rXEKfI
6SdV82QRWQZ3mJTQ0HdgFXJFFUJoo90EqmOn6QEq1nEzlUNt6dEqDDuu9FFJfmu4yIxN3mtwgDit
7bCZ4frSn+djz/t5QDOi1x3Yp1TZXcgEL31argBm4ZY3tKS/2WPuwllJGJnx6WHDOiNMqiOoe1gQ
dVKEmGv4wVkC4afxeb9t/LuhATxq6/p4J8AWnVPQWpRmK5vARlA/7dortuVvvYdMbB9zx6Ho/yfF
c24AstoX+X6Gy0xdr3QSDdjutlv6i75yV2/dDc8zCeSMTrAVe8iQ9aZGWM+nJ3gY134RnLjxJ1SK
fWnSjJoyHhdiPb6Ui7mySUyaSji/CH/KHbqRsQ2xV1zTeR34oqzgX/6g+TR6z6dxItTnLSyx0t4e
15KgRU4M7bU5stuUJmHGBxHyuW70x1bd18YsAnsS9GZZ9f4sGEFUfniH3M+RAoz73cjrqIOumQLR
WW6eGdZR/9KHylkQPahsqRhQ5SY7w8XoQN1CqnYDyccxY2+48rJ3Q1sd/rqYSJt8RYlXqY6yjXu6
AM1BFQ8jN/8DvU6kQiriANVIrqCWcCoodNU39+Yff5RzdoH63qTFuyNHQWfEohkflOFEnzGMwLZI
n2uCkennfmLk6FUxs5Wl78fSHMcqDw2vuCj4WfdJXxKMTquPm2r5/tWgLMYScJux+JRLStWsbaV5
2wyG0xD38n3lMR7YxB+hbulJcHwkfdUvhI3g671vU3KrIYN5aD25W2MRApEzl6hpspxKi/o12h1F
hzyy5QKbHBFZ/RWPEw9o/qfjJElrECMDg52CyPv5CGmYgZLTrzCmpcVOF0wlM8+f2AGZBFq8Jcny
4S8uV72XLIO9T2c3fOSP6+DvGmDetTTHuvlKON+D2FX+EsiwL363TI4KWhyYtlhJhEnKMe5jGbGA
wK+yBT+Jzk55LHz4GdCVSxCOCzNZPUoEPEdyDE1avmf1TCnNarCsRXvRY1CiKTvb/X363gUlfkCl
buLommn/Vy5OgbukNUpI8abfw79Df84Fo6TIt1q6BlEmPz5IL7V+olKdy5EYreoq963zooSxFbZ4
Y//wXBf5CDEhMVwvJiDXOvPpR5Byt/9JBCavbKU60GT9ILNKDQj4/aFDi3iTDGMVYN0uFhoOLZYO
/ko/FZbQwPdelglN9XtBHBPvMICqH+qf+sQuTBFPmt9u1HvkwuXGCjEIlaRodu5ljNNM+fQFoNfs
Cc+AmEoaaux2EptOB+cm1kKpiTuKymKkPr5s1rA7Jyzohrt1Wx7kto8dlMI2iOsxw9jhFrp4CB09
a9rIrJnFz6gTt8OPzTwMVPJa285AtXl16TckzmLBnCmclI/5Z1dAOlufaJonwpQrKUxMnhIJjbkT
uockWBTjJClN2rcVjos92C2c0d421BLu5t8yKmioqemofumj9t5rJ5Yna8CEUNeC+WZYFn7gZsZi
m6rGGMJVcfU7qsjI8yOUClGHXtimbB2Jam9TR825wF8wV+wRKeonCFuGbmMG5elvg7AYBf1Gjg08
xaKbRERz5YAlf2HTCLuOKWhjTPeysl3sR62djvolR4ntLNP0disLtiaP0JynsJ4NGH58DM7YfQyY
a95B1oLvxjluBzClY0wKwgkzGou5FrYgIdWqmeyXIh4O2znTwfMFIpKQMc4gyDG0bVad3XjHmvwN
kLWyexyI1xla8dxAs4Abo2OD8Wv00uQg3Q1kYF8minqkT4gu+F6rrHRV/zcpoa+jWeDK5utTsAET
X3UtZQ6GaXvIVTUcuulvvojob68Yg7IJT7T7aEKjurhx6tYAjJh9hC9yrf/olsXOfDcMok7RduVx
yXWRE38kmor9tdqxAe9H9tJoCcMita1dT/6vrdHjk+Yg+YuhfJQLRaGXsa8ZoqjYJwUbeZ2/rLM1
buBFrdpUffARwohSd2hiziKt2bGSamfxclG8RU69eOyDHeef6ZuAr03kFVr9AxkfMwB/cWpnrCUI
NnKF/TBEuXg93cWcfGper+hWq2f+TKZDMPiOpxWySxed9ky9XwGstMjeLx8OcHS0yH1RFQsQFpTh
R7RuNIM6DQBZjf/2J5L61r80x1EIpZ/ME1I+XqAEjJuA+8oeCtJq7L3Rlphp2cVyRBwcjMa55hrV
pWXhjnPgWHUQ7iYnUmiVP5AAAuYpQuseEKQy+VIfFbGr/DumXBFL+AK7Rk2CAURMjENKOrM3hbdB
nAKlFO0lyFlC0q2+OzVtkLzimZ6Blfrvtifxo25gehogDtjL6QOBf03mq6YPuQSvFftGiWb+QgGs
I2LOPWkpJMr31c4tqWI/7hSKfJKlRRGE7inwNhuhw6vohAQjceN091aVYmMAUtG2X47H8Sa0k+S9
uqzUu71evcAWTW8HYVAZ98GumnlmtCP+LHqfYh2653dlco1XISx1zJvCJnRKj7Gymbn4u6PulTYL
nrk7xohcVL5Ytj2iU/Z5TLHHt8+IC6KBcI8gH6pH2qe5Mv8vgq/10VyANWEfx/ZsFMCRjhAIhMb+
hp26bJkjyIgv9NZuokkL0jHp0yVwjuUyFl6iWMvDnPnSdwk8g3n6VVP5nNwdoImgdk4vZFEAe1bG
fIUadJvLN16UYMT9VKFsKVI5Nn21gCB4zbWqetmRqTo3TSDsYxELUrIlJ+E8jDxT/N14OKwNAmwn
+SXajyYLIJjRCigvQJnI9RbVF++f6s0Ll3zjXJKlwlP1ySEuAuVKE065FpSkmzH3JAAlmlkq+F4J
WeCbsHcj3zxnqLGC95zNDJUniKn98fEBM3Y7h+Tj1tOrblGLy3bF/zGIQQ/MK0cl7Ib1HkhYFFXV
oCMUryjpgImYvSPR0U9iIJSt7fvfPU09Pbc4yJR8CHcgP1sbipcxYBvo+wb5m00GFa6FZIayxRgR
CIHSmzsq3C7biw3BgvX+JCi8oWUl+hKQjGmBJGQtYZ5VrNrmeUQ0e6eTxR2SCctJizzkFXEZS3Z6
rCRK/3jEjT0dEmzMhNHgqB6nxypRM7v/cV+WItC00x+RyQYfiQ3ry/LgO/8/urJ3VUpO9wgA+0Nq
CpMIn5YD0MpgST1nzhgFP/yyl8ribzjl2JH9ziJ8HVcTxbSCMDYkH+PdhHoLlYGCfJwN0owdAta/
8c2VU+AR/W53LRwo4IRZuegiLkJfKbT26Pi8KVqxkb4VGou/PEBiveks+4MHfT8xAiL9uRdGTVGO
HdI2VKD1I+i5ZQH5/hYH8Aj3+wY6Bn34OvbFxzniWMw/V1W373jrTSvzormSg85wgZ5O7wrw9QUA
OTN07IXoIRwKi83Wt2zh9ioKhawRUsXQBBs0+tqaE9ETo2Ri53uRBWihLuPQORnVUW4cdYr8ghdE
Bj3Nr3hGmn5jVZIDA7uSoJbAUjoBIMjUOEimJTO6GAujkpwtvkTWsNMspxpi1G1OU3iv46trMLU2
q2TJdPFY3opFwEHCRlnY/I2QORxreUTOMXZmwdKIL43XmFHmfJorodCx5zVkEIIeHi++alrEGdK5
r27wv1eAYPbrFNCF00QQlaq4HiKgCMvqF9Pe560eQcZGnfzZSVuYpCrl1Vv9CcsYRlw/msLughew
qSmcKcZkabkFdl0KSgn2skevwoKMKXlIV47YhPAyO/7fFtbPq/V9QuPG3KIIEP1WsmuRqR8heVxK
kLWxuBLFCCrKcw27mO9mRYATE9yfe0fWz1oC/NpPPOfT1YwVgGjNzYrokjNIuMM9V3rZiOFqXSbE
rBj0/cTxVqpI0JHnDPECYQIYGtEpDhNBg/LFJCBhy0JdVfawyHbaxdfYQGuETAghuZFXkR6Aueeq
5ozrfUGsa79+VfTL/79js56qiGVxcHTcR8j+VuZsQFfvZreCerkb2MbxhbYrTvSZiD3oL8l9iiSW
nRoMI9NEB2JzFWhHuna875vxKCzVuxzVqBQpIQJfLv3Aoha7K7e186Z3GNQiNyqdDFi40v4dYoHe
pwNiTcRnhta8Di/vyJ0uepybzLTxBkN5cM7oFfYvBhtlexw3bndU8EeG4iHO066ini88vk+IBXTp
ACDs8GZ4RtRr4eBge+prAe/WlyOBG/RheehXKOnBUl+UryrOdHkph0HSjUnFPT6PD8H+QLMuG4rU
gIjQClaHrSpauwiq0C4c0RjyDSE/H95Y2IIFxxOx28lcv+aCCxpJyIDXJIecld27IlYj/cRfhxqH
4N4qhI3/MgE8uubn63Ft1gBK5QChrpwZkVKnu2ejnQ+jbdCH/g7fZ19Pl8DRrx/3sDGX+GlUo2Cl
pJPndiebx3CLBZWZNuDVZm9zPaewdAcbIXPnS4FbxN7X/BmCouwiVXufp4OjgwkbZkfAMZ84XmHY
ITQRK2uJlzu3gGYGs9gd6WRe9xSNBPGlFnEFsLY2ddGzCZc7RySi9QKBZ+IrKXxNDjK8LBLgJ4B2
lFjwx/Oru9Wkt8MujNtjSptgP/gju7Wh4o88tIiwncmPklYmF7Pfsp/UAiPnHcCDsBh2bdYxcUXS
nliJ/7c2QwCzj6sSP6lFjRw5DX9LizdTTzA1y65h/xlftsMGVlk9ggmoHUtmxOnUgXF2Pnw/MAOl
XNUMA6gIQ7VVQ6GPl4xY2ZlDoxPA2RxPHQulzL52ujz+YJGF8HOrVtFJoEzZ9BnfGLp4EOSFBKNh
DeMIlrsLD9Ue70bXXxRThv61XCZH/QmaQlLXiAU5wrUzl41DwMnkkNUTAHDyUqCLDokG6aZebzU4
2Zct6yVWbvc+MF7apPZSZezimjzt/tnze2xss3qVIk8yBjjaotEfeIEvNsH++Qk0FwdBYEoM4kar
osisl4noZPnwxjSZtoLvePn7GdyXu28VX1XX9KV0+pWf5sRiI0Of52AbrRelG3Lj1ydEsc9kn+uu
4qtiSIFauOBZeLMFNy7y+DLFd252OxL+ZGgzRWpkDCzt0hP9oYgzOYBiUuALAUIBo2JgMgWE2VgW
z2Ts6mHoyGkTN+i90v4IWIuDtm5Pk4NyiCOrezJ4ngSH00MemmaOdd07CkLxUX/iV8reucASaQ9h
o1WisVdxRPPFNGBRenztUf7yysKPk+7Gvrdsv74p5/wOqUOZqnTxhxlqa0hiY4k2VYmeMI4126k+
FDVeTwg9V1Oxv0GtFfFlphyyjZuDioeyfIruehLrxD6k4GWAB6py7lOq3KAESwwCZbAKvD6mFXvb
kweE/Dg265sjpTjLRwNQsu2xF7m61feYGq1Yn2E2kTlL1CeLpEsg+03Rg+FtQaEvlfkOI5NyuPOf
bdFXP9OfGGXaAJ95WwnyfJSQVtTbnpyYv0rq5qwtBQa3Nr+GpGZlt0ru5VuLHGzP1xo0+WXiKt0E
7uirAEyuHYd4GVg5p8pOcFdwVXBd3c6YSjDk/DoAaPBqYr63ZUBpxfXHNPqXgDORdOi+o/BKPIVf
VV70XIL26jexaFJ0Hlmpb2RBBvFPR79E3gFBjdtHcZstVc08YXZZ0IW4G+ZYmJ06gkNd0VYUJ8zO
CpR2DS2Q6AKFi2nuP2UjQcgdDmbh6QBn1r4/YUylEB/liDLtii4xZOQVcEn5rJ17Jx5fdN9uE9/a
l5k+LiceD6IQZcRhOABYgb5Xtf144rxYc7adf8BANnKhUaqJOEJvO/Re9mZEK/BB7rVMdOwtMItJ
ajNSMs9PcXh8hKEuLy8ojMTis8wnDQ2bcZ0OHCVlSwmrTlgy+0aUpMeogEuSt0vACA2UC4SmLkT1
Rvl2aUPp8gPdaDwJumbaoDATglOnlZraRRuxSUJmPmJd49shqRz75EjzCqpMa3g8vbPfDTZZew5g
BucpiUvEN1vXknv8Ndep1H0syHXfpQRQobYoEcSlytdb2KRcggJqpdCHSVngXOWDUcq9YBL+qpt9
xAjfmN6DG1LTTKSDchk4Og0rUWelfBw07Ch/58PgTx9RAcm17/BRPFOz15aE0uoTyteyVPpnR7Ae
CxUcse0LzEYjDGUi0IwQpJePPrRhf5iisHoQCi94DsGgHgrLN3vxcz47miCnr9K7hgYBspZjD6UZ
z2rNDZ7GPks2vANLHtQAne4Uj038nUyKQJc1Mp7hSUXkK9uTrBe/aYs0PfRCKph/aXgWCtsvNOJ0
Fz269CGabbYxND1hmHs1johUKt3FBDQdtMHDYHJsK8lI6VDiCpYtwpbpCiZhDs+Gq1497uiqYAdm
Bsxzpg/Ra6q1g77g83m10LwGW+bKkVkE3rG4TU3dR8DTK2ymPFNVjDgf3q0Nc/MCoU8e/n3kBtEW
eTJvAs9RIABMz8Z/82mdSQIuNRWJaanPFCBxf79tYbGavchJiIJNVPHwdcoye8GwjfgbVHAI7aWI
yygb0SaLm/jeW98P4PFsDOxOWEvUxbD13MAzUY+lo1GknbR0hTQAwaMkPXnmB22J3eySMQLOIDqB
zbYx4Di4IUgJy58ynrTrSEnm0Cqp/hn7Z4co4OTalYoLfNwfuJJmKu3EC6UhHu03JM8rG2JPYFm2
v1U9X/pb0izOyqT7ydR5jTafcOzBjvDuTVRERoSqNURLnJn6GC/2ihG2f3yN9EVCiUHDpGSlPfmG
T6+bhvwq50nijcR3tZF8NAdtmxWotwl0UCP3Pntou/ZUNoNP1n1vO/Qh1qv+OSJohnqyUtzuePWj
pQtkOzNh/us2oY0jwej0z0FuW0i+Ji2vm1sWBAmT/Nf9cBHzGSqBRLpwbk8BTgzfoipVUVO8JZc4
uDCiIInydVadaxCstIZc4eG817LHDnuTR6G0DBqCFpkZu+n/NfAlUT37oEyjLG3KlUztlPv367ZS
g1VNiA9gI81Ko3hBuwfgKtnaafvvmgOESPtRkqwu/hVRDYDiSm2i5VeFDKKEeXOEAQxzP/Q/0DnZ
NuJsyNLV76u1GTt+3D+2qZT5YYNklBqJKzZ2t5C/g8abws0vCnmcmdkmBY6lyBW8C22trivDdAUV
Uz5Dg0owoVRHUVek7GjoRIbZFakLGZ5qS8QbrvXzB/MDeo1/Wdeqde3GRZDGiFqcGn4cF/Mt6Bz+
Y2ucWa+wMEdF1tbLPaXthuIF0sXHKU/Y87+DIzavaYRbJrWt5oY9tyB34WCbiNzB82HRQM6Vy4Lj
MBnrpcz9jp265z685HLElsBIXOGTrfPMBSu0bTJJ5AHMrbF1ZY/A5UnxgIMuxjHMA6z26dK6s7dC
8QobQbVCYLUqivB46APVWeAu7a8mS9hUgWaFIPDGsVLzpC41gm+hTzpjrY9+9tr7LTjbe4bsmFNl
u88jAQOkSo0m7cimwUC5hOPYO9DBf/T12QqUFRGYyyQf1q5OsnuBaPuGQrfXkl4FLmnNOgAveUqp
z5SFUUE7YGbHslNXuUXVeH/UyCgOs2STDXfPJBdLKiaBOfn/lKthVkmFJ02Td/IGzw05qd7MjF5s
sdUoK43ZWZG+IcjUylkD1ft9ipAfeP21AR6pK6XNai1L85McJXq3Ljbfbmx/1BcBH6xqpJd2hYDY
ksoJ2k99uPu8pzeJLhG2GKhqYiXHbdqRevhDjkK+PTApq92mhR3Zc8fZp8WniFccLCwht9iAlgUp
KDXMsmbx2Oo+eWXV7qm6EvGpLPMELBEdhMXaeTTF1SQ3WT6duc/Ax6O7TiLQC5GVdi5nFuYUKFZk
vszhb6Tb+25CqFFm6UeTHJPiYXWLFhJ2z+qk5QiJmhURZoGpTNIi72HBnafcJgOuFNeIsv/ge0xa
OuVMDiNgpBGX9J41pfTm8l2PlxXhr+wH6PqntqBSiKBUf5xKQCgaQqSFzn14wmXWFLggow7FQ9PO
5iy43XxmrEOEXcrXblvOVQtOzIri1nHctYqdroXY1aMgOa5FTWfMlAg24J6/kHWsmn5Q7Zy9xjdH
ytQ59WTRRPmQ6QpWf2h3YqZBLufdYJyKKTv4oFyIcdUMV7k3ZJmAiOCH+Sy2JmjnrDgO/VDNf8Y1
8WZlsJPj5a3t/e50j+O/6UIiZay1fng0jcyVUpxEmKwownFKOqbW87Qczvyd+jAHFmgRPURjeSgG
7tFOTGsPybZLuzK6uSNp6gZXAs50FsHyvalAHVrJGca1pu2jb5ahvKi8Wr3sQvaih+nOmFpjAS02
P9HsDVEGmi06Ts8f4xAgldl6baM17se/duIg4UXJdeGtSeaJw1ltb3b7p+fsQ3ftS9LbiazE0kKt
Q4YIUWLLFMYGv6qjCxwu/nqYd2jPuYz7taczrZIN2LUzuxMEeXmKZPnRCdMLNqIyIzM3nnbtf8/7
VlX0rTzgKBfhIJ0pbdWBMD1Acn/IZ8arfwpg7uXSEMi4KousIUj8mr5nTLed/0pUHjpUAtv6RACc
TeuNves4PmObAcFRWsXeq49su4J961y1FK6RMk1hdEG/aB5JT2OVREX6vF12LdX76k33JawA2szp
jKeL3JgFtklIYGhYGzYiErxVns/EHCFWb/SpbAs66+AenF0QOj5Mot3epYewnCG+Uyu6WldoFxI0
tYrG/61HiINbtHnmnCB3S/MH2r8c2PZ1phhgW5sU1BtZaswmEZZ30UcCmXyRs8h6o1myzd5lMIWK
NWVs8cnODZhrLag12kQ2Dyyr7xjiB7PrcFueMTPw5FQTogQzKIpeyaT9OcG8875wMGQAxha8tmnj
J0vnvGkeghY2mXOYVmzCWefqP/sZz7HqhE2upU8Yhhkk/VGZjsYWREha2hE2oHQseDg5bmxhv1YK
ZPmP4DKcfvYXO4oxUL+ANHPYA3JAOybbTK1rGAuTEF477Wdl4o0Tt0XzaMfkAdmW6rIAM/I9HOuE
mNkfyzE3eRi9tBPN2lhnBzMOAdCUoSoF3SRchaGF3EwHCuKQSR4DGfnh69KtMi98csxDhWZt3Hhs
14FRrF1Rem2o8JKstv4qzlqcABoLXSIHdibxaC7G4q6JDgiidraw/5IqpY4cX+CHpAJZIXmIIS2S
aF9Z20WVVQi01n2qSPczEfvLz2TGW4SlK5FenmVuiJmdjcO4OmEF/FJWrvGxXErHl8YJkKOsDhxV
N+2oEhyaqTRpFBet9KsL2OuT6SzPD+040ksAqTV9lXN11vm+lIFQ4+aD4oYdo5vf4CT4h/ChRP6w
9I9/RoiOH2A+OS3CSVrZkcBCthU/gb3wC609T6QNAQC/UAGbMtIb66ABFH5elYn2GNV/LMXIHHHj
vzq7P7LSsWDI5+vdcTSXkYHTChbeZYhV7+n1el46xPW3qLXCws9TBmR0UTTWvKqv1AMCMO58jXxq
wWsXe5qq4WxmGVquO5xDY/bakUlMnmNC7QDQoraPIipnZzERUfTE5apI1XMzR1xhTm3miwsc3OxX
gP3ZsKakXOaf6Pp7ESPH2aOOZsWDnd/dPpKBwKbonlG5hfB3XvoT9ifiFOpPiIgePiJu+0FmaAPU
z5MhYGY7w0bxAuTpHWMka1qjZ7XKdOr+BRoepTm6764y1SCRU0120aGtsIffrbvn3iu8L269v6vZ
Edbqc0+r5/AWWRyViHNqCIG2sJ13e4iQAJvJDPup+zSxCGNRkty9eXciGXu2vG1sZkSntSozTBMd
7laYquVAgkbnuNVm5PSsB9VgfIOFVQnKUsKMnjXzEAvODetNoSeAC9jxqFWe2YlVezQAGVg/DDgj
XxbdYI7U4aNeU0tHNXBkre6Rd8CLq5bVzGYvfAtVxfN1v3h5VhT/rb/jNMxoH3yVgPnnxRLZCJjf
bWXWxxbD0iO0Dj0Fdqt5/g4EnPPjU7Ge0A6jC63Jl0ydsnG65AYFC1wmeO6rQ6K7ePDqhGeSRGKc
/7Xv0HXoueqcLdcljXr7bD3izU2Zp8g7LDoDijBf7B/W+1WLki1N10lSRrYALHCqSQm5SrfOeb3C
+HuQczkEFwT3YXyb6l0flnhaJ2m8ipQMM9IV4NhbbvyHRyEkfOPxJKd+UTZQK3RmBS6GCWJy9tiC
8dzn2WBymfB1YhduFCM3t8BFSZZ3ue40yFn8EBOtXgLpfFNfuhJg6h0xqR8g1Oz2zu0+QuIzGYAH
OpoiYV/PRPJaJJgTTPPwVAT/FaKGT6M9W9QPhKtHbsPP8o5215JidwEXm2DrMDbREOVAxzw5zFSZ
u2eKL/V72w6/cjh8C6WtVaYV8wazmvJCvanjgsOp/6SfoX8tHLlDDGTBYZRsOs0hiw5bvHmsOlIR
e6v7dheUS7HU9u4HBaKr5kmAfD8HGpiTf2/kYj7AgYrwAzta9I0O+K61h6RIRNyyxFLFReoLuy0C
lRyYVcpM4e1e/UfM7EUC3/H/h7IReIMR+Gd6/ffRaF3ydzNcMb+ftr6rvPPL/VGHCgOcfVNQFihT
Pdnlc+cyIqlC8RifF5oernqma5fvzhBY040OUrx7P5AzpYZiPE7Y8wYN46A0lv7jLlqzef68snLV
1EdwRD+z6ZM0/NRdTlLTwD6l/YmbWBBXIqOSKC86D22Za7OvY+Uf55icbVMcwz4Gc5GPf3tQJDqt
Gjm5TV5vntcEzQC/XT5RYqWIEP6gJ/3ElQtgvEdhDx5GZ3USu8aCQUAbFxVDKVsQnePDricefOyt
A4Gh2qYodODpeBcaD1vueWbVxVbL1S7Ix+eDfvnAfbW8COsnbdhtNzz9h4yCxL7h2Dibx58dTriS
5SdOXV7yGZNMGFk+xyUBpCfbP3peDCAsnqpDZ2uD63DNNjdTtLZC0Xqxds0WdebOIUc6g97u1dbc
OCRmVtwi1r2CZXFKh28EcR3vSNnpWvxafIzwGtb75ntblgs+yMEM0JreykRoZAzN97bKY6cW3AE3
GK5RlnqUwbnwxr8HuMvxlC+7CGvzzqkIyZvVQNIUjxqsWpKmpDr63s3rzruxKkkHipMH8/TXtSg5
f1f1ilkvdA6pZeGeL8w7oHMdOiWTVqxLe8egx33Ap19WqfL3AB21emltSlO3oMi9U0+2DDXyv2Ja
DTfMifbbGZIfJW7CgtjIw47QDcuYFyjdaU5luF1Z+uG27lBclnzGSvF8eMilIFg6dZYEVd0yBTo0
GoSQHr01YJd6nVxpFfNlHNWEhBaGptM1hTWqy1NOwPZKmLsJO4lHOsSFGTm0yYGbQLW3B5T0QnrV
BHHeHabQ9/dlJ415dIdAf/Ebm0j1AXCL2ZTsqkN+HLxBuyChR67KoY92EYQm7UG6nPIcj6qLYM6k
9kKUQqjfJcA09ev/Z144Y8B729S7f4ecMBfhN7Tz6rsZWU4J6zF5f6xWfEOE8bro6I/1oCp07E8E
+kGUECAHlHXP1Rh5LYP5goGnurh2fluX3RYZE3JkAHjPuy+IL7o6BEh5qLUqkiDn0UWMa1diAZ5u
+xasdmJDttNWTuFWxIKLgw1Bz8cdtivjx2447rfXhWsOOF7Z08wi6w2RPGkn/RoaAyXABMtPt7zN
1oSPAUA0WYK751jHo2t94OteClY9eyBCYHLzMWQa78Ve6ERo7PuGl/HedCfGCOG+4uSXPDdxCd7p
F0yBpkoU1AuJydXtFkFq3rW2qWpRjCvnVYCXVcf2EanUXxGjvB9ORofrdeBcP3exNp++P0kiMFvS
AcpTLKHPXbT62ESglGQDcmyuGfC0JZpo+lUn2mS/fITodU+8I1MKqzV9rmsmPwsrfDD5JU1C1sFy
ymfrV2q0WEfWgkt+zCz6fSOochQKL++tUFNr0De0QBWaW65y0QbfO+n4ErEMsG3XR4NJrSEE7dTD
snH+EIfAbeSv5lGeRsI/M1iiBRcQD2jkohD6bxOJWGpdPs6DYJZacrzPyIdqKM8UfRIMC/A8lGvU
R2KtkCf9kONeyZBWFQSRviOQF93pcsvfKekDlNRJSYdYr/QP/kg/3eUsm0nblJiHL1nheCCnPTDO
42M4ne5ZFpGOuz0rR6JwBxMVxFzzgOv58kU76X92XsKU4TywApxP2nbhlsjcmu24+GlgWn8NXUfX
mQ09kY3j+FpQvTswHE4Df57tB4PZ03SN6zDKaZY3RvNMDPORd3u/3QHsQF9XQq+wEwegIGvjU8Xy
Vvjm8uTx/NE56vSncHLdKfBdVroj4mahfp34ZCjKrFbXFvWurnBFgJKmZucBnt+7pRFF1TpOinfv
K5x6ADr8BySCfqviqd8xhsm3fIwVAWb7xl51BB7x5Qvt2PvWlagQwufuhCph8z9KY4Joa2ZfJvr6
EGRzRbVspnr3SJK5LgyYRcYIAUYoiyLylTyEJMiKizQ71f11Qs+zDcWN10lZI2MF+iGxYEDfYFL0
B183E2vmC57B2D42eHJV91QbcZwnIdBa/Xw8CGuRkaS4n6qOCXvqdoewAl1vPdMrigTugRu6RWQn
GD5hm03czqd10Q1+0Dl5BITVa1vmc44mrRZeprysP16++unxv+FOtjot/JTQ2UgPh3J80qfVHGmW
ptLDNOcq0FR+QFufgAhKfnOV1E5R66NybCK4o8p1XYwdZErhI6V8IIPWxDH9poTcQdNjXalnvuJC
rfkB90gBMZFgOKy2ZeCDaXnkUn4TtW1m8QpatHi5p5nMj7fh57KVp0kNg+44V1sR/iL/Vc030TFq
M6dP5MFhy+/6TrHR4lt1A35bYHHSjrv8SND8Y52GpU+3VFDlHsi4B1szpJlStmPmZSy/8ET1etCP
KM/aIx1gUdNe4+hbAxjQ741DaqiVWSzLekX0UGYOnvUrPQ7p15jzVPAvktwiD9yfVCmddXl67qT5
c5GZn2FVvxQodDnDewV0NBWHEzw9AkYNBcsxA6wAH1EFHyB2uGeizHG6PYBALrsmyUbPq5WSm89m
S0cAdAXibzChOsPWUNl4LgbOj8sNFeDkhQ+QSIZLTgycZdEjL+vRmH2/R5Xyyh8Wj+VSRVbcwgNY
wPY6SwasVvJXKe+wbTJB8bHflnvnIyv5poQCtU+nXDZXaN9GRJ2EfnsM9/SP3CXzFa9s5l3Gs0Hl
emtjdmKd2I9c3XzdrydZeS1vvVFM7XVs12BxPFo/MQ1qSm+6/DmR0w2t0ARlh5v7fiyzufHYumrV
rnhWTnQEtja3zoMoB/KCAW2TinqiMMw360fjPFEsQDSzfXZNgEnTeQA0nH4Mdi4lqUU78NLEsiKF
twq/S2tqnLGloxFG2vC+eMSDCo7j3/t9lBLt2esVuLM+XksCYAyTUsuCmJDYCZWBvZl3TtNM3N2x
pI3uY64X1FNHs5HTOmH83T/j9yiArJmTA6bZdt6LVR3mGoGDbvICPG75xz2s1+8u2Anbu5h7bMFx
xacF+GfkakVqudEuI3KNjyNCF+GDgmeAr94gpSEwsEYzcyQJ7SUVkn4dj3V/Ew6aQoxxoss1ZkaW
Mm9/AFw/7//0W++pta4YV5gp6EkFWiO6QbuMEdn+ZsMEPh/HHDc/Qmub/2QZfZCHKuanKK0vgQZV
cKLHl2pzSbaQfQvD1TuxKy8ljs19Ii9qYlAqFYtY+SCC+1kC6syZsPcOBQBCOze3oUeT6d5u7QfX
EHLxVhxc+fry7Oqd7I+Qe0sZN87PA9KXe8QbYRxtFh/2mMuzKYgznYUOT9guqUKgoTf0Kzqb9NR0
m8b30IGJ0vzkghBPQZhbvlGRWUssa/4V8Eq7uGldO2v6iUDDMNVW6kqQOCR0andeVQgXiTiIhRi5
d/wAzfUPtgbeZHucKi7UiBnQGug0kTAS1Z+7RWd7sSJNpq16oIo3oV4B5/rRzDjlATrKqUG/9fXr
z/c+7m8G3uLay0+E1QTBkACQmuzgN3xGfpDTro/COHt2g0EsB3klrd2TRD0ncnHHSpdcq9uFAPUE
Wvu7r599PuElgToPtqHmYn0w6qbPi7h6uZxXPbzoDif1P8fG8hFppyS5CgEvkQyr8JTyJzPDB9OL
48HRpRMrNrQ9ZL2Fgs3Giv275eUAQ6wj9TpPMf+e8K0yU1fDn2jB12PfZIBc+A/fia+F+Spr+EUE
DWvAgxe3cRkd74ETE8zHnX7yjdqrseiolXrCbfsNa4ux0hFfwbfJv7TVjy3uxRZqhtoGwsgzqsjC
m6XukYgfZFGPk3cQiF+4OnSGRV7dOLdTUFL2RHlFB/8dSxZIG0aCS70QJVxkrBrZpjOwMNUBl0NW
SeopxS8GRK8k8D8FjQ8RzvmJA7r4AH8XBzGmFfHYueIiWRpzKsK5n+4tNY9rVWwF0BSASg1yacKE
Ry5tptCAqxkNkRkN7N3/xOz7HMEZRUQdJcNbN82gJPNZVEZNbjuEhn4i4OOjJDnVy7R7wPZYVHSE
84DxhZsC1bdwnWNxG5nwb1GsdASxn/reLGSKY1za5qEwvPzGUN73TgutTgCLZx9lurAdd3+hrdx1
uEasAubVgLoFKHer4F3RyWTe0rvjJVeWtVf50r1VG2CFFzcrZjFfH9z95WqWUBe2Bh6sBL1W5jfi
xQbS06GXjF3qMufkAslWr5qVLD2rBY74+J54kFMAmU4w83wS/61KPNL2bIeO48k1ghPH6GjFBhmB
R84vIrfs/Lp2AD08axX9SC+FEo6EqId590POi6gLgePI+D52b+H+jbLKCbn99ktl4po9P5iFymZX
D0CSlSvkDT6Y7KdBJKvDhLjE8LBtgIMiz60HfgH83zLLhw0Igl5NAg7iRD+0c+f/gdvFAqqzMovp
DR9fTsrCmDivHTP8MIp/26mMZljrTJOcH+LgRwNpUFEpe7JGCSicgC1/sPACYIt+q28IqRG9R22j
t2m7z1j1L+BN53RfP1HyH73+7ihHIeUhVrC9etgSwlA0XZRiE0wWia12YbuUdMJOsnQJ3eh1LmIk
GqSHa/rPiQfjOSLgO6TeGvUeXQbyLUUVbjEWq+z5n/bzJC0IBaieecccBU5vkAr9nce7veEClWNp
egsj8ezfERQZAeuyObnhtamjMnbEFoV5VK7HFDVsbLb/HnIUpUdzmD7oU0eqsisPP+PI5sEpT6ps
kqJLu0bVgqGcJa4xzz1wYK/E1KU1FhNBlN7QrUZfxtTzJIcjhdOVxwDAss/4CUd5XnueTWS35WuS
rgp9YQPmicWaiVzaCJ1zchq6ZWnj7UbV4b4yFZY+F4Tkj7YJ8le8ydiKyHuSV3M4UUFD8sOd297y
4vx5rRWvcDMtQhgID4HxmuN193oWd+SEfkEPz3W72TxG8q0mYBAKCXN5hd0ygAaRlx98sgZYi3DG
IJRVg3YetVEBwYacwRlkJu6jydiQPdkXAYZPqzSIau70e6Hq4CucIuN8zggKFe+nQ6SGsCjSDA9u
OJDygL8Nc+7BDeoGiBqaiexf5onys5/T0HFrOHd2WomyYdJyH2AkEXHnKYQlwfaEcpfI41mQlGLk
T1mdWaZ9C+uq7RYUPQzPvgiYsRdXp6iZGFG03w3g8nQ3BXo1LGpwv6zzYqoXHlawEUN9GyBIo236
RwBGeS1lguNRPt2p2rwIAdg1t1ZNKPCGjz+kGa04Vd6sMfjFNutrgYQY1Bp6dioSLn0YpIsfUznD
QMnm9a13geAMnZmhIME52ScPc6FUN/0+/yGaxczuPPNNlJHp4iCO1yVxDT14ew2KX701JroddrXb
Ti5LwpIsSQ9DZutOxP9RuWpo5TpIln2/rxtNPKMr7eR+o0Pxzu5XTD02E1cBZGVDnaDohSCSqB5c
SbR84I8lmlGVKwtor2a5b3d7IO7NtRxStF161wiT3SPTXNq+Y5UT+L6i9BG6Qh3nZbhxWF35GzaL
KKGB6SFXzLnavuDbTWnIYwPOegHtdLv81u4MbOPcyGMKHinXQmC/DFMuNAPDLoKsyyB369NAe1jb
aFbNHMGQTpUHwipLyiqzYj8bSzXbVlqVHF3GEOZv4/M2IuFZ0X1Sm48zA+XUEO5l/7KwI/Vjz+ry
woYDL49Ner0b98rAbvwuuSBYDqt+Ic5yCbFtoJ0vS7/rMDHazTzf0WmvVSOsp6mw0vRITHLAF4KJ
n6Zy2LRlFvo4bhLaA9iW1H0gR8Sx1po6ZWX0/IosXESyOIhByi2AhGn9bEalVK+xJC3YszTN1pkV
C2WYathxpX8/fSLhNVhZINrwk3A2kSsXK/wAJ9zpHF/jRd6kVoqf2HX/2oy1NLuRonmmFmpxebjF
wzQ9hmDESjIrcUdkS9LbnigNy7133YFQ3swdSaiJRcNvYhI6pn3GB3HQAPKMqX2b/QztrhjAjVBl
WYdtkWVc5mkrul17pBEAqn7LpVgq5QaevjRCqPQ2tFk+HhuPItLWqWyEdwJUgB4GzWJWm2xYQT6M
nWTj2K2uMJj6UF8p88hBXEgpzBCesoMlKj67mx6Mq0yEc3mw6eHjSWl2DX0owNvoY2zcIyw+/V+z
u2EHlWuPyAtE5noQMwbxu/rlgfKQYoWM8f4u1hVc2aqpjVxDj6Jm6rVhrPW/EMMbESszliSfWv5g
WwfEtXQvIMvGV09edPMO97uICugmPZKNi7Yxrhq48q0rTG18RaUuZH7zDuMfsg2LlCrIW2PizEwj
YP/Gj9GEt9GJ4CGnKDF4Xq70Y6FJuJ278Wub7TAWS0dcjF+1EaSq/BpwDKK4S9WK42W2Sv/YARCO
9sKA8E95mCxuCf+70XXKqAvZhrpvW+9tZ8i94yhm/QC6kBpwGWEhxGmOo/eBQUixU4ggEXqckMdK
IQjJu1TsCAG4lO0YH8PHfB8UYJvhdYEDBEfNkV9Vzd6sDBqoJuJyVbmqhbngmxD0DFcdUedYo7tf
Hzh8BShrem8ECmP+b88jK6v9cTBpOMTArOmWszXGKz34zWeJTzc29ZYwjCA7HjAX2NucOLZhNwR/
XjdgfuZudbz3Bc7935O4KyE5R6pyijohlrOSUay8EPJZhmKGoWwPaxtn4DdArP7Sd67CMfe5HAbL
lG8yLYDW3uJp+ujPc1OGzOhX7TbyFXdCZZ1e20ol4JPBoLMaZlBEHTgutEWEnhdnh1cKsFAK/sEi
/wYINpHpRRY6z3CR896+n95D0hLz1rVkw77jzFZLpEdMO+9Ikwavyv9Jdqq/3c+54fjmkNT2fflT
Su3byhMQJ0eZluta/kHgiSxqH69boEQpJsYYw+0CTdgyPafSxFMGEV2Jqwo+1UmnuExCLVraGO26
TeyoTiLpKTp4iz3u/U7q1+0fK8JQvSzF6iv2FEMAbC/zXFTEPz5JlPDuxb5+06dVP4HyplD4yHCz
2zcyixzBVSrj2BlzlnUIbNhk7gZ2643UMLZBbpQgudRfh45YC6q3hzp8F8E/k3a1DjuVAsJfdRsc
aOeI4Ty3NGIIlpd8P5r871z9hUPpyZ6EsYhpeRqIIDVnH10fJIUGu/BVhPIvq7cS70vKgoAec6IF
pect2J9FinZeiE5w9Naay08aADHa5lMpCAMUrDb9KXBn0qp3WsM96ckr9R9pCzDqkoxjYxDopGJg
mn6ATlfYt1pbk1Xts43xDmVBJXzoqLQQxsD6KOImRYAW7oaGZJ3IaD538ri0laUdiko9/LH049Yw
x0qzpOjOgOqcexdyjrbq6xqIs9wjkMKN3fX+Lk6iBwqjOG6W4xylJUz3JcHTRdKa/va/u+XWz7b8
4bNWIjSYts7OudZTvqfBhu2WVNbnLJ7lGsgRcsW2ZHXsGF5wyu5c4iF8x/Zeu27BLRlaM3dILIgz
klH8MjqZhjYbF0QWqa77tCIyyfph081ZkvEG4AQx6uG1rnmpib0uygl4GDdH2qvOibvcEb5sK1j8
li+1Osm8atLBojF9j52KSLy202FV52RAom/+qL3UFuHaid3wIHCZXz3TW2H0hPXiHfqtACAQpeg/
ER/TsJKEK9m7EO5kBLvOe7g2Tkppu5CJTJkYkAPpgzB5Da/DQekuJtCCv/Ytyp18Wq8Qat9XFJxw
jLWe6McNTEvb8aVq+PdI+7YmpDSaQQe2Lm/qdUsIEgWnqoZqb9sTr84fGhEFj5igtnbm91+nzPcv
z/V+nBpt4/viGubKQ2KE+rvRU5tgoLhzcRFp+JrrPuRVVmO73hOn67iumcY4+mg3sIqclz8nsxMY
DshE19pMOUTr18R2YcJmfrShF66AwEchBWgA9r9jx+JViVwkKN7y5Z3hUnBOwzroW4VU7OG22Kvp
bY/YXqo3lCpYKZZvCWxIt4yPz2f3Xz4wfhdFKXYBJGg6IdJlnLGOZL57lqA/5WrJXcnTSxoZF//J
uRbeu9V9N3tD8sCd+IoqjVOnTMuE6Pe5DivbjPBjUnP/Fq18nQy27DO/ZcmDOgLJDl1LMBtQJut9
yBFk/9WEQvbQ/KCwDNIZuQRd31v6tv+VPKyUFhlIyj9kNDzPExtqn/LzKIsAP+iO9cX5JLc5MENZ
pvyxWyaFHajfWpNaUAmH4cNebRhHI56ODa8F91pxJdijpJZVvbfwxwDAyAVWsxa0o47jyVthPE22
8UDa0u9ItgxgimPxJlEyjPp5gtaAh6KM65QVJa+NO61Zxws6BEAk1ov7MvOw95aDdakXbu+GecpT
HDZgzw+zsqj3BG35Rw4FHEQzBKdojI7VtJJwtTCvWCgEETABSpdPqzl25ASe/osEDX3txIQXhE48
SEPB0fRqCG1iwKXw7QMMWclh/3g5tGSw4G5lgbXCtKO9xjSukCNPwGRhZA0+dGDi8WkqQvylj/IK
RJUczSUNZJRLZQ1Uup2g3bSH07bspK6Ju7H+/Ip8QtpDLxc3nzZYwAVVupJqwLGYqeVPThtsDeL4
12j/OJLlfkBGKWgy/Y2vTimvW72njUU6/mx3+2aT2FS+VnMMm3tyct6eraYUJFbxq7VcI1UeArNn
zhwykGhtEdUR4lvZ0eOTFqDlIvfDSDIw5eXCnT/ge2bH3TpmSZvFfN2IvwFvi3KU5prKcU/1ktcc
mHBQ0gi1HLoHLhXq6K0PwKhiym/Gs12maaEwmzLogxkuTTloLOxUBYZA307zYIYiYw2ahkmviJU3
XrBODkG9MUAQQDqryRWtkQsw3J+kfFV9ahXxZtlFMRQ6eUc6u/mP8WKBmgBte+36nGFkZRgwAP27
Qf4egkNsYwXUoa1HNQqmx9+o+jiMtT17XnxC85st/QqY/XF1i4fdSFjW3heTLIjqA8iIxla4C3JF
aU5C3TuCQC7eP7MIsQAYb/s7IBaZsCeEwpxwriUsvwJM77KaCfyEokY81YYFdsjdBB1PkoyH82e7
AmoAn9FyKFgvPapxJtz/a10CD9waDwYcWpn/ryDchSCT5vEvhQr+br4PB7sC4VNCnKT5PG9NkQSo
i45oU+nBSRZXOmv9AZythem7bHA3W2Lp7J4IUUCVw/3JUwZh1Fz/XuYRnWg3urftILB/Kp7o3dcb
7mHf9aCojguj4/lZlb+RakQsYCphWfscyf6CUtNn3xuaCmrb7C7UTKv+Y/q5ubxPANmyOkyvstKw
cXQMse7MKGHyiPzaji0SCo9SZuzkcmyl4Gx0P/nXfo7epfabAe50gADHeYm5qhAKWj1o88jWk2wl
7BxC/M9A9NnYnOTfN96Ntwu0tq4YXwSYTeIRkDqg6QbyPllTCnO6gRfIsV6yJRC7eq3mhfq8yC1T
O9D52mWGyzmeMHH0r+xPRFe8Iy+4USKIePxQjMoY/Pm05JFZVYke72uKiiZ5A7AE2I8I0T5ooOXD
U3CSKVn6s3ywYg/cRSOZsTZSoTHvV4KaMrDDtMVvsJTxKW9oBKEEIrAE1nUrw/HkUoj4ebUMfo4H
1jmbKmxX9fqLy6FoUXRn4lT63Zp9DCH/ALGwpFLvsLaLfYj5jQBPdQ7r/w+2kwyS88vZHR9qv2MC
5SBSXjBh20mhv9xcu8q/OMpInDixxHCLDIkwQ3XqzdXa9+EFJG2tG8GO+au4ehtlTt+4dJH2Olde
NPBeiA/DPZkllAxf+6SNaFhaWYVcBD3MPWqGWuLBoC7xHBAPEyHrmQVILgAhJ2Zb2UsWyxUZ1aP6
lBfOgvIHiKQ384jOxNf5ugcZIA6T8Tc0Ks80mjChP1+aPh+ZypFL1Ld5/I844tS/h+FVNp9R1YNj
PR2Q+vEig6lnlspxRquEWoGAi/TbOjowCsYyYDJczwdwoptNXVcp7ajJQyU98KJCPD3zwhBDcvgH
pCgC5d3aqtBoZRZavUc3g1XPJEq1jZLgJRDv5effUcxujm+cEawDdBNrPJHyAUDJPY3MhQcfdQJ8
2w17x5EKo6AvYQnimnJXhbQGuOq23to+aPKQNZ6a8BYUjSG87HsICqatm7+igOaqt102MmUEhd24
CN9qlhILUlPyRkcdi8aP0Ti5wOLGoyeZQMzNVQEQPZU2MSyCt09cP6ScD8M3UqFcLSdHudij+hdo
jUKQN9ZsQQ4tAky9MxjVmjAwlZpI0Kd2zCEQV64hIFnviZ8S491H0KfZYS+DshHop7N2TjXz9h9a
dUH/j/Yu0i/gKQyyd+1l3Pc2hs7cxQy8T/fO0xE0ao3CatJuJ/Ye2jVwzD/iuJoPNq/k6fRx5Bx9
SElzoAJDwi2b/ew57+gLHtUw8uNpnITJVAODRK2uhAVX1vpEE7CLQUNZ9luYAC/utbNB4KMzynA3
FTC4A6B/1DxlZIze09qzU8LpjlL8Q9+HVtgpkoBjnboqIX13BDBGCuF7cfOoSo5pmmiRyI3MTxzE
Z6Cq/j7MCpJh3cUxHKbNgIvAG38wzmopXW/ABg0iqdfvxTgt7aXY4fo4OV5DCmRqzOBSWiXIZkAo
IxTaXD1Rgii6c0i0ErHL5WHsZjTDzJFKf3JHWDdx7qc2QqGWaCYcf7h4lB4ghEWa/meipLPaFXV4
Xn0psTRHd1Nu+oziIQRIqvoc4wuz+7iK7R5ieLUUQuUdATbIy19ZP0m6gbYP99amDPb+FFsFyjb2
BjTcq3a+Fr89TufQGefSJl1dED1aLnNh0swwayvv38itFmua8Ocjh7hrOVw3bEskl3V9y59Cu8NX
URHnZZ9vWH22o3j47YRc6Q7U1zl5PNXaK9y6AqpJ7Yvmg4i1xK8WJpx+TyI8EBOzmw+KGg2V7Rqq
bC5/bXZ2D7hSvyoi0EGFt/m/OHLxDtKVbDCvaPhXa8fHX84AX1TyFKwwXf7jq9CgnfOjJtgdjVhf
2JBAa7MQpfJbwA3b01f867OzhS/KVAp99/LWhl1o5zeFUNiMHVcLA0uQ6Wp+J9gpHlvtP7O8yFAZ
mqyJ4ryhYzN1iO+ZDnbqb6/FtxifZYGY/chQ4HD8sQoTaVGg2MNKIwn+rvSB9njxVUjuxy/kpMqM
SzNvRuPQAas+g2RpDFHLA+ApcJeXzQeuagchQ1zqPFxGYaTHkOgvTB65iqoDZGy5ij1FYCzE70+q
pq7QyBH41mPtlQTjNHbALvG9NBMX2HJlc3G4Y7XSglPz52hiKxZY2d/Kl25aSSbN1EQXhD6WymC+
LIlgXeiJSnN0BFymhCwmfiJp2YfDUjCTgqwT99HZLeJVFK9BOn4oEFIFHEjTq6EW2KspIVy/V1Sv
qiU+fvnJxdkxKY1wUJDSlglgUvWyb/XxzHgcjXwTLXuBX5v9OQZ6GgGMWD99x4Uf04ntwYWpQVx7
Y6EGyM6vuoD0xAtS0r/BZ8vv9dEGaLFPNYGDDXU4+QrguzRHI35U8uf+mWz4vwDF9tGMO2pUzSGn
yJg+7Z4xPe4t2455h6YSNbbSxYGYpBIslEgZrQthC67vgKI1YNcb5ziiWYIvHb4JSdhBrBRdqGGk
fOMgucx9o+9skTewXgsaqHBR6WurARn8ULazAvXDuF3jsAit7B0mpytJCkwb22eo1s/TxyX9INjc
nweufc/C/c0p+G4/J8IHD/9tTsl5vQojKQj+8ghHF0rvI6Ng7GSGUU8V4Scb1GzcA8M4OaPAdH6L
KWD3wvZ0CPtPX3VsIZhcDSNeDDjcubPZdUNfikMv2Xob/9PHF0CPyeha5eghAHpL0asE7oKg2yjP
0T5RR1897MmeveY6u3gSJSmrRA0F40+wGa+Kc+PB0CGtSmYC3i7uX84LtXPvDPzzCBb0loutzXKy
MfkLT8NzC7lDFxL6X76Pdv98ZD6LrlvMmtS0gMfFPyJG/uBLMNCuca0Fp7/cW9wUmROsY8eyVsTL
vELvvUqqR2pFr0VfWTrOmg4lFo+YbqlF2KfSSfunNBsv8DbcGGY2udnz439j5S27U6li7JWez1mz
f/IyjSKEsbW7CiZVpy7jpRKHyRTl6mGcnOJllZwsaiJ5ExUievMooUMixjx0wXsrRb5s+/QgAcHL
V/tNLx2zTger0ktdahcjRM+1Hlb2FncYqgF/jh1K2d2IjFiavUbaxbLpYtkeq+Tl3m7Ib/yUpTdZ
QFSEFfJJCS+vxI4ZNthpCznvIxzaAW+elFYngUEfT04cf0TcWvZ2fCrXENdXfde8UBZcY1KVXtu+
M1GWCMMqg8szF/3Zae1h8e1LgzvaIc7IuCeGqTgyXJPRG1aZ6XvEoe935quV0gUH0LwZw+xhjj2W
/m/4pseCgsLvuyqkUKVvNrZSMDX/I/zxuwWNePYTGBRRcBo7q9lskSEE7RSlxceLX2She0zlf8/V
Eof93fqPrPriNJKb5J64Y4tfrDvSmdw5z4UN8BhWY7IG+npe6V0IL8gObvuABedUmoSyDH3V7Zzz
skyS2LtKViT7ukkgVxVCVDnGRPfbUjh7yGDXaU7u+fnCqVWc2ebJifvP0Eu9YosiB+K/nIcwLcnk
HkAGw1EEuvkm+AdaZB5NFJesQjleXpkd5ppjti4vceBpZH6nMF2kJ8qNx2NyR3OJFlB1noZaZjeT
VROAiZ1n9OukCm4i/eEnuIWATHxnieqb0r5F34gbdgQaDQn5bAdNYOe8dZvQh4MoiK7QsiJlADpq
BG3nlll1dAJvqYPub+HCeIKnKjLghnWTSx4tyuqa4aeGvqw/ra4mUWGG2RAgwJsyh+I7KBNA92nW
+yM8TVdJB+QJZK6iCdAmJensxFHhX0xBcAY6vqyOAAWGSeqiLBjlM4ZYuKneqFXIfOanx7b5TwSo
vv0l+YBleYMGGJgvAo/zq7mezaVx68ukEeVifhhc5EkS+RZLdSMZGTdahW2f/6mjWIv1acbfFcNh
gmKy06pGP1+Nlx4kPcwGIPtn9pDDdWRGJXC535gzQ++xkytyKSd+2YpPcJEYN89bG+e7zcOtKDRx
b36Oue8IuzvDoF/sAlquIIjq7488SGFc+9h2xP7Kxc0Px2lGwaeNPNYCWsAL3KgXijDezWY6BUZp
rw+PEmpoQwcoDA23u8V2PiInAdNC6mEurGkEXrTHUGagsrHFZjEUSZZvtzb9HLu9BBYiObdlxpkh
CSNih9lh25tXuWOyRpPOAozC1s5AewaXFWO6mxEZkqTZR/fSvI8tlKotdVqqxk3nAGU358AUwbQd
IfGVJE9Cz2PGPlak33EuZ07LP6GHyAOdl0qyK3xexO5F3G+vwBfCImf2Gz7NR5D/PR9T9HInfWaJ
M6gW7PqCX8AfUetccgLWTq+0Xo6v7DhAVYGJuV9cpEWvqYuHOuKUqqauw4uUu2bqD+bJknKbS7gs
2UG6ohfr2LNQmUC5+K/TgthE0oZp07fSREJ9LQ+WMvUDF1Q8bVjU+0VK4XXS6B42F7L00WFkv35u
J+SJKd/EWh4ea2gET3DMzAvYX0vTr6VkYlfkCjVilYNZfvk5JX53c4FqAZNCpbWfZHjoGhcc8V49
GxKbKXJ372idvJmnxFXN5/E2vgpNS5c0jz0trDd9GYI50RXsoqcbOevYsdsijLM6nMxYPYZW5eQB
RMLqjHyD0buS0BqkbBE5vELK23DDAfSsCBQvWoDS/CrpDBfLeeiFgy1a2d28Z5e6b2YlFZzQ4b0R
g0bI7KUtWY6FpJ3d6bSI9fbu1+fD0XVgaVpLSdseKOEi0EmKztxgl2yJBTNmIABi1yyeN+jBiJsm
GqyAEcwiSOrWU61RPjDVmyil++4TFuxQPhpo1b527iTsc7ktXGRA08HNYrMUnbjJQ/cz7oKdsauW
RB5V4R6zM17/r60gjRnvNLFk6es/8sY28ywhPcDPw67M/+SH+rUkORoy39bg3fU5N0kBCvFAWkW+
rXVtSGnvMTU1hhP+B1DE+gNfyniKnp6borFymC1z4WQF6mZSuPIByLkTxBz1zrf9W/nF4G+0zEQc
47CvxDE+e6XPJJ/5XnDOKCnQpBCw0Sh59e6IkQXQ9B2/UMbLujGj7/AUQu+/4Mis/gLLkF2SFgNU
Yx9ZfecDNHb6Vy5iD9HCkRIdT9K5mQXEbm5txH36wQDBUlAu4L0B0OcK0JRpzupCtDjB5b2ngkEf
t06Hi/LM9IZa5vkh9wbVvScmZieiKMVzBdlyvo/aEJ88y1AQEPpdQYe7k9Z6LBYvrkBei7XJwnaE
DOw6IvLI1Qxmsm/smSHo4Z7VX3ius/QcjQV3Thef5MqWo/NXGtA4qoxAaZ+HHpS2gtqx2gG29+ro
BHesjbLZ4LcdIXg74pmDR1Es5ODfxrP2z9EsSLUU2muNyPnTpI9aty2Y/CFZCJNqOvYWAf9Iu9v5
NREWE0/kdHxwkeGlkCt3uVgVrvqPuzEKPY7jrbXepi+ADwVK59ueujQaHD2P7wxzk+9ZJaNySP+v
wBaleH07lIHGgDzgAUrB2BwelsFjIf3sdESp8ccCGWJUEWXaXlG66PZ29Y64RvfkZ15jeZbMbG6O
ngivlcwPhkmAzHUYltqFXn77Y0QQWYYljp3fgpuw50vyUbcZc5YmSgmFEB4KHf2/nvQoaZmoDz3/
vy5ir+4jKp0YxuHSD7eKFvNcQSMTl3TMLL3Z2fFGmShYG4/Loo9KMbONjFrgKG7zZRdqbyriQfax
bwCpPbLfqEicO9Yt8R6OlQr/ux+cmB1JdUQoWROh7qJBPAWxFZsSa6CMLP0CVK8vTj0CXQKD1D0J
Ezht+5HcEhMIhWn29Jvr/f/R4NZ33NF5uMg5dl/BnqKR+I/nKjfr4ZMf0BN0hDpOs2zFqDC6oCI6
mlB38qpuCu/4VslTtNDJjOxY+suzICvLG852ULQQ+GqUCZSnsrQc3Ei2vHKhtV1GjsAtrjDHEUk/
WCFnNM5/vl4lkLiGYefLKZK+T5AzZi3tNwsw17YiCKcXnlrMBc+nd6kzRQtODKZtkP/iE3FjJAYN
UN6PU7jDbEiPl6DuWUXPlhR9mncZPoQGFhPNZ1PHBCxSh942+ESKHFSdqJhbPfF4ureEpw/oqnKv
teq3Zk3KW0pVyxoVZG0skKC0xMJDsCI1ZJFnN7n+oMYKxt5u+LVibeDGWtPfOXDOoDlfW3W/5NFM
wgsya4JAbdjocxIb+tkbIo6mK363dgysceZZIJ2Y6KtJf43BPDohvOZtJyH4v9Lz1WJ/Io6OL/H1
a/JdDR/lCXy6r1MzUQv0XCIMPGhZB37mCRxYhLF0LUWK3sjJj41m8mfhhtJFx52xlT5ih6/iOyuS
ALjcP669ukmlcO8N6ILRsXxELAr1bfExwfbn73GUU+GhG0b0PcaMiBX9IMogsBotc/eQOZp9V88w
+g3xezkTevta3BZ9u7eVDTt4dL+vDTftGtu9n54xH+1hnACdXzCr7ZhcYtPK0QhODnSSz469b6n6
ci9cp4qAaNH7wTWFjjHJwGlMcwIWepGHoYAVAPbI4EFs3Tz7yflIC42peENbrvI2AMC/HJsf27f1
FZYiWdRRhs72Qv+a5XppvGB10WEmY+mysL1kfGeLde3HuJVqMAFf2oVsQ/ryw4Giip7/qDiR4XtD
M7D6ANJKG9lMG1Cm2K1XQSxqEdFokRQUjMkyck7UoFX0240GajKwHGpJBACQTL7WUSno/KCkPVJX
SO6QZI2C2uVp0BGCOkb/EtyaOQzUyuLvvbz2vuSxc/oVuNEjWCWJ41TCme4AqIJRoqIw2mQKVKi/
LtPzSdvT/bmMT/193207+YV2XIQstJMGb9SWKdtqkyYH26KoowD3XKPJ+hQYsshE/holrzlTQMdb
WpNRFAPpEWyg0OVmZypGmmMiPx/cwhPt4HYqn/Tzd755IY/Ef4brd/+Hm5XF4QVW5oM8MI3/qJHc
LUjjdePkbJoyop+U7A5RhidWTuAMqmqF1NnsUADCKrvqs/df/WWcS6paccvx5PnuPJYpUKpbalip
CsYv1kCv7E9OZ/fW3/BCCff6G1bVBHoaibTHqNkMACdbqW9yFAHF4lBzf4JTg2DDd3E5eSMN5MoZ
Uk7D0/BZzgOcLOfywDyRxo5bK7a9IMRIFM1/6cl3ay/jB8A0vtXvl+FOduGusVv1Yh3dQkvljfdU
MXnPl2jikzDnrh2Y/eBI61Eh0r52ob7O8qTGVu/hfzCD9K/IsufpiVwKIO1drN8tnjUoPBHIwmd7
fgg0oUVphoEULk07GnE3L5laGTO1OZFIn6Nc8S3tlH60/PMyYCpK+XJf0pfORPPLME8XaIyIqP7R
oMQ6gjIFHHcQao7SEcbZkGSukSAHjQ43D1WhDdEGgE0npC6pqDOS800dUaQ0goW4Mes9ObfNOX8Q
ah50PZL2nMsRP/NpDQd276BQg0FOnxolHE0HhB9Cgm1vf7CRU8biYr1ejqzz66k2yWNtNCC8jK9S
BPpiCFk1w8pYqWA3v7k/3m/FlYVhWzn1I8xa680bCTZPqYQLpKqvr9BNJxyAeT0X2UHLRtbsgN/R
W5eIWrfiSxRHM9Fwy7MxfRPeMe0bU66t5PVXl6C+qPkauB3WPZfsqhWOkoScCvr4caUHDRzzDI0C
wxyJwTBKobygXrPiIcX8HTJ5zKDlhA0MpR4QyaigfCUKY8i0zQ/v2RHrunHkCPrzq+/igGzUPcuK
MaXTzkNTSYezzk7/alnqF8QZUfIHu9DkutK0XJPDOvaxxX6C7K9KcjSXqBUBPSepLgA239BielaK
cLTXDujYHdw0RL4EsEqHval1mmcuULH5bc/dG000hx7UG5Omtv6DDyZXkWmCeKnIH4cT2Ui8vdfQ
DcAy9R1EvsPXqh59Y2w6/6tc5zcD1gsO2k789ChIJIntD5R/9gdNP3akrM/H76zsGrbHuLfbg84I
SAiBiq4AsG9pNqykaREoCgMyYzJs3EUsmDH49bQ2fl7vkY1W62MzXfyF8x+ibZ6gQdpt+8mENZ2j
RdkGlglcRldgJfHHM2N97+V958Ks9VX7ZEq4pf8jf5Dd6piar8VF/O+VkrFngcfrBMBmo8VZ//AS
1r0QuTTxUnThiTJiY4fRvlfnROuOsk3xAwzKJBaDChbzMc5Ia6RnOQtfP7bWQ+tj62OV0Hw3zjcX
fY06b9TkGkE8q7JYzEYaXv4rUjrgbudrhPVLX16pmxi3tcPI0ycbgxiUwFeBsABsFludrFWY1Eff
YI4+4B1cEe93mVmeFcbHA+Fz8/f/ytP219qU/t6Ff40YHFckhYb5WBJJPogOwYgSTMyAuIUObBPQ
0yJMEg8J660V5W1jzyRRvfzfzreA4JWYtG1X71fs8a/6/+CmXf26i+uNcY5BjfojJ83CV7VUDqAU
bVqF4KuZ2jO1u7qk8wJFhExiRVTWSq7eWobt/03jfSErm5iS69NBAus0LtmtFWRumdPi7iqZSgjI
Auy3ot4GSI7OkO3YRUuFkyceakVWq3Socn41/MHsrw6b6aKP6ltD+gBsB+2btmwdqA1yolVsVVTy
WBbGA7WHNDG6AMX2cif9Zj6FtMwUq7Q0u+jH/ATxrVfN7/g2IwqRzJIqDO0FsCLq5ndY+mLg6NEl
Fjd0odpyAkIFsSYfcsP2FFjOVzPjO/H8C7nNUOursRQlGtg/nBo+t4l9qELgGS6iOwb3wjw5m0c/
+5Ou5Ng+i2aEMbHrnBBIykfcyB4Rk1W/eOF320WIoxvY3XsO1zl4OjcIBjBwTrZIZeoJa7OdFtS1
0tlJJq2NF+R2cbFvFzfJIOfajeaYTEVCg5EY4eavCbBIjNWOmVolsANZ1KnOjAmW7GiBrBmsZUNV
TLZZPYegTAuwgLWfQ6gtvrrRlfrnJMV5WPR4jUSGNb0ekJqTg+0/sPNwFkqoCj+CS4uwgXoF0Qkx
c53m1z2LwnacqRFxBnjfhBUdYWdkxrblKHmlkIGOj4NsE1Eqt8/WTI98VjaAdEe+qTrUkT5HgFyF
Sqff+Z4/qfEi8krZfXOcyZJfwGf+y+HsIG1QxeJ1PEOdUszees5LGdoRUngxh4Ll/aWBysPX8/9D
chXhaYqJHzN9O+Fi21Z5+Tzmh+eIeplk5YAM+SRrliQGhLTfTX6TDd+lxmIRZx8QCMhj93EONT9B
UN1VFSfkIZ0Vxt/pJxNFLA4vaBoALCEnMbLKFV2KpgkAeOg828DkCOlNLGrgLdlgjY2X5N0D7MLD
7k/rYXHjZOezTQwVKhEeAuCgdWCUJQIeKh/xz61ZMmSzg/0Bw2Jdu2r87iQzw7hhvcq4CJl4rqDx
ktsPw9CGiYAZPnXCTSNI0qSmUPnwP7+F3ynC+waaAexEZG5rrqaNHqMEH6L7pxvTSxaHa31raqWs
EcoHZvU7xklOcwxYG0l7rnQ4xULDBGQnas06icQcy4jX5QVzxK1XwpFPbS3BLCOhemZZ4AWPopog
9FdM3RxWADNVodYBAtvlDQxLtdsyWE0+yUMds8xuCdCK7SJJOG3M/nFsHPVX4M3inzh4GsJq3UEg
zPLnlFrfR7ZaLZbihhMxYdMWCA4mS2+bVgkMNcmlx3Ho12UcvjwKfJg/DaAH2Q6voTpJqG0wdqJT
eR84ZPs2GBbe453du/4OhEUxLVWrUUq5jzOCKS3xCWMOd4K2O0pvWIatRPYMkMny3T5x9TcAPgsX
mWMESkt6tTzhUVIoxqJtZ1Nn3AtRyl0t6sV6jjbotOUWT4jH5f3s9RI7aJ05mbiQ8fZJZLxZGl3q
Wn5HoheDXRqSEas5jnZ5uij1AQ1q+dDhAXupB6kLbH7NBBbq2aVKjqoN7S0xl4h2+8YpqYWMTtRF
mNdLN7CTDC6x4g4Fy/QGJgL7yQMCz0regQMY1v9UO0wwuP9wnDhHal6bYVx7OOEqT8BsFTFF/WWT
8YNTaamEihzf3TUbTOQggVPKVU+uuvNZK4DO72mPKsfmpsur0qj/v1UQijc0UB1TCsEGEO7dmyGA
KSruhTC9FE1rP8XincH+e2uj8qLP82+2ItcY/pIrZV1NKsW6bzT+UOwRUbOikysEXn8PAkyhrtK/
od1UTxPltRXj8+Xz13p/Om7b6r1g97vIjvh8jVeVmTkYDEHWrYJYjlRJb3FSHGtIjevGGHbuDz9v
vjwqdZ1Or88JDi6toEDc8wMb3yr2VjnW+8Hw1IRlxLmjJt2YpFe3VBdoKzTig8QwQk3dPPZ+m8Dm
tqTtwhJRaQ+H2ilUfa9Woeg5/di98E8mxiIpgrvXRxeTSwTbJBNFrbvadGcgXk0kucBa//16VeFm
FkXSmIer0FRh+OBj1oenTVYuCilC7AhR1WCyvg1L/ehh5R6R0UDnbHlCZbXQy56IQ/P/SHZR5cMD
RZXjoUNuJN/zEgIYosHHIeCU61cCjz+3ieIL4sudALA3qv5lZtSgjTR0derxLUIWWOmIPQleFoC7
wo+kaAAQe7fVtEzqZWUGRZ5Eoz8ZKgB2P7GS7/2uKkWOnkh1+EIWlFL82faQBPR6cq5aJJdM2B2C
ttN5P6U5Y4hopsT85c6rtNLMYJmifJHJ0LCMFsY2AzvJjEACuID0yrwn/QCki9nQd/mpNp8/IduG
7G569Q2jpgSmLJ31VF9mQ4pBj3tj9vFtaw5GxmwD9i31uUzgvqsoBMvawbXiX9SbMntNUSQWpgxh
ShScsgNu43fa1kYqEiTr5yYpn3h2TRGFKScO10P/0hnQN8KCE94Ud7frCcsZFzBXVwpPMZ6W/TPg
ycCtUqq9wdo+BILnKV/LKi2jP/ayTvGgeBx9X720NksF4L+y6NU/HfxNkj9smE4StOqP6jp4etCC
yLMgfWzRmFebuUgURu1JIHjUc3/a7urwtjtoFupfeXkuO/bb+T7bDTNRZAPF5h8JC54esmUExDTV
SxEYg36yAaDRmZYHvvP/V7vhQ07tO/cOc74NkFT2hssD2xeP33O63mA69U1UzFusAEZbrIeVsZXD
Yddhl7ggSr4eJT98OvcWisQloelIP3IDN9w6QEI7tz2KMXCksc88GRJBblaopHaewxy//ZdD+1ww
S42ZciO4GUwnIEFSpEKA4UYkuLDWop/NOH4y8ku65R1o3c3aK4K+7yay7F0/+13iaN4OXERIju9l
TtPJo+wU2lVGhGk4WCgm14ZRrIqM18mC+pGkjxCxy/yshtzPXolB6aUI3QhmgO8voX2h7LssWxhA
Sr1VQ4PTPjmdMEBZnHGQqI7qTQ7CjuF4l/dl5nBsoegiTr1WlvYwVfvB+hiTsOnBcOg9MWomW19P
zAyqN1Cn2iQs8xXa1Z50TqT46e4ktI8Y4j5wCwhqZUguvREm6Bns1eE2Pqav7eZMDRWnXHqL/9YQ
EUPh41VFdrhkaRzVsXFplKH17AIQE18eI0pnA4jASL/u/HAnzZimn8DKbDV3/0z9/nWK3D2yBsq4
tsifcuoeIod6i5yXmoqabZxeS57/t7Udo36mQc7L4glq6evBPuhS8hltVK6yBb6W+8tEr9tQebaW
u3V61+j7pNTEhnTXeRLJ/Agdm+RKp+XRCTCtUMA2/tC0zI3tomD3acq7lGsGDoWPjwMCO2x4fAbR
YcUIZgyzWKMTb8Wh+TPTS8ghNFvPTAGNpj5T+sdn9NQ1z3Pu8l7l0UnjxJIEo1NQZRyjHxrZ+EN2
iPoRiyjVeWWfzD8aAm6VIb5qwUwJQorQmp0ktguQfHPs42ziLoXQGPXVyfSdU39rjRgU+rZ0q9CA
PCVVEQX0zfDmYIUL14bfGG9qFXe8R6zVpAoY5VA+eW3p9mQrx+VE/9T3VaIKE3glol39XR9GExL8
ixmdGksv7tWGfvekQZ1VP+vI5t7SoRblphtc1x23VHf/85OeH7K/DrTC60w2f4TV9vmAI+a1nMAU
+6DXJALMraT65b2iSjJrLU87sno5CAXu0hSyu9A4hjHHiGnY8x/mJucZxv+IpM5sg5EMi5vMBGW/
nqeMlnFHIOX1W9oIbmrZdsQDFENiwnh+jd1/VXfOwP4wc2EqHzQFA4F/xAO58umu/LfSHFn5ksjB
w4/tv+I4rN29bWdqE5ay9j8l+aBUlp7Gx/D8wdx+UajRy9mazD4mYsI00GJxQz5wnj7bSj75/Oka
X4OUesUFIaE0EhDu4ZrDSr1NyG1TjwT70HVPDpl8KeEMQ6ppGQtxXuzHwDjQ+iELtJyJ2ub2tY5i
sWjOkhpMbG+g+uoyc2ujHTtWnV//PzZ1LvmHSb/5HDFhjv7VNg7X5B/hUdANLhsPmdcDJzgKaBUF
D3IO6rCM0tpqdMyL6UsoExfheaJAdO4CuP8GRIjiSTYNq+/gSLlLN5d9sCjzNTQu9kQb26iESWaZ
7E3659TnaMz7RyNoka/AHQQIzGsNLx144Xg1+pYYHAaYEH9BAVrHtHEv/Of5LWUmU09LZo2FSW6P
jhITuNb0RdqXqaBS4GMVDqQX5eXFKj1TLdzJEGyPFVe9WmZgEpTfQtghgHHbcTpmjxx4n0OI9yWw
N2Lx5d+MSAqFm5nyuJiOGdGqpMA46RU/6dx4CFZAzuswit/owI5jtrsmEtvmKihYWyUdk/dZY/J8
WcKmMxV1qC0693yyaBb55FYLVce/5sftWa1omXtJF50gRDPLQcBn9o+3p44yYxE0YKNSi4zeaQX2
FnSJ0sX5vwBKf0W3VoDP/UU4Euuo5lCJ1OEQUltJaOG7md++i16MjJgBAQiegRxfjxzH6bX7nhSt
1tLZ6oUiqHtNi4zKN5RR4PteaDTjdgwNzMQG1vk3IePuqoJTJ7Zq3+5ktzXVVSKxFNXWBCtBvq1Z
l9s1Yblew/NYYMgCAN+RBZ7D9lbR041KU7f6B86+neze/Pk86JdBgqgEm8NMMKTHGVAaoBFfoGAz
nSrZ3kQoJgeF0914g4JVvkuBUgdoWTBgilJUdCoJsYxmpi9a6qQ9Jx67eCIPIsjqJB1Mp4Yn3ZPt
PR5ZqVCakLLte7Qk6VteJTe+QejIqi/XvhsSlhmMlyqvtWYTKwJm3WbNVsn+zZSUvr09bejxAuaC
VbhqRrqux4f028AQPcGIyjkipOH3e+77bJILtmuKUOvAyZ7z4GWmx6IZ0riyjPyqB8LRyiEk9xhq
FBFOLA7nIr3tZbAV0seB07jus4YBA6CFdpn4gIQPagL4Vh6GPQsiCkEtipcZb519uZ9gyOETbfX4
inHgqkVOunpFrhLKdd5mLsBRuC9dOqCNXq9YLPzZE6u2ncs57L8B0uCvfBnX1U2ITpIHgk0lBt6I
F52gYTtLUAh3UARGOrafSxe+Si+NFRrJzBCV1SZ6WqeZ/PqAN0JHgRhIzyLIjc3j+hHVEEUBS2OZ
tpPFJeU1B/2RzeP1hbzq25/LkPxr9m911rXv2xGjqal3nS/tyY4CkMO0V64DeMr2qF9K7BWXBX8f
wqTuCtoyyWQp0APHT099P8a5leLuCGi9FqKbE26ZH6v3F/GQxUdTvEWdM4hC4949A3i/oQDXbwo8
ZcWisjU/JTiRDefSqfW3dGbETYJ5Y52+wv2ZXv+BlbMAR3/8qSM8PzS1xTqBvijmRYg+Ps6Y9W2Q
Hi3t06nVGSyfGBIg6tFLwz9LwS7TWFry/80OmsDMkORfTLL53fF342HamGsLy39QpJo5p7xalohB
xF4HbOJHKXqfFko7Bphdzu+6TYd8p9yeoTAG3mKvZyqp7FsQ8n2ur5DVMy45fySalIiqw6Ag3oCG
rekAXU/pOLab+KT1dsuZ26238izg7f1oh7wXZEMz8rVZ+L7QIztT6KMpJordaVhAV3CVnRTJCxB6
i3SArqJWM+yhjTmnHuPnxCznf5B8XyTSqrYbaeNOqnUQrzEkylauxZbZAqburfbcuOtY3OunpJyp
S6SCjCSp1sCx7wdk7o+hwmiwjqn6/HogykR8CpTabM+ybFC1j0ovW65rLhpF/n8reS8JSszRsJLW
VU11wUc8xCDt+6il89aD2qvdJ0jFOjD+Pzmsin5Jz03QsZhBjJFPDef9q+OEZwteF4r2UtzgMIr/
R9jP4VZL9W60H2ykXkxEZjJ9ZGLAkC5zqsfVcUMYreuI0yCGC9chOrGB7xrWVTZ3CF96nCShYAqA
epKs3nk86D5BqogKVlgIORSeQ88orjD/GaJJk0JtacPZtDGXGPb5lAhr69SVCTv8WQwYP9mJ7s7I
VIE5FF83gabr0O9LYwiDMe1fjiLEMLO6KRN9Ydpk5QhpnKawojli2871YReSgO/tsnvj3e96KDrG
fZzWmhO+XAupPoX1JX1NUswOnGHK4WPoO6K7uiAH/uYbUFGBbOMVyeB9ZSChCCrZD/VZFoUYbiyR
ylIhRBfvxIji3ZHnXjZvH1oClFQypeIy/2ENyO2gB1OlzwZnpapimVa1bTjDFZkGLUxXxPqswKDG
uZHHWr3Gu21zdEw2fEtf5vVCEc+tuc6FVvOscZNClSHCBLQvW19k/NidpFuKxvlTJCw42Wu4m7u+
QSiBH5Usvxy/8xqLxDi8GGRsRyJyXox5nsbncnFnCQWngYlGSTXVeXJkWER9ZzqDQo5hA1E4uVjh
QwdlQrps+3e6Ue9cDWiH2UFyCEToNsst3QR65cLZSmP3wtb1TDt5KLYtxxsaIFIY6qtTTEOCHIlr
W6un3jF6bvbF8gwcm6iPDIr9JrUIAIcBlN1TjYURliK32BeH1NEKuOirEzeR2iYBZqmLve2cZ+c/
l+e+7xjv0r2Xuk8qDuAy6TnfYnoJo6B0ZAnn6rDGyIiF0DjcueWjuBQjtgVnh9Mgp6JMV4Q0b54+
b9tDfpr7lkgeE6yvjSaMuCjPiaSkuo/DDcRtvxTRRORdhzUTToCDNQYlAQV5lXmHzEsfELEe8a2A
Pencqfh9IGfWUUY/TmPthz08yfnGg89VpFuLlqazJPLsLQg/Ixwy5GgNctJGD9BlkmNQ9mqpEIya
Tf3cMXB49J3HHerOLicOICGlV8uqpMnCYsb7hnfRGhePjN9IaxGbgf5y3wgPujBNm0RUfw+bsXiJ
vxFG6AKd6FiYDueL/oxvFa9mbHXcVPMyJ8vCXEBQr2ARBPMmcwA6Ou2DE0XnIA/ACnqpEgnBJ5wv
/FMl8dSTLKHre2S4tKhriCshOlXNx2I9LAsTuFJq+QgWZx6hQiU4CVzlrJkuIS82CK+7jBnjGQXP
/1oC7HZGJlNhhWEN1bY9y917mNWkuL3nkkTH2P6fug/16XWjwk2aLVDTWg5uNzxU+31inDxgoSiN
qVEsbdscB7My1x3WMBUK2iChnSJe6CA1N6nM2RvqrPwppl2cpzMtO+H+8vdkEyxemktrl7ssJYcq
0OyjDoq1CZXVn7Q90T4U6BxfdjOpHDZFMYEeKnPCLWVEY7eJ2lVGZqwWKuo3zeJ0rfqI5XYxiUS0
7qKtpsFjx4wz6HVV7z/I0QK6f+i2Ms065z+Z5ElsP8D0fKERlOB5EVHA1zv0GUEKtvwRSi9hSutK
NHXPUtRlsj/gUcT78tepeCD1E9ro0JJDFMgqrDJ1OBFn24FrrSeNGIfGI3aST373IgMSzUqYvxqT
4UBYgXqpcBI5R673oIiYWDbYcjsnMlU6CRiedxlefhRkU9K6mh0txbZRZwszwUEvMO0YxiTzuPN0
RHgbVVVZaokLNGLqa4Kqgd52pJlLDW+Wjsjkxm3MeZtRu+TyUCyxQfzL0jAoRAcZUzHj+wcAGCwE
Sb0blpYGVDmHXvm646u4RvYoGatuxsKqyfLzcp+DkCpYA2qNfU+10Xyhr2HJcbpUK2hbs/31b/Nh
IAqrhOKNtWkrFLe0oOYqy6wyePRq6f7zL6HU4NlLSvN98UT3i40T7o85Y7gDZ7iMn3wSFwm0DSg8
WBRXydjkAfeOYkoYq3TnpjeCFxF4f5qUibne1kI7s1/UMrNI+bI0qOKDDrCqk/2yr5e4nhwut0Ca
0mwUpMq20nG/ghNWahQhSqdlY0fFfL30js6suq2jC5epU6WkrnQrPOLQJoW6CuGwk7N49NdxgUDr
83mcxxABtmjhdqqU3xSKRR7C/JivS6OzGTNMoFnarBFFuL75DowNFutpkI2MM87QxoS7qZF6azzA
Kdxz0UHSjiYt33gjIgglLC6sGw+e79E6gxIVl9E78i+F++yjESo7eKOUhQdh2XoWZ3bCiHZXNy/g
dd3T3gVTqP6LLMjwhY0v0YmdUMPVv/x5R59ZhPG/7v5vVv+dJSC+pqHrX90anKDxtwraNyAg4R8O
UW6uvwiX0w+69zF4m3d3wOwhzrZ7KU0sovbKz5vZYbtbrQTZr0UVUd4PSXPrv33ScPBG1ouct9Cw
x4w+pozVPYb9XoLA0rCAaONGesLKMp9GYtpHFCxCCP5E9rojxn4B6IpwpJ7v0wjL8Av1d0ScdscZ
aznAgOYlzlCDtPqYf5otSkfR++3jMb60njp7i8Fp3WMAf4kITadnZaXjNu7HLFCDpTTycpGGg3Wa
WkE91sQKBDCTBhqC7uYrX+Kst417RcUw6S9NqLoBJ6GZCqVbcXflhRz0aJIN5g1+pAlo1qy2jDbb
dTb8Ui+/Xb5Z7RQoPfrM4hfnLQ3l7HBzSjrFxa5BpOJ6dhwUFd8dEV9UzvTdhPXhP9cshPcwuZiN
NL7tAHy/o+dC6fkvRFqhaLsYMoaegb7BU9DLoma9CVUFCHmjOgb1tfjsa7FBhlTNxBh9nuVpExqd
vryGkgtAzyIkszFvL2Znd2UnSRF0KOtsGVGgxZIk9/53naIMTP4zA8I156FcwVjo4fCJBCSjWBEf
gBo1oXY/ZmaLMptRB+SCdNSYBEcxctKMX2pdxPf2PphWd8Jxf79GRoJ+yQV9qDiJO87+MnCB5mGc
94j+0Qsok3ulH3s2NW2UT4HNDhDo7oZVnpVFQAuSE/marWRnU7rtmD0wyw2RxSVXBs13dK4Oe7V2
57RpMVrAKlEelO1Pipi9auXBwOZ6P2EJ5m+nTCqGZ1vIdWZ4YR2dgLXyvJ/8YByBbx4kKqBhZkVm
URcQGKWkzOoui3ICctaCL2+KzYmDqGIxkgvXrEE6knQx52Zy5CyXwVESgXr1CAL+C8KqleMyZVMA
duuNkdVWEH4EKuHsmxDQiHGt5fcyMIddV6NYwnuiAqofBT5a90j3b5ad1eKtxFX8e+ehLd3QQq7i
UjJsiW9xTxwsEogc2SYNtNKga5AoR2B5+Hjfr6gocMkFR8/aOzSOtrosx9c5zAS1DGYwvit+vJi6
UH44g1xbmE9GibqlJY65kaifs4zmWDI426d7ZiTbMTCv/50QO1oZtqD/ll4I39Y/7xj+cyqBqm4v
DbtkZ1wiI4TnlZaLrNFGYH0G66wONBuWUV66ZNB7M/5Ff6Wcq46CCAgxYCDrNimYYHbPvK5oDZkj
qHe03VphWXPh/SlTloA8QyDx427S9ZQvhvy78RA2W6LHH/fpDKMNQ5QXo6762CBFJno6kXEmnf8a
Z7MRtzrrhYW2+U5qcCdEe0aFMPBcvnPXcVcseoalKaQirYVXz9r5QXIQRBiGVj3NhYdWzA7sjtUj
3wObpJOhUEC3EeqRwzHHRriYVX516yNcLSzBROhGlSjS1FuCvdenEDZqJoUn9Q4PJmuNKMjV7VzK
2g74JovssqeNe6y8wzSpjKnrzS3pnkK0Q7BGcVFoLFq/q4V+tXmUisGBc0x5L7it1bauf9aKBelq
BoQEm2Sxkchup+M8Dcj9/rcay5Et1Oy9jwnkdghsh/B068h3aan8Led62BcLHgnRPAbUhNggqpeO
xUXkerIYVHu8ZT5hOY+0FxhpQjYT/OuJnsOgY0s/eIDwkTkgYV+N89xri1WYbzFi5G0po6hcWKat
KJ8WojaR67IhBbFlr85kybBwM1+L8iMdGi9FKRuMLIbg7E5kv42Tn/ys1jNxnxvXy8X8BTmJsYuZ
lKv99RTUvlIYGqqOtV6qdp90Up9EPc+8o3XDtGcYRmsCIpJQw+3y0Vf1CdVSHZzu3viu4RtLWiDD
J/HLNF3JNzxthtCC3v4xG/0ZsgcYP+cLkKpAhzKq8wiHKCXtF5TS6bxHkzvd/SkxDo+VN7nZ2XzQ
6TI1Mog/XuIMhJDrb4SbIvrVLWqcGYyyMufTs4xgR2TFwVvbjD4lO3zgws/OL5lPkkIayBtTE9np
1lHCw4DjQ/PXpjWzkQemisZD0phvBm3epUNVE2ZjanWBGSS/jL8EQEn3Ob8yR/H/g7L1oUe7qPH8
jCdRWqwqzF8pkd6zDL37LLM9g31vhr0sYoRdFm4ZpPGmFokrF84jZPHkHWSOPXyfQvZRqlYjtg4L
pwmw4Iw1d7iVc7PG1Wn8WO4DYOhSeLQJ1uRINlOW8S8q6NpEdimmtwnsLwetPOg6K8GqDOn2wzPt
CAmMBwMyyjEV8ZlRgESk0Ps/vMDxKausc7fGanTTpeOKixnKK19aV+arVKuIgeKO+tKxiJqjqhqF
AQkB9GyKWyD0wq2hZo0TJQARqYUiXqecgqtqMqWqc/bYlUdaoywmk3D0WkW1WchYzJXeH+gy9r/K
P/hyj0FA40p2zCqOfr1Q/5n7hSkQUe2QzffnyXScd+cnb7daCmuXlFqskUwKRZvctxYVcLcDhDS2
NpRrsCUjIto+mT7JGk56tAlnqicNTsW/DHcvqHJf4Uv09nbL4Cq8JjufwL/ggw3wTEE2fGT4cdeL
hoBoVFK3LMtwV20bP7MfIUQUHemWuGceFncYZPoGoJhVjbmjEGmVr3xgS6f0GFrg1O9KitPTjDMc
bZ6ZXc89j7VVZjYcwvVy6/roMWKsCwMYDR7kwAZZnNBLjvRQblPq2pnx+cct8Jj6BiprdWcgfQt+
vmckK5qhaV7yAyJjLnVGRme55qvuRe1nHYOhBGDFJovva+nkE17ypnEpLlC9thVEdsWOazDRbvfg
w+3KUA/NCemL/vHJ+Lr2PsfU5+sOTBwmC5/trtMbv5wFyOW2MJ3YNdylkJO5pfQszFGhmAnHr1lh
p2QEWtAzvkRWKUDaai/qjNxqqBK6cn1nUkxhsfquxekf1LJPLsBLA6UCWqPxXgWrTeV1ZalRek/h
F+dB9Bql2rvva7kzCuPyCZUsCebkPyPIoMQxUneoR3Nn9A8tekBfVcZ5EGJGQWvQFa95yqMgxL/g
aDETuDjc0BamxKIahn8PvmImaiURTnq624UJabMsugUDoPTpLRpkTZ8Qb+yoNXG95wFlZv15Tkka
cbuSXPTExhB3bLW+3j09GT0y4aQcmdF4wEDz1Z1TxSbZzDcUHj51zrXl10cw60UwDJskT3QIHoLn
G7EUBQdHTUBKe4SU2EnZZ99K3poO+0CJyfscpMRIH47t4xQxt2ZYtvMVacGVkvD8Pz4uhtlFg9ge
+p2YhEMib9xUgCThyV4Z/4htKlx5xCWo1t8A4Rka6m/E8SXMVKmOb9DeqkQ0EFm9L6jJ4Y19l7JY
j/r1Dj7XvvGhytF06H2THj21aicYAfcf7wPBl3TwV/aEqgck2JF/a2I6yZ3501Iwzmh27dZSZTog
hbvgjDCHY0d5KOQJS2CSJemoUdo74eZCCdO1oaeCEJmCPbtpz8g422Wwh0TOC6DCvGRwqmXJ6v4L
e7Yfa4+hCkNc3MvUCJAtpPM0FtVxDkVJXKAikJU23ztO9XSJnYadOVrN+a1uULmKHmycXuqtAS1m
5ksn+oMBdFo2Cxy429TRt5/rUH9Pc4uvD9B1Q2XjW5rmqsE7odNLfUVhB0Jqpaq3UPWyDUdRg30h
wNjjBBqSpuBpP83T5uDm2GETNEMdZSPXnCFSHpaOmL3inuMExuSm4e1ZeQT4ajdsY92cXZIsFuln
GX7x65SK7O6ZTM6oXgvNshN/VRjY1pfOovGOGApVXduHGr5kEJMTPPV5/dS8aFOVXOUFchxa2ARX
u4tD6uXBRQFQ39XwCVRDUj0d5ZYx16/obbEDIzK9HhA+NVy/Bm8tRw44CvUkXpN46m/9X+1MNpjA
hVXdpAu1kiBAtD/gRMb463FlP7Zq3XQZEyGks9YP9JIxhINB/iRQXNmT37YTdAGP5KNWaov8wm0e
DdCONQk/XDVnfbXz7zM6DJDrhsPA7M1oC4SjlghMs3h3Ad+n8/k9BAfyKHFdihB9coJdAOSJDV8p
IijqlOJ7OxtDf3CmODdZCfnXfxb1T6lHbZSoJWIK/uogB3gGU2svOzsY7tDxer/D0R0OA6fAQwxj
FAJLBdJbs7pwbgg5cYdD34h9F1aDuZD19FhXI2maw3db0Gg2aXdQh78GLKdEss/E5WIn6lQhoZS/
a9pDM3W8f9FYxS76JWFF+SXAJ2vMdYWXFPAhMPtPS9CITElEyUtyR9/1d1S6ewcXA+qoQKwXMVKL
ZtNTRUAcCvfHZ5V0joq5uCBUySOup3mMFOFFGoGo4LotfAi2zPxKZ2ZL2nMELOsVZWtUmTXKIXp5
A/qauNQC3y/M2lqcktyNCGthQOKi08YAJ5ZEh9ssKWAP0HiQcZyTZe6OBg/CDu9agtBCjSwReIaF
Z5FBa6VnU43a81qAGXYGk2LtU27C2Ct9/Vr2O/ddW4lOfY+e2ZtlEmdxEMzVNKbygYYgNrUQ6t18
T+CS1EfidsYbG2RCSkRPZDHwr97xH4kNf0Xm/+zOhMJPGouNteLPIYGnyK0dfdXHFRZk/f6D619X
dltgpsTxSZ56xMlNdNc5ti3SxweM9bXroJQWQfhTQbgwxXlNVAbxqG2Y0qQucfbS1ypwkkuyRAFx
0LbfeyqHKNDT3KVL6DRzcymOb/JnJVA62Kke5dw48USMqMj+nZAOpE7n1z1HSNpLTWAEneqwr5Uh
C405qp+IgOlyg/0CBfYpeoD7Vmfbh9bEulB8ItWSL1qi4fbwJNc9mTJNY4iDOdnpexzJ4ZS5hGXy
j2QVd11Z4SZQj7bq+Lzhn/4J3DDQYTx3qD+TPwVqFUEcZ4cWLvKikKsl9VDouWTcCMACIMKfoDfb
lIZSSqDow5HRBkuyVs2NUaG23PIClscLNb4ImGhnNLz6fcx/ZJaEVnrw/OoTWdo3/a0CGpjg1X1Q
QUBiYZ6NelXZZ+pdXYiqkN2Oz6xa124KDlJkhwhAzCCdZB9IL0GbeaKNx5OJ08FBpZjXkpYwRxAH
b9MqJQEvWVLkBsuJj05XG+6iXGJ6SAKEQi4v2TnFpNoP0t7I1MS4r7r67lDetJi7csAG2v5PHuJZ
fYmYx5gahOl+oYHYFQwPUj8+vvQLTA27F5XTdCN2rwTsLaCymm7NYLZ7dUyU6XTkxA/eNQPLgt/T
3IET+tst5qRMNj0lP9ixlqDjiIPYhR1GyNBRugG9twxazWg+KIEabKWHdyaQARCBdXVk4BwvqX+f
MyvCkybemNpgI5wqybTB8VKQakE3GKbWWq0bmuCPBOuwf/fLvLhuiQKWVDUKDsxjewjAkFq0ImgF
AjrPaiUdcjpsbquRwSAzyLQrcraCKq8z7PWI8xy/mXvM9ADuFfx2PtDaHnRlecyu2oVG4cB+mGGg
W0S/hl69tHUYK7cwOByjAK+FmDu3nqFn8Rvia2NGe6YE4r6Czu/mMaqM2bcBFquUa2jDgNzMxpUN
yqXcwqPwYcBknAzHbAKmaqs0FDEme5AuNyJ9Pe1pLGEcdiDX2c+eozvb7+EMVzK3ysYrCbx22ETX
U7MmTicMLKO4zLrtpwZ2WnUnwnNTJIBStVquVt/QZv5K6fI12LgldOzaLJZ9E6/GtmyOHkQCWTSn
33jeW05eZUHXOpKJWzt5oJ8y3BpvPkUi9NeuM3yKvMpoDbOKD9knbNtpARPx+9vr2RT491aCB6RG
o13q6p4gGnzXDnJ0WNTaFFJRhFxou7m3iduqTu/1F0A69KR8xvE33XWha3aXcN3YMvwF3CyLemIe
at1UgZgJb5nqy4O45YRjRyfMdAx/oDOcb3fPwVu6xgaRcSeDJ8lx7jyb6RdANOMq50w3ALNgxfuV
czqVe2TdiYCE9NirKH5FnimicHaQryDtpuEvp4917GtOeOIsvgnxReaOsvtp3RB8h3fSEqtoyCKu
yhzi1A9xefeP+4kGA3RqQfT32ZH4KyozzVFXvVA2bOxeuTs8ZRHJWpT/4Kxb6sa6H5JPnsk8yE5p
+Ks7By12U1phjDa3PlE84/XANm+Ri5Llx/dRMgkQLgRaTDXs4B1rvQyULbM9MZf8NnCUzgzGzRNG
p1EQTSId7bOLcZMosNOwCGLQ9O/LArDZNcGCDQswNAw87xdLUiLwPZXchE+Fo+q0KqfPukNMsWML
v+NpZVYFCFX3cy6/MQ8ivkPE14wPSuKtPX5lIgCfh/SyDA9qn8XBLh/0Sn2TNtlKB5iSQz54DOJ5
ZhaqiSk3ILciHBO8Z54kx2DdHyQtd0YSX9Xd73IhZ4iuK3gh03te8d9Z6U4kP4epNMEOUVZcwMVr
WaJ+oU6iW5GIz+XuXU6+WwZjmTZBBZtJVcYM829GkwKhv+yxW+rWMxgL8H51k9RcEZpU/MLc32l8
w4mLcw8XlcP0nNDIa5458PL+APHOsdw/h1N/HSG+fZy5iRxkGaOpR8tmyeiEct5GDaH5aMGy23rk
sy/Epra9nPfB9iJ3Ae5ztOVGgQ2fI7yrIkTVPX3HHyrtywzNN3IDzfHISBhjp+6crguJrpQRUlHd
0RW+PjmKAb3xrvq9c/3QZPfxvzt4+cYFThnsO13kVGtuFEyG3GNRwgTHWHz4bdCjB60iXOfu6m0b
KyAG3fudkHQDOvTUkK5e755duBh1wid0Vmx7Jq+J89VRayNziU8z2LYk5gwmQmEXV4h0OB2tu4uV
l9xsmUtHRqh4Uzh5UeGjYIV/Ut+bMrJLqbbYP5OkZyZ4Nw/elea5YWgaRQz99kWTqUt6+h7IdFRa
fQ5ZKl4WQmXoXzjktg2johBhG8HnsiIVTzoZ32W/EBVzBvAsMNUj/88en+wp73Dkp6usF6Fup1Yd
dN14hXFNvMPxZqEIpuKF2ctC5T6RoDKPZ9Eh64AbDX1oBKuXbH3K1NlwaMJEZdniZlix6V/h8VSy
+WBr8/238xhFwWxUrPVRPTRXO0eISbnwy4bwbDSp/g+TXaMi3oSsRJ+/BmC0Ijwa4qvQI9AzUfrT
6N5XcoIfIhn0Khwd4Bhywi8BHGVB6WyYV5FZUgY3fHrYNsNE5XtlGdiV54VMoD8utYRCMIy00AOb
ebpmRkYw5wJY1qCjV0llk9P/Ts4Vs4eSXF1CVZGhYxgLi+q0g71SglhnZTetLITOWOgnXtxlw7sm
Lb44YTPAd4N+x28gqe8PHiECGNggH5O/NQWa8HtXiZ0Sp8oLNN0z/tIyFhXeYmHyXuIiPXZl8zKr
ZqWE9tbgXqCQCQNbvejOBw6oqW7MIB+IB4kUQ5Mx3cRhpMbbbdHJF18ETHfdNGMbemuhdKz0b6+P
//evJ/4ctJO/UHJKmB8ew8WgR64HG67+cUrGhZYw8PilGYiUlMd7XSQUipw+ZmfVm5Wlx8qWf9tT
2/ejKL4WxXdpOC908o88A/VjsGRUeyoVi1B24ixJgVppkCZtTTmbiRNhDAboOPLlPze5x1+jZG/Q
Vt9u64uHsIaJISGW/U5JWOYOEskbTcJCKK7cA8v74iKEL+pZO87hcRZHsSsCjEDtAtUTkU63vVwY
+hDbXFZgtqO/T0LjU6j4REmO8paKxPFr34un9JHBr4Mrxaj6XGIJqA/c7vXz5xuyxVbC14RUgN9T
sA6VJtW2MpdJnVBP/HFu8Uktmc8J4fVCtCP/CmRH85ud1jfvmequLvoyn9nUWsw+GCdW7UAGI3gA
FevItO0X2n8YK1IN/BtRHs7UfFku13dTueiX9zLpI9sSWsDcNgiOj/iWhPw8WfqOEKnv3RMfo5ny
iCmgWI32Y5zs3rJvWmN9lqQjHN7UsOnVHR1XUjwSI4fwOd76glh0XV6YekoIVPZgFXUM/1TZ9czb
3f2VAzziFdJRFoWAnlcefVjK2NF6RSLhnXqa6M4WujBZj19IRlwoFK7ks8rUvwa4FqdsT7kCpr+Z
xbqMpCDyJFHp0AAKnNOdp+dD2UUU8jkyBBs2PTzdKv0f1x/M7L8INFDyvbdHVKFZnTlDu0kje9Yn
6FMoheqDtIf0XlNuh3vhAg6rcKgcNryd894ntQQPGcaj5ww1iPOcc4238RqCLVazCIbNSlwUTUhK
W2KvteHuNPJ1stypZxwXGAcvD2TZ6915mqXtgon4b8hjkTOoy1H9guBwbTiD3lGTzOENdHGr5cl9
xEJNoYw0naV1tTr+NYD3jQa2ouSaRXeDZSN2CmftoUQWyMvgFzGRu88lThkDzkBtG/j25GJ4lCbV
1J+kBYJZ3/NAhzO0D71IQIJM/b9wmedHjUnt1Old9HPqRYgie6UpdITXL6UiSaZk5yCMWFDHDjWG
jhOc3YhogA0TV4NW0xRMKZG50lZ8EEpEwJgjtlSMul2/GwKHgUzX7/c6L4HeKNnrn0ueVcSmsyPs
7Um43+6XnGtq03jBUYRFkP9pDR4m6ptP2v08T0o8jxMk++E5VFsOJgZcd4m9JtlAO7zwiEss+Lcj
9zyn3YLl5IRlN6hYZrZwl2jHRLsz0+EkeCuGPukm32pqR52k0BtCJMX3yHFpWmc4NQTuPZwpChFY
FOQM3DIRgIs2P16bgIwzSo6s8tSCSYWi9J+4wSQMbwrfKkiseg8lBpbH/xklPbCXChQVPT2MkLqV
lw4H3Rr5/0SJNvXFYE++U9BFZU47rfMRWxYxFHpTOpM55nkxXo8DrgTVM+e+B5p/CR+yiVefauOy
Hse0hyyABuKX5QXA5+CkTwCCaFAfUqszXcWm44JyQQjItfo7/qzoglL/Rm769p9fSEATcieVmdjU
ZFl4NiUaaLiW718ZrIZkd52Hwa3zE++B1iSiqTxVwlSUC/pSqe4gQSY9rQzZmGfoftDNNlEvjJhi
8AhlCz4iOqZvL0t4WXET/pJNVlXz25joDrqrsrxj39HKSgf6rLXgCtXhV2avrcVxvCV5bBP1FTex
H4aEP/XE/1m+3iEY5NX9vtZ7fpBR7WoBGltENobd6LW2kB531+cVIz9XP9GwVDbaWzkgGoIsazRX
VhnJuptOw+LqLeVGWYcvSIA0BgM7fs8YseU0Xboijms4QtmAcb1SnWSQiffQ/5qsOOokkEBbHOWU
Wbcoi9VYF9dWmxI42TYaxvNDu5tSOSYOfwg4OazneBIgjFYhJNQOT4T4lvvbcPiWn3+8B0FJoj6b
sIRu/KOC1grVqko1dOPCw/IUMLlVJTXvZR2nsrSHzqVqlT7irjbh4kT/J3icjsTbY/i+S0/3sVff
li5MDktxzsP6d1t8jdwPg/8yQ6jwN538FYAzUwa4qIGPqGtKf3i/jyA6Twn4+vAfUO9isWg/cdTM
hoN/WXrWwCQxuUwLU82/Yc3xU38Xcsd36uSe2/210fFJiC9wAmsGn92lYEoqXNtNkKqHDBf6r/lJ
aEIv3TcNG0zN8x8Z+h4Baq2CKRv1tPLrPZmv21as0aABwDAUxavhoKgk2pceWzC0Wif7fXqGRSie
MILW1jgRnP9+dUAnYngJGW05XN0qyB8LHvez1e/WpX9JG44EmTpwMk2dJBra9jYooUHLoBzLcYo4
oQAIHpgK4hUUdnwjrlYvGnMqoewmoiPFE1krZXD7Rw0gPUULjlrgwZtp2A5Czwl4NtiRmm6KmrzM
f/Hokr+Y+5XNiwyYvyNMwtlSzh7h/07JT98t/Fu4vqV5hZaTAQL7hqzU/iYH//hn31hvyo+vppeM
zXuJPh1KO/ZblcguIYuJJfmzOGnEUvGrtf22tCV3IPBUScHgXjmMBOgif6UkYOir1vhQ3OJG3gFm
awG+WoIdVeBpwHbd5EIOY4zgCgzFkd9/55yq7PAHg/jLF9d6fT+mpjpiwon9VpIoyz6gonfjo/4e
B2QvFjicKnm2jRMok/iZ+4FSZlKoFYB6BGCWsfvHhKAm48iS75lpFOdFtRbZNMvgAL27fRfrNKTS
/XpwLtwUtuYowUwQfuuyR0nBfU4wHvpLwAL4scYJ06e98nUM/EecEMluUeGJoNzVCv+UhEd/hD0y
32oX2lNBhS3QMMPjXziVUUcaQYgoncQNmgnRMl612IFXS0CrJZG5xQfXqjIaNJnUTrXb5XYBoyMb
0nu0wuUl9V51hMzrEGZ1FWTsIfSwPFdT3sIm76mUnzSYMogwrwcdzBm8+D0z754TaKEf7Ymb4HU3
WuE16dd0mlY3MM5huihQxGGjS9tu1E0MTr6sw51WpJgmX7TzLNSuXaOdIPgBHjKNPy87B6XJKjuy
SXaxBCWQYToZYV+8OzBm6HGK6Ficdeze3oMcISmNy7RWw6sUqKpWlJviKP2C+z07Wvftzkhnfg1P
4OxOZAtPP1LIZAbHrgCzJRx9ICueWY2SiHJqnlsgGV/KbkHYAVjqlFSw30VEKruLXQklM7qRDuVz
1iJX8gd64wcmapXm/BLz+gO7hfyvh5LxRfEvwY39XssZwXzFJyQLE7f4/LVbGKh+lX49gNr1rzfN
PplfUMe5ELoC5HDiMry6i5X2Flb1B6fKGIBzUMeU7+HXJcrKQb6TDG2eOBJN1ZZKfVkuhm+VX6YN
5i7pudB+kS9O9x2I3LQ6cAbs1jTbfz2QHjJRqsPbDbwK6ZxHHTf3VTrUypKSLAtWtJ0wfggOz/pj
v3p37Ey9mPm3Y5Cf1T9zeHCM9xyNaOihJnWKp7IPU5a4TTN6EolA2ooXW0poyQ3lkgMXiQIj1BJW
Ps9K8Y1HkIVJ2wEoot/Cv4AABFBf3HmVBvW9vBHqsrObG4mFWKxxCBIOQYa+qZE+ITYNVHISL96r
oOqm1R4a8qpD9j1gLK8SvsCTL5+jh9TWpiVpoMaveeM39cTO1vNT6Lmb6dV2gxIuEre2VoHQqQuw
HqiMhdLmZxgJFrAdtLqa7qu9Xtqe/ZKikYhiRnN+w69IZDLMbGcYmXM9JrHUZeURF7gCOqbxMXwC
yFkHT8a6rTzz9eOLF+Ga66zrJGYo4NN9iZBU29VGL7POLqKw1ELdS6Ndq2knOxPo2AbvkrAIUCOs
Sj3dOZxKpvhfQVXoWS+qBALkkZhCiyqX0q5Dm68KVbxobp3O/zmALgjS8DFvnvGfnohFiEeLKP8e
S3YIRcCuNXjDYq4VLqQbmrGoCdVnxr9krGhNYp6I2N2/9RlXZvyg/SdPY79z8BbxfbbmXPDcW3C9
TXa1LWzP43tEF5qyBNEBBAGRQmhFL5lcwuNHh7kMHFttgpU1EwWRVj/Ayxdy1Z5/l7F1YWbD8+/W
h2rECgYC8TNR9YBSNGRyWADwof6lA5c2SUSxsR9qtx+QUGFVXtw0iUVsMpOMSm8Uv1N+2Dg/Sov+
CgBw/CqMFmkhVAvoDdLFBi/lKWCQjKEOQrYC4LxGppjQq6UMCEXBzub74s7TaMcZ3OalDGtcDjTR
cxzoZK86amKJm8LExExOfviwvhoTm8DqJiUrsjbs1AgLkuUn5uSfgGI5leNRf0aYVr8so5JQ+/EE
qZRSye5x7QNjNvz06uIRSaHCwg2YNLI7a2nDV7tUBOYHTztkAklAX1Jk8uI1ue4H4IHzWbRp95fX
nuFBG3FviWELoDWUQktPgK5hJzrfkFfKBgTJuzs1QAerHEeG9tYpcQc+KHa/M2io4IpKwZLvaDah
tCJegJmjgiq9AkRSLEDKf6spDb2sUo5TaqIOE/cw8nmUKQupjPgDxa1pbiBT4BEZbP4vb8TYvx2p
SHXLq/XsVVx/KiUqwQqmz0Iy7HJlCDMNa7VBQm0heZmHlDIiMI7eBnmS2g+hEPway3SobYTKNnO1
qcJLrLcof7UM700hEjrJj0Vm+bu/ks6gETJuMNWWNTc/kjMWIit4CkQqD0obJJWlBRGPeoiU4f5x
ap2Z0/Gxy2NgOq9M4/vHbWrteB4ej7XGOwNIHDEJnVxT7HJeMLxnMd007ltzjjZsD1znAVbiefXZ
+rk/g0hD5d6s79y40oJoMJ6zhqVKQTgAuQ7p3R8RRfe+1r/+7M2aUGYZP1twuXBw7ZwbU5ndAcLJ
BFS+e8sy6i41gI31o2VSl2UADRlWjypiUYF4GwFjKFyVWTdrlfggw7gKvE9CWH2LGUjCUFH9U2qV
RjGdnTs7m4vyD/gw2OlhZC6pzO+B8KWOjUWs+Xbm54g26J5MEDGNpGuwGZEpggMxrhNR9qzWL4rT
14SJXqftXU/J7ySL2AC8l66Gsf1Er/+BGhZ9uW8Ja6quXYaEoIMOf/Cmjkq9gNcHVjaZo7pPofid
AtNbCUMsHWovJtiTKW3o4fa/KKwT593iodrydNDWL2b9aTqfkXJKxUJLCKMkFSWJUfz3Sg5ZKx9K
lwYot8riKrdDhusKYhNBZ8deWK+Z93TArijaz5KAfxx9haikgMeXdvWSIvbWLdbHoND0LIHQbwsZ
WCzsBeQ9Ka+F/6my9m4CfXQDFrcq8vEEsond3tPjnrI6ZoMB9sjm8hqN7yO6FXlFXey6DMayHwC9
p0hDw70T4Y1Rc6HDn3ecmCMniJpj81f6Xs6Pxy1yZDewUylZXCmujzXx/YaY/3lfHQu+ys4Tf3Pf
1F8SHD6BFBt/jSMwoYfeODDBl6sn100SMf7CeBW82EbeoVifEWhNvByc075A0twpipc8nD+HQmMj
jRy8d5nir6yXRY4Gakd294Rx4TqxsplUcAXeeDu41ZGruvwN3ZkpnnDoAij7pHWgzsp/YVZyMIXS
c7/mplO+j1CEz8LXE1T//vlZaFhASwSPZ+0LSTWROH5a0jidAAETzE8vJoS6tW7+7qj7SAerUbv9
eHP3hixSkH7qFvYezNmhoMXSjvT2pLyJRuU/rAKJmd8b+qRUlklKl87QH5DnQD436hyYF/f0Exna
jgE/zXxE0xG0RvyKj4NI53/gkTKG4qBPJ0qaAXG8WR1DWWl6AVJcc1I8vbi1DEejSDpr9sUm6qvm
u4UHswHoqKUj4mb3Y7RyLKSFvg78nItI/FnvlDThhHg/vxvC049Fn2LlKyfDVlm+7SmtkZbox/HF
qWHnAVJns3cVCHNcNKm5dUaVOdIvAWEi2uyoD/l1/wqwSVFA483i+NXVjxEs6ogLXaf/45OsCcZA
sCXervLBdFTNERvboPjao0e4t489EQ3LHDql0YaofqNTibwbwkEOM5uJPZJ42xhdmfue44hybgxX
7XGdA16VOfyzV25N2nZNxwvp3KB+pmtuS2Av6ZzQIsXtu9QDg1Gu3xik0+UE/2pigz6HPMYl/JbQ
FNvdwjPd0cPg+Y5C3aFr4LurhI1Nx/B0jcBNy12iomDsicb/Y27AcV2uagezByNDvB5VuQgIQ2tE
laSBSEqQqLrOrIp7/jBSo6dsyhPKPGJERJ/J7ADmnDYMX/nx6FRpJ/XW0vhZObYje7P0yvWwEeF8
Mlmx0XIMvePIn7xRs8qDIz95GLTksJkmMRP6esbPlDjPjSmeqXlglUMb4nzS4CYvxElmuzp8R1fX
Wxi6o1v9Ji+aDABcXhHfBgr2cMGLNXEOvxx0GTzdtDHINBUV1POWDWi69CQz1qXy8nlgChKh9fK8
k7JEl1P41pToWecorxGXQe3tubWzm0Bvdg5SQr5SuuZPb2gnxqKQvlO+6rZELPUq50DJUaiQKERk
z+ME21SJS0BTWOcddBep0SLNdcEXct+Vx3uMyoeBainLXOXV/1dqZ3JvmbiTUMvh9BC56EZeye1u
ZefNq/1wRqrmKz3nV9INaRcUwjru7HS40MESlLu45/Tu6SqwUvNT37/q394cvuhPgJDgf3gkj4Ur
bgX/wvOTB7UKBO7HRsfFJTYRrF9o/jeuv7YQ102quH9/+58/apb94PMbelNy8dcwDR0/UQsB5y4A
Xo9/q0Ml8QXaur2Oa9ADfW7LwBe4rKW3/EXQu7Y/UWl1x3JWAfAfP5SHi/R1qGzWTTW5cOw/X7HF
cFqO2kyRgomncVvAVSoZ+KIP9GwBU6h3nGNjJ9pF246EJ7zlwXBe2ywagPaGkEjd//qEVCL0cqaQ
Vj3a8cYFmXKmdwn8nWQCiEfdXa/uU5hd9FZNj2owXi2+ISesg1TNJRsN1IVyvQqh/06xCBphBAzY
wY3LKhNLAnCc3YrThwu5rNrXqjtojVAUmCynBXce4rmz0ZSLiNzT3/PPxbmkHoX5BFAjGGMHKCxS
BKRCqF3WSTFxhLMRZxbruQ2iyBHLGrcYEfMEFbTiLBft/XaWK29wWUxm1lFgSJgOQyNkEMfzprT3
nvazlcIBwCgmX4b+W6exYl2OsiZmtQalIu7TMJU3t4ZhsoSFxkpnB8Iq9ugh+cAV1c66FOtAhbmr
aCyO/xrZPHJ9TxwaxLn+Api2ffIePBb5mhsFNFeUlj/uSei9Jb5TN50QTZ6fsSB5MbynLnqFPpX1
7qavjTDbOM9tuIDszXBtS5376WgblX/Plp+pTNYBz1pRIZjvYDI1lgm1PVGipE04/SN9eTbHp42c
SeEkoN8ij32qBsn+XoC47BZJg0pKH4m7I4L9KtXBg6rWQ7UYRD7EkTXfqTyn2jV7NmN94N07kbGc
Xbd2RhYFhjNwQ44cXNNsXpoukw65se+rzWrk6IBlsq+kTh+KaNegUl3vM23gljRy+R5cNSTbdYQO
Y4e8eJhTvy54r9EM1CA7OrDf8WhKsnmBO/3fbGiKy2sQrLGAs6aLei+MoKhhlxMp6eVex09OXiJf
EWVbv/KjByKLuhIOHEEHGzRkEgk9lNGUmAoyM9V6PpxwPayZYm1QY8GB/+zgfklMtBp33ScPWmLP
YkpRgsMkWUHaqeiCRPVPs3CTW6PLZCnqQ9dAC0x2m7aQpDq2fE1ixR079Dcem6oraLvhzfFbZHWe
x7YZhglKT6QvPy7VI6Kp3mRuCyTrgjwVygyKOVM1w4G0vvv3IXyo3rQicnnKjzunVyyyaCbcH9PQ
kZHfQbPHV3aDAXm06pTErbxYoGUgAECW4cAa7zu97gPT54BlqG4+JfHfxnOBZwT2GbK+fKQpu/xK
rq3incoOeOu2KMf4IX3lAg1HzfRNiqwhTXqLccHd8UoA6d9sewzohuDd7FrxasIE++i/lz9VQt4J
YC4rsj4fHfWAkEdOzAjUPhIZaOkjCoqUxeSs0AoN1JtAvpZ7ldWCDvQmX+dT8amZAgVrTknVEjqZ
CEOFvE8WH3Majq4vVuOwIpIKESFQFoORZ2u8nl9T68NoY+vMASBl9hojxi2EYw/GFLJ1DwiAFwwJ
o75p92Omj+5oeCl0k06Ah4pqKlCB5VgbCJde14iPq53rBHQ/mZWGHJdxBZJ89SUfkpVQVyoThw9l
dl5ZX+4mV36elgpESDFBVmZIRqA2GyJRatVI76Nap7uZGWV3J9tSqt6Ktcyj4XdYf9I5KX8Myltt
Y/+4i0ixTPR0ot9c9l1iIN+zdEXot4yeLzZWPdk4JTBacMmH2jQOyGu3Ce2x8AL1okIhSlSq8BUl
r8wlHlXJDgT5fACmVMxykTHxfB93tsAqHcqbYAorVI20Hhgm38aGaI5bS4MazapfWJh09IcJtMjV
4L6qPOMnJqcr/Y8euMH5IufKMKfukZrv4vynCy1xMwvYDWiIYTlMd4RobPayCexraaJo7gqVrMA6
OuYKi8tw2xq5PgK9fGCuMumecZVmuisa/1tq2mmm4kZX9RgTL9NLsRhJv9IE4wdoj2bZJZm3gaVh
hu0Y+Xa4vmkgA7vdOdyp2j3ovCkhf4jD8qsxrNQq55Ksm4y4JVFIgzCv5a8CfQ0qbVxf+BsJLyC7
VVXg3bRprO0pbk+U4DX41+0Zs7G+GWepe+EanGTTneKQCGkGlHwiLe4ayLITFp248q/O+hjVAsp8
w81GL6gFIj5qCqJv/mju3t72Dlheir5s0OhIWjcuHYosQRaRnRz/ABb0I9WVJL2tRtk1/BbSjePK
v+44PDdul2khvEx4zjIhplSKPEH87TOwc/+zsrwmkmto9pI6PUjMvly7qYZBTjTlIAf9uYE5bC7H
JhBt8/R1bughgTcJ/XEqYbOki5zTzxRWd6KYNrYxzuV5A7SGlCkmM9FzTu9c/jei1oLPmUkvzmpK
hg/obQu8AFqfOxd2SCblrp1cSSqes5DwymUa2VhyuL1YWD5kXliIgOSYzenDelcQZMxG+65BhybG
8gHDJ+6pQwmvi0J7qRbdGsGZybwJJOhAArRYCwzZpmUSoxnB0gHp3a5EqYWviOebCVGGnSNjUUkA
TTmLeyU+i9R9xJOCs9Z3+60DgGjg2t5nthnRmsUZdkEuldN6F4zVGS3jPMQMkjarMq+h6gAaqUF8
euWT0USuHZ0IQz5+HiOk6lPa8fCX0EwYyiGkSL3RdJShbCO5WD8iO9Z4SvLps+M3uksJhH+NUDYS
nhhTk1ioTovbi5BL+wvecl6eIGWrAf+SgNO9Fw5rTAi8rR4UDjhjYATp6/NvMX8OUCDYI6sgTSU5
vqesrA+lSvoXNfy+C0mt0SbLLyBemkA5opG+uPxg8HCFR6N+a+7GgMevxlycyd2A3AMGWMV1frOR
CdACV8HwJ3zsMZQ6fl1tYUogtnbawT3bjde04mkrNveW1zOrxDm3hmq6W9NVj7eIv6XZ8nvmKXUP
/YfrUa4Ex+7aL5P86L101Qh6LVuaY0EdtjsXVz5vMtkUlNlSFlAnKHDwu0izhHh0S/5e+9R30SEU
hlm6jhYuMqHKHxytErrFcJ7dvDQJ3oZoAzgdkneVg/ZJv5annb4cfdSlKapr4hqwOoVh2L7f+9je
EueU8WzPPYiAWO8wzymIYsBUA8GtR3mKyrNO3hTpEmgGr1liAHlWDWH8l++WnbL89DAm2oqZZ24t
zeQ74YLqLofF9iL+hsapCFANS7VEZE1cCqLrwvrvxfE4cx1jWB0/2T5gMI4KgjSS2ksxcYwKi5wj
zDLumJt3p7NhDEt5ZUnEzSun26SjlVevMbdYkT5PBNKUzfxSCpcCP4F94jZMNjLdm2JxUeH0E2ax
5fM84BhpNJRzBtx8q+hYAqXFzgveCSH2slxy8nbIYv3lYg/oEOVX8qh1jX5BBSLIiQEWOFt0L2i5
va+GIgFOO5xufPAbevBQ3uTFq0Fb3HE4bAkrSBnsJea1n6p1c3aWi2BVDFtjgklPRY9oCOZiEGSg
1tBB12pgCKGsZypw5xK6f/7JjM8Yr2nVYH0FssWD5Suv3mq4muSCq2bHFoKASxEbD/nX0HjvWSPQ
PxwofP2meM3pVt4Mp3ixft1Vl9LeM6i2NOzG6FDLlTeq0l+hNAvB0D+T7dbpg1hyhvYZrKG2AcZA
wUMY/fhqzbCz5OgDWGFSR1m9vWiwyXAiKu/GU6tidDIWPKQI2RgqRDDrzjPPadO3UDX3oiKK2ZJP
gEmzCHRhIjb38z8h8eyi3+CZi+ZbznbnVr1OxhdSwkjHTXBRWJAHpXE0/sM/J3tqBHDXVb1GU7bv
1Mi9+hrqGKMVNncLPctsx3CMK7YklvxeE2/I0NoF0xFe2gcQQM4JtfpuUVlr128bhLf7tKsRDZyM
C5hC+OxfV2KPyHGd6ENAAhmw2BYuP8MfXwqxK0DJkQFqMtCKB/CYWe7m9JMZSt7cHb5EMekXnI02
r65r/jSb9Ugsa/dSdpY8cFdesl4UCfihyxs9vlQSX4Nf2f+x4inWu/Ap5jMPzlP0XRS4KMhxzI29
JAlbUOFXUPRUPafjiLN3F6cL+IR3pKetYhqjrzxxpN17W5fa4YbZ9CLFw6Fs75ZJzh0B0dyXt3bI
D0aZfYLOx5Dy8824SGMHZlOm+fMaq6Y/Zm5UhT/MIRQR3UGBHsON873FYl+0hDxvMRAggb2IjcL/
GIr80mICFZGltRjMMpOmy7FMbFtz0BV8Laeane3nEaVAPzhDZkkEB9AH0QAro8dsNl/Z84Fejy0s
ElNvGsHEx0Frr9Hi0QxrMtUhO0mJurQ9mbH03Yzkln9yRU/qEjfh4Zkd3dswZK9Z5orV1KAIwbdK
hft+iUAVbyLlEFOAHoez9vUj+if5m6RJixvmoxNgZc4uQE6txAEGTY0xQ8DVsajzL+eCYapdZwuo
9yRXboNHrvTCW9otqk9a/aeKzQOmAzGiIDaXvHDOZtGiUWJuob2AKgqkztAnz+yh5z60TGBDoSrK
v1dU9a1C38nresBWs88oCDzAh/hdqHFWHsVAcKTUnJLQQlPiNGvDE6x6jmTlIbox4fH5y9e0tmPL
4oYpAstAbTcwJjo4EgFXFF9TwDD2oRXVRBjN/brIFuoAo25RuHjGA+NIr5MLcEa4Q712anxoXgem
u8A2JpyDzycPzOCkxZEC2QvgXz9xnqTo72265P/KYAW8yIxmoP7zRPe0KrKUp6tHQAJDxnzW+BXq
u2gSNCOlts5VFXJW+wYybkd+ODhUrz/eDBJs+VKBkBqLcgBitu03UepGBt3Bfj5ZGj3JRSN1DXtb
QCtsxpUKqktkBmyHNZycD/qQY/uptUJeT4Hv9XQ7j6X/lpP5ATE99/yRU1U0mlHURafEapVDZ7iJ
q5ufb8jqsqU8iy16A6y1sEFO9r77YJKHccckeaLCXAgaHHcqY14AgR9IS06fJV7hPSWnrxHyugNs
mEoa2prBY1ZVfKbYJ7qZFp/9fBsXD3+qJH2KvAMPIb/E+gakzO404QQB3l/BCm9f1QhJynuY7cQF
6+HYVldtw490gPjQ3T8dI8Sh7eFwco9BxLD6lA1q5akwvzPiyrB9r38QRVM92+0ckmvVQQWfmLn8
8NYsIHP7y8nH9Se4Fv7c3kI3XkYDiKoiL2RA9zg8RlzsJF/1QjtJVT0U8Y7PPjcktaGSKoSbIdCP
KlQvKGpV21Uc/6X2qL0GM55wFsnRmZw1py9jSOuRGGVQHM5fOCVjD11NtOplz0TdLYf+jlHWPaGJ
6T6dsDW26zpRkpqu1nc16uKfqsv93YDtMzaM2XK36UQLgfjBDoNR694iRTsFhN2rJMpTpeXxl/ZV
8iwz0495JugtLMSGFZifY2wY7Cqnk3dWnR0o6KLMrlDWVsTFXA4VkiYLej/7KsT8/lI2ts4bifEd
pYx+xb3KihAhi5ox82JQLb0dXOKeruvbkYj7VeA5wB2jHsvg9Emjjebxp9lPfc0rrj8LBhCewbim
YUfpFprYEmAJ5WFx7kVhi9nbJ1k79qeUpOAwRC3ZHKxvWRH8nj9c4cWN2PNbotHj4uBYEnRkM08F
cTzx+tuPhKPCNNKZJ962GJKw1VVkV/e5XmB3yQUZZj5WkeRGEei5NNl13PTtWI645do41CWcHyCY
CH3hsiAn37B+XrnlYMbhC49Rdj1STZogM5YNy/4RemWYFJ203K4ASUxiLJE7A19LEWZRUhYBzTp7
hEgeRQLkSknPYsfK2BhbOdunANx4UlSsivmOP+J9Oo71hN4JkBk39sTbbZ8hj3HsLPZbgTweR7Ww
EZzqP+6OVfh8z2WuRDBxDm8djheHVs9wdTuiPQ73lD0DJ++KD/y/1axhzeMCAJoOLqUl5ITjiPwC
OhDAz+DknKrcRT2hTGTYNTDshJhFPvPpj5gN2LlMa1Z3qaRGHCX8LckBw+xQooEZtPjtCmMAdsA0
y8VUlkJ7BpEXfl5/UjISr4VY4Mn4FKNvh+oDBnGVZTtKgzEuljrCTim/hybl8LbSss+0oWX8gSBI
hLaMcBhFiwfGQ06KC2KHEz+jl7Hk9hu1KEPfJ7jZjO+Zp3dl//zAk1f4mVeG22BKdfSbysko998d
E/3WoofQpq5Ueb/ABsNSzTttOsj3A37GCS0L2L6y693Zx5Z70mHNHDV425n4wHJKz7ZmbL7YYa95
ihfA99TZ7/NmvkOlZHak/8ZcOI9kshfkZ6v0JXbZv45fI4RE/1HdOM8HBLWO82UnaV13QatgcVBy
fQNC7O1C8B6k8wA33+Pa16qrADIKjhelp3d4qna7hyDKygrJPkFgWzh5OEZkajsm1v0LjdAoGWRd
i7JGMOJrloAQwsymvGf6YUJFcIxg18/9N+r4Spf7RFugAE90SjkFu55EnOwrzKJ5BI6EqDYuY4aY
CtvzZ8gWU7fU0ZfANTyjXgq5QWgNCQp8r+K9/Om8OM+3N4PmRoF8zzok9sHqMxq9T8Zowqdg1HG4
zxQDTVStIfJPCUoU1KxhGkqUNMvaMCHo+yHX2CMT3EI3woI+E+HoFpEBRq7xQ/6u7LJnbxGzbO3w
QNGYaKSehSiI7w9xs8QtlWKoDSBQhNXcchjj3OCsj82LunA0nVyA4eECLvXWpXBxKCXpCcf1u6ju
4Fc3gK8YrBmIAxUrQyssLhsZcId0qu5L+U/HVkVAto4mIEDx5jrJZjjMNNwvI1HTUw+v1fx7F63F
a/thoTZqZtgHUY5cZL3KbXdpqfuvlFWJSY2TkEAhwe83c17B7utdQHfPpuJQETScixaAuat1KnNG
sP81lQGSLqa+DcTVnHLzRI72yyTwIwyqeNvyVT1l70HAWdd/ruPuqNnt9BKhXF1wJNENpen/+H2l
xnAq5sxXDz+7nzBy/xf+xCcAMDPdC3Mk/pKIJ3pf6majBrR8PbBRdH0DirbMFe/dQnydYInorRPz
gz+nOlLlr36zyZyRZy74fYREsRywmtosG0DiC4ofO2/fqFXUbz7c+ofFHI8HU3tSRys9BZ2410Kg
AI4bF6igmCGUBarSmSMiYy9UEQAr0Uu6lBmxAfGnkGmQWC32n/X8/MxNK2UAbvKZJPv40vy5r1ce
bkjYqO/Gp3iFusAftDKMh9GgMLvoOPU1Ao1dHdosCN0w4t91e/aVRsQ+7oxXPS0xU2+qOPAquzYL
liUhiRVjzgJ/wqmX51vkPC0A9+vQFxHsVhVongf6XbQybEfJvC/5YT2wRpJob7rD6EO6+jCjubGI
s8MWaw5SRknYCvLltQUAWbKGRZ2EY6pVM1Ol3D8gRCCetC1YILRiR4WNdWGszzxXRYVRR+0127Gi
JBHLJY6YfwBoqmaba1u7yS1apyEY5IB7Ax0OzgDY+taU72zo9yO/DR/TbdBbUIk6QdNf1bL/4C6A
lCxYnALKCdIayqqGPyKKmwsuMkgUnuLkaamvzaFmfxzymyQCG2iFvdS0/KvcdNrdRgN1O4elU9oj
c9tBoxbJ05Af3X+4aBkWkm2kNL9LKS3VriAU63UCmyLLzhmBxNoV8VV+HbW6TKjOO0I0GK2Gj8aS
AakIWkH4/RCEnieSrmeoOcrBwLAng3Ix5wVY20VsNGz9TSGzgAZcIxm+k26w1sEmhCbACCzf4I3p
D6a+Z9BzAUfIQYEUptArjMVqA0YJ0CfBXq01litMNx4HNzXR+YLndBjO7U/D5Ua46atmXIo1wHVB
PH5OW/8LKnnkHxJqMrkPcnMAtBOFGlIaIlN1hil5YfSrD8pnfQ/DUUE4EO9X7UqrbJZhfa6dptCf
t1d7wuRFBkL3IX01XjRtxiTbIjoDJrvJY36aM7VW5NGLS9POCmJ1W0ZxnluTAtkdUA32AvRxM2vS
7s6YE7F6wk967u++fM4HnTbjHCxAmBgfLJ52HPwOJfGDqDY0lwvyXQnUNC8D2JAn/tgKLad55VWu
x7B3ehXF+eH8C5uq/g416PxDD7zpxTQxNO7015xdDkU8AQymQS16D/zFksnZRfNSRtzmxgDREueo
GnbfSufn8tyPYv8z1Iga64QmRj4w+S2GKqGGElBpyvfXyVLq7uWMIj4ktffOjPN1+LK6gHhmsVdO
fkzWd22KLQRtQnnSyBW1QUg/ozEmsW2PupGf6wh+DsOxu/G+ygyWcZ8/IIEU3g49F/hr5+fJjA9O
69DPhCbQ8yPR8UGMCkKRScJGsUH3gspgA7QCQlyEJGquvOPsl0paoUnHT+LsxBxlZGC90hlpvnzf
nz82yjZAfPDplEPUul9xudJSUZd7PGsqffKFWHL/aQxxbDZ60bmkOGORcaAOOKypVvlGzV7itBnA
/tGObSlE6SfunF4RAyGZL+UzMNMRYfboZWwEO+JqF7KkXhiEU5Bdf7XvlIumfjoNkTUz2TYOcPjN
JMWb3bsJ78rplXGtKdGJGTwmwPZ3OEvUy5H240SXPJ5cSl2ZEFlCQshrN0T/geOS9WmchWtBFsm1
xfFhLlddaUY9DbHBPiJzVDRqfRJlQudHMYcZzF4E46TPVCWp6XGqG2w3s7aIkdMKMqp6kHzORZKp
zItU1mqW6TZdVMcUm0Tl0KtIB802az17noySUTojazpZJIq0O6n/Q7FUlo7pHHvGqNTNOIN6MHoP
p/MiAHK4FO2ZIbaqcqy0AbMAMxx7O4z9HlO+68ziA7QvktPxmd37ruXVB0n1zfDB74rO3pzCi0KR
o3PBPpb/kczKIP9SQixyW8LVb2Qxjn7Y5XlM/ZH4ZUUjqc/89+ONkE0HcNBzy2aRU/ZOsJYbj3JE
4IcTVDZV8SCM86XubRZLHiecKS1GQZ5x7R8D8JmurftrFjLo2/ykBz/8pHRDa0LFlrP4abKOIeN8
m4EIsqO2O79QZcn6zCmo9vdqkF29vrVT2z5oFexTlBI/f3FqXA7skfIgxwjopy0+FpRGX64QxzVM
BAWOf+aMHcJdnRFXPd5AKjRg1yyYuGQOhm2y+WfQL7Ta9c9x6t+YHmjuFABK7F0IED0RTNhrYp4h
UfPP6eGOTATflkwOuwIZluoSXcr0CAf7AqBiI6vTOf4AvyFrGw8n5WDo3n11AOYv+Pnyxmo+7ejO
UsQnJh3AD8qj2nTk/4vCeL3lf0A072n0KoOzRy2CSZKbW/yqYbYbHaiQzSSv+QYY1fGNX+U+wLWB
gEg9QgNhCoK8AQpi6BxyialR2tPnr04d0t5kU1XbxNVqDuL80+5E/IxLUY5f/4kjjlxgi3VxeQyX
E9q6Bs04AKjImt6hfuGZY1qNoMlAoOM2CKrS5Fq6yaSwiJfpnCaVyUWbmVkNdUG3pPG75Td1WV43
XG+hYelbPugrFe2RaUbV01bPHvPiaUEpAwTSGSgLTjgSQZ9P7f4fHX49CV55kCTR1uACB5/h+99E
CGuCGiV52rjHP8jSq0GEdmDnD8PKjbrzrhOZYrBxGNZvOSqsQSzVMBBnBDaCVMqQIIqWZnfyB4fE
vs3RwE8fz9ejfsQ1ZyFT2nsGl69z8RuHHm7pculZwzvDn4cZAUFJns4fWVm/rdiZFMLUdHAdOFHV
5T/vSyzNwfq1anQHnJdQ4y4CDH17CUwvK2Jam+aAsvnlXc5CD6yeozRsh9/0RdN4p1xYkk9AaEYN
JyHR1WffusZZ7hIKNfj73ZwdHajVqcXzdRj2NgZwLRLORxLQnY8wbcgkTJ/MOF61EEBZ4K+/Y/uv
+wRtqoQ/iaFbmqFQXjq8F0x3mG+NSenq2IKiRRJqbBeSMA2zZinSE/5to5xx+Y13Z/quurBY/Lku
BINn6if/rbxBvyiJvPzwaReyGG/MQ2/Nf47zbc/X8KJ+656r8BHGJmB8Gpoy/slVo9XPBaFnjlbA
1ROaN8YKqR8EXZM9LwLZO2VDMuH1JCwc02bJCEIOtnHOWszuKhtBxM2oOkhU+mTk7Fll+BDnQfYd
yCLkijs8CFPYJMpAAoBQYwEeoZtOxrFeY7Wp4XClK9sqCr5kU02hwXkEECWvXPLhCpMKhtHMPEbH
LL49SFZs1l7qADA/cDAol+tDlAA85DsCoPWhsvqK5wQkPhubxwGOiSgaYJyEnkULyT9528V/UadU
C+b9EiRKvdN6l2soDbacdmPDVi9n1lhceQh8/15/XpD86xpBXakjBuwnTBjuZxg25bKmpiQ+U2Wd
XN/2wtzumXeUh+85cJLn9zbsJ+RI2ZEyJd6H++j30FH0Itjhkv3REtYImBfkgegfg/a4zDKHkgbe
m8oW2QnFqe90gTNcRaUYpTwXZ3LyBGwSWmqedlu/uEUHldgXzTNHuLHkmztSWDuKXeudFBqA8Gbr
D1g1YhFaJ/kT/gKDQb2l7scgZ2E7duMwg1sMuydWNSG01+VOcMeyWu2l2oqu0UcW7CUcybJ99c4D
I3CiEfS1n5lDHE0ADA3QQXKL2P5/D4K25RtEp4cSucizqf3zrm+qBBdI3Qz99tDIMLygqBpXnBSj
7UDUASC+JBULgs0qtY8zGIAx5bnFhfJD8aDwuJkLGCbH6ooZeNi/7aKIVAVOLnDneuquqIqbmX8Y
QEVZb1qRR8qrOCh4KkBzyUqxe9eShksDORT2X+GWqzLT9W6x+2PfyJM4VxFb8BdDfoXCQXfrRV4R
vakxhhADBMQQT0iqg09PCKDu55X2t/OShTgBNOBJODo9O8flCmiCaz3cfG25hVfU0QmKf5oMArkX
murO5zMRQ3kYH6nUCaQB+Xp1MvN401O+y3BjLlVYWeaDZjbgXvEjeZEM4GhUBXM+UYrYrofVJb3I
NtkK6njP/RUyhyYqU0Xj7v6S4wwgXO0JuSt0gdW8Fs34cBveZsOf3PGB+X4U6oebtHhB8xN7tlaV
ta8C5f3fR8ItG4Ek17YlMjK4XX068FNms3+WbcKxiQ2IgWziShd3PBVMcapttcEHQFouRmi9Mp9F
AG2UL8+G2Xs9n5OKkh5olC4GFT41lUBkl7IyB4JxNclRuF+fzsd/2Br9Z41QT2snSoaOdDZeQwaJ
FUgGzYrvmcfzonN1PWmyNzEyOxxIXXIZU8coFYzhPi/Ev+LUNTtdaOOYlkE/2k1dHoWNrCpgcOSn
H0Ma+QWAEW8rBmopg7CU1RHfm93wM7yG8I5I80npP2xpcJE1dUQBSrkDcuWOVMRFXxvisNn1zfbP
H/fPE9l4UaJVmorTpXB9bVmPYST3esQHCYCiiBpGG8RF1OUGzn4AfI/IfqRXAnk+p1XX2xcxr/Dj
79vm0xZmsBAw3mYgBh+0igq/BH6j4MOsOUMLk5Dgzep3326dw7LY2jQEQ8JAIxapc74yLAwgaO2C
E/FFBZBFr9ndB0R59B97f+R2qvy5k4QcqvmXq7VRXVr1y39mjjYnd4b+CAhIURPRdbA9zSM+liFs
dscXB5AT7NFbH0WL0ByTFiJpPM53PWPK7YPG7bbVQSzU+j/U0pddoGxFT3r0zhwKoDFkPpxUQHXu
aUNCfIlWvT6ADLKmOAnEV4TJxgfb2y7/JbgQp6zvpX8MMl6JpdxidZm88BWpp+xXnKhOWng3pqn6
Sg+DNl0I8+I+kL6WRxjLnDs1EtKQH4xDH7LemkxpoHzaJ/YNru+OmpfHeMqb2AVJ91IKGobBPqQ5
vr/Jy4RvdvhmxHJCaZla9S2EXKMYL4ioZXX3CSQxAngEsVHiOqUb5VGU7rYimqsHf12T6mNTVaXK
NB1EHjZPw65lQx6HidQPmJNrESQUXhT+X+SsV3gPK+UnM2CoIqwZtpQveMo5fhw+qI/rM1Xobh5C
vkG86EtQSYn5KqW/JQU2SILJVaMcgPJsJ2EJa37WhGFRTMfzwy0UEE1Hwf2Cd+7lIuAldn86TF+e
X9BJ7L4Zzq0EOkodhkW4w9gqgUVFzylg7ktLmN4DhIDfc7KETwxgBhUZ1NJreBCzFRY/ahvh2cGF
llJj1gyKEEkumFc0vDF2rVyoj+PATP3l3ScNZvxXeoy0wPj79N/dEnQTd/wgXaxI14FSCn5uGNFm
geg1lEmhKIrg/9f9IZ6Dh01N43MzgLWNrtkDUAj3pb7Zk0UkyNgIAE5ZJGGjU0JTszYgN13h+B9y
iztG7U6QK0kzd18AwIjMmW/DgcsmJ5lF7Wh1UjXUE6F45GHeIGX9OIPmpTkUebzvO98WjDoWXphr
e0C7veLiqhOCtmQVDIYj1iONYfw0JPEXa4+QrDStdSF4+wykj/U7aNggxLylbmsODObFLrJzxl6k
LxroUAIu3tfFFChVtnh92SZUGmDiIed8xy3vEKOu8jc0gaQjadtBoOlVeomE9XdR0pyxPjz1DGzU
vFqdvGV5imdh80i3JSBr9sKMMkfE7rb4Oqz4VyUefvuWtBy1vs6++R38lzLDLBpZ90hSJ32dnCic
0lKLGVvqbVRsIKu8y0nS6jjkhAoPUrkj2SAORo5gjc7UeSc094+9kXbT+ZbYWpdIJ/k9kpKydAZz
NVoUvPE6LItvKuanBW5A0H4uVE4eAThvA2DmPVrd1T4ntaH7XlNktb9M+txx/2Q0xvqgWT6toQls
zFs8PCzDea77pESlfXHaDiXQfSTJ04NE4hhSyDFZv9FQhBaEBdexg0oZf5PU36cSJIkdGnrdjOZF
28ItcQ4yAPzTdiR9fkRK/U4kip93BFSIHzdvOE0uqscLa4AP7Qp+pQuUMFyoEQCNYd51WNfkrjFJ
TbqaowEygvC2u/QaTbedKuPNC5NPGCUcE1Fzew6vwjAbgXg0zn/YrSwJzm2CBempUbiY57MuqvMK
Czbl43dM3u6Kz/OHkbouleVL6lb2n0GtgBa6GQly/S5BHWseMdmu/MDLSU+1DcFzRNOUUiNUZPJG
NUO16E5hf+P9lloegHXkeHjVm0rNk1fP9JDKgs2xSrFhtDBqus2tY+M0MKFADo4DEMyMDRFaEH0M
oXy71kUVRmlrhx4GALSMVbJ9acBrOHdgKYXgFZffkC4Z3LXhVfhFRWIcM2kUfXCH/KMD2iMCEZXb
WOk+lSjO3GtKlzBwzFeb5x5vemOcIC3AP0DrfR8957ockZbLSc3PCP04aB40c5X/Y2vQh8TuGU77
2DY94RZtNrkfgcoUk3HkriaZr49gprbgJl177VNUt97Kq/JWou9a0Cvc6N6CUgaP9MtUZqi6Ar25
ayF6rz4m0OwjGZ81YwEcvDWDL6rRAdT08KC/RRBttxGsR2PH6/p1T7ec8DIavU11ZDQoCYZ8kg83
A9z6owuR1TcoEO4yIJ9saK67bzWTWD9BMaeUi6Zcg0DJnondMqaLxHwIK0PRjuFNvtPoUap2VLbg
JnlNNrWHl8ICVX7eigQ6POrjiPg9c1puRwvGqo2FIk9PfohjtHTJFVSsPYgv6qRH1ekmJWOVOFUw
Cow70DSxycGAhnKuP8oSOSPGwKECwfxRH0ZWUyxp0hD+b8U7Q13mLlBYUgVuoEzBbZjJqWWq11aA
OGbw9xtjfb6TLLQGJ5/R8GqvAc1MmhDTHwMv7dVTW4kl+qe9gHb+bhThGwXza0nK2fFaO+EmJyHA
mREegGCd9w3av9HXBPh8iVwrF+dfY/DEMg2cYi+pHcW54hlxXCwQJkiEAL9Ed+aVFz11VF/pel/y
dlKG4ZbeWxs1p6m8e9E+4af2XW9sWCHBNbhop2c0dj0l5DgNoqpTHz6lAZR1mOUuiSXnCG4hCAqV
joH/lnAWajsExDil9Sc5zf9fideOhi2E+wIPNk8sMcVP/sFnAFR+gXSXU2WI9Rj+oVkxnB41oQba
S9GCOSQFxdWFgW7korOc3iZfDEaOM4fabdTQ2zAJlY58e5F1Zi9quIbepE3JaAhjCsBjOuGOsIY1
xmnEEKpGxpWEYaJ2bBd4otTJXcXuojMJrt8CUYIvCOt1MSsdGTrTXc6/3EOp1ygFYrU973ZlaxlU
04T11j0eziQsQkMbqMQqSqHnpoE4xEvZPN0BfdrF++mzd9LTkAITEyP9EQAY4MxnOfOa8FBdhAPc
+FZRfHpfDO7veobmrvPvf4rNmH2HY9K8OqVfOGnpHTnCNMBymMbkBDXdxX766jaRk0lmsw39Vs+3
4ocQvqi8z8kgbJxk25DZHhtPdbDjxC/aGjs+aHh/YNuDBtzHjDvlPLa70w87iSbTsCf6dekl4cUq
7REextljb9KQ7KxPjKwJMzbpMdkQnNthPhYlhqktDudDjBQxJWNPDIRFeUN3RBn1OvF+0KhdMRGX
v4tgykgh+Jj3bo/tRhg1a87k1DsxeDZh/BqyuDCWoCfTyzA0IcXOmcfTxSaH4Zd4GlJwskOzXdTz
7HI5K/I0+dW/vmlqMgIO2HPaRcU3h/Ch3S5ZyMV2VN79FjWSRtl/qGWo7ewciMgvIzvYxfPwLU8G
ihiLp6d96TQit2dB0EdR/iI9z9rNcXCQ4aVAM5s5hm3puWkrwt9gsRDXa5b2Cri6S2UWWlJC7VM5
VAiElbR3cT1RjeAEbPNsV+PP1NU96857YJhxR92E9Zfv+dq1HcDnwVw7XmyCTKSnSgWccTb3c56A
vkrTqpdNLGVjKVPL2JVEWCooNu5eZW8SU0mtqjkbtqA+2GQu9/FTA/piy6sKXB0k0tcr8hCCwFF0
DZjjtIxNb8YR0th6W1GSYnoqywVwFYS+oVaNozpkBDcqYVLyKMlFDXwOIRf5eplt6g6jy8mcZGu6
nMKZCwtAwySdPJ09V4sgufWyerXrNzT4OrtH61l83QWgBzPt3OtsarTDqQmzZeIm7K6maFSScI5L
0xKkOg4Bh+x2rrXqt3nesrA1bKmFQnneefIhT52MwgHiqZ4jn8tQs/8DEGAyaFfPC68td5vZD7X9
9SJ3kPnsABrfNrs6AxiffutziLlv6XIvZnhOypaqAHRrkcj+7dqQBVfQ9bI5IVMnGDsbko0oe/Yn
mVrDaMY+JlUTUq1g1NftEFuShsZTB8fVGQhFVb/dLS5BWD3OxR0fcJZo8E/XnS/RK2ukmTYe21gz
I/fAVRzHf56qknaikelQrDP8WiHI//os60fSM8rc+SSqYDG1FksV18vJgYIbPJLg08JCIGEwnkQl
kJ5AEvHZR6XUVM9gx+XY5mCQe1fh6NRyNf8uCEIohNBt3s2rwohXlT5nUjH3E7VYBSu60XmxQ0Xo
KQO526NDrHFR1/7iHdgGNMLsXcD9xJ+nn5mSlht4LQlML1AsXP2FQfTVB4mjh2IgixZWE+36IZna
KFR7VtRMZQGLqfB3bVmvoXjXVkQAXR8fQonVE3ctr4h2nKtj5TULf8bJBvVvh8mSY0UvJEnphYfJ
oDvnLhfJ9AnsZ2ySukloypgS8oO2XrTPB4DKqNEs+UG5ulct26maODE1hBLlUozULRtPvptptOqc
49tHXVbeQmRF51Dncxm1OXnkyOTBToiDecCg/19cH2aWLXTr+K5L1uyOEBZ/NP68McgxV2sggI9r
Zowxl9T0cpijEc9Szr4tSsj+TlVAUARbjrQXT59qshyYsqRLr1BVxHGaaWTevinNxuV8gCG8wSMM
1Lp7L0ojpG4BgWdIid0jowxnVfIydFARedX9/wlcFlVEpLW9vrHGMmHikFAEk7t8D5WgVKNbIeFx
S9rzAYrivG41Dv6fScwC7cIjCJL87EHzDvkwmYl3K6bSGCBUwbXBTu5NKoo+VTKTbKAlGVOf2laE
Z+bzwKrr7TVHxvYv9qoN9CyPPy86a6oy9hEoj8QGQu+5Ka0gn2Ueez3P4z+TRf7iowAiLQLL/xvK
8lBkJXeJ9z9Ymly4aysj9INmRdJNPDY9XpVVj3sM6ZE2mHr0UvmmQwcgm1D4tQ2wMZBj45wJ4ySS
2+fsR94BEjCKov0bbuLFFJSaEH7tylxWk9eU/2KzWhsRndrii5FuxMaUoqRO7OyQ7cQOlwCA51UT
L9Tvb1PihMdtlQyXfHMjH5O+Ovh+7tKnb3SLHuNx5vkJiWu6NKNc3PbeuGHVY96T0MV7Ut7Gg4qq
g0lhYHXAzFWvu0NZoJrqUkyqZu4WRcjeNTm0qxzouSY7GstGufB8PUQJvQ5vQ4ULf7NSYJA4xHFy
xsCt94BRonJDCUw7gpsv6GUbI6cA7n87e4pzgCKlOvUmHZqa3sDcJ5EPXbJA/AbhhH78RdZowQBh
iB0I2LdBPI5PFhiG54pYHXWqkRI7flSGr/hRBKeS9GHiStQDnA+66yBWj7SH4H7YPdTB2CMSs890
LYzARr+N8CNS4nEEqvGNWyHxco8VsUQsFTCk9mDEWEnZjzujYrG0g6zPjVL0CKckm7Nz0JnH7Sjv
F3LHrNNYyWjI6lvvHWNiJS8rwoA0TxWR1UwpmohK5kZYajTD8tNC3pJoQ4vWquB+3T+lfwcqZbvM
tu++3X2OaB2F+qwKKXb/+kl8YPGrqrALl9frJBZ7EjwoC3Lr8DoVTkz2pSxwvLF0+Ta+1iHYKFn+
BNbgS3TX6QHJmyAuw7uXZQk3Z4GRKlbD0aibc06LzQYh4uFTCR9nMesquzGRDr/SMS7dW1ZkDYqB
++Un3pSRCa33ntrpY0sWhBDkUuifQJfS5OCDli/HYocT0vxVBwWrb6kQ93KGhgdKZS5rxqkpGfFL
mIO1ef73onJ8olWV52/+YBPQHPe0IGPCcB7JYkfDIvTXCpraU9SXjopbNwsx1T/WYK6DyI03oQiA
O0VqiWPCa7uuUe8I6U9sIIHuSxl7Z4tSxy+7k04NTHXpj/TLXiNqzWzQoyCJFS3vGodFHz/VN/t/
VhauEL8Zogkifts0yxn+BIOBwUqQjotXZS6Zbpm7IOGgwCMzVABj2DiBkz27kW8n5b1LHNNxxwtZ
b+nYU+6K55HDmz+2XCI8xE1b4wHRPZQqGZtNoqSJwqdgOAnGf1FSYifGSxUkBI5aMCVyPo1Cc6JK
QTwpLY4XdJJ2onvbIdyVxZCeJF6M/SWpY86N5L30fFtMlbwz5CMhiMtU6KPrvw/oVbLxo2kjEacI
B3DBetsHvBNM2k59Q2e7kyRn9CSfDxUgwJOVKIx/rSQnniYQdgebw1PTPYta0ZLoH7ON0UJChiup
IVpr6HlrL5qTmziVu0N9jzeDY0Xxxf32bQZzBgAuhB9BuiVQyzST4+meWrf+AtRmxsl7xHeR5mdQ
sR/HoR+EnGCkGQ6lpABCivnChSxO4CpayUtVKRODUUSTaU8ve4snilnLx9icejK77Mu5KA3XDcd8
aiEVMGF626r7poslsUMhZclZAX0JAfzhMXrLYTZpK2B/Nzj5YaMKAwNWNWz19JcIXTCgvB8llQnA
/vuj4f8EX3Nx3Sex/cR2uONi7AUGYt++YNPbhmXCGjuAdiA2UE293YDaAdejwm74O7N6UQ1wXVHH
EmdL4kZJXT2i2a6Q4isIGfYEYerR6FY58R8O32rXyAOr/1od9T8zj/jlyf7YfYE9393jwfmhwzJG
8Vx3f7EXzxMqUHSFeJ0mLD5SWFO5ukYPqdNs+B0sip2LrFYKa13yvbulRgWjtnN/mOczgX/4TeBE
h7HqoZm7He2ullK7PyK0Y1c3G7TevIXhwjayVsP7C5kKEQU3QJkxkck8eZP1rqaNvLhs4MBHJ71X
1S6hY2ETI0mNibn2g1WNxdP/jJHPCztZQc7357QG+t0yWW7PXskqNIB++oYH1D33cs/j0ZbpNZk8
EN/g+jZXl1wtx58J2pz4egXLm66X8L1Ivx02eyKzbTM7eVGufwesNFcvl1sdJ6QrlXVouA2oBdSs
NVITkD9I1bHMtv/694sMlcJEQwtx+B8XXIiqDL0i5mK4jYldGq8gslssZxMNOoAUeeuhvVweTVH3
vTjeVh8uqdd9h0iS6l4HeWiqcIzdJ89CkDkzen0GOo/r1kWZcPdnkagRbWRsf2o9oriFiErMPIFG
qLyT4Lbdl7RYUdOeUqWRauiGUH50uuizWQict7exGpBdqdpYx772HjJA/wQLZ87r4OxB8iVuZu18
1Rio00pzuXMGCk92dEeWRK5FOND35ppva/v0jn8OP4NFUhf1jI09F9R6qE3SDPlDUXoqVo6bgnVx
IZ2GwXBfxt14YpJouUxTxaXw5mOB5JcXXnguYUcramrd+XtsWDlxCJ0eOOxpH++8p8j5E4fHy9lK
n+Ngn3nJza17W4+nbTa22n5QICStVyKBpHKkg9i8uezE0Rf9CB3ByP1PbIWnmATX0F/nxEQM2poP
6vNxhCq9xoTXJz8I2lZRnlXR12+tyqqPT+PeuM/pA+qGWGKODC3LlW/WWApkX463icLl91Hy2Vc8
4D+ISq5ZUEiomYbZdUEgrshDh+3BGPQLO1FyV95/d8CJ/+OPigazOj/aPqEXGtYdztOQadZboEb6
rfh33BawK0N+wu1XdFzHj3SPVkavmHVGaYaxrqCSPx5Yx31QsOJX8q6RUzzHBgYq61rrbYxgRvJL
U9b8RCsGoNI9dJCk0vw/4g6AHUP3hFy/YGlsbtyA5YPH0xf4Y83lf0cWbrQqqcaTTdV5ZxHmbIV9
u2NdHkBqPSSYt9nQszArhhp+kF9k2gfH6Zb2goifWSxcmnpiJRVuTQfL0/JTS7v6F9avD0xFu9aZ
6PeY2POII6Y2v1XeGO+ohfEO4yOCQsB3ahtbhKQ5/hsu4uLq2c3SEAe5B3Rozal90lobhMyjjy05
eisVUVIgT6PMX+IiNaWsQVeJpTmxQL8HHL5ZtO5QQVno8MQUpsde/iQWMaT+2BN+vq6nx1Um/wLB
OsVxKMYwoWl10bdqxvKiaEvObvlb1LV8TW8OcwMbDXbXcbHMWSordE5X+eoq85aLivB8CvIlUhb2
pZQLjSgDZcw08nJ5uCVx3bdCS5/KbknsT82CLeQIp02dFgI78Ae6mTGgfubIwgGUb0k8NUuhozj/
W5wHyy1R6DnfSmNxle8iE7ZP+vFGs1Q0Z3QOnJ8CzpAnkRFQMB1F5e3RkyY1XuomBFImS7jA9XCu
gZuOPSzDUqPErG//43cl0Sm+F8dlOEP7sQcW6xxlRlhK+UVlXZkPnBBr0aeQIHoSu/USEeqXoQ9X
QG3LIotfZxU9qs9wsgXgYTN0okGz085OwJ3RuGDppsju0YCUhSv3PFx1hSOZhu7T80lncMF4+pKL
KobZE9L7QzCtW8ajtKLKpe9YNSjR6xsCnFYKaawugCY00QlsJzac6f9318IjWadmkCX7GQ8QPepQ
69a09WQJHX1MLcbvbd+KaGzHqAZKBpTw1gfKX/dQxcLMUckZFEwtDpMTH9QXRBFiOnBdCfWP+c49
Kdn4GDmaAM7yojEUwHmRalK+CVfJxjZhZrXrCHIk8c15VACL35Bfa9BE0u0ZTrTLGpwleQRliD1W
T/K+oAaXhY+E3cV0DprZtuGmonfyCawvKmBax10lJZso57lBin7YlVWgnVvk+Nfjfj0ucuB9LS57
UB+azApMmK41wyabc465jfpLim7nyE0xrr+8jLqHI7lkPslj1QnyPHYy7FnNBLmdb6dtg+WQwPdV
AthIX97QXCiDZdlOJj9Tmz8aUTZaZ1ZKpY/7cgqBNCE5WymWzUFgKfY3zwC2/n1Y41SVmi15kOz/
8ywrNaX+FZLgushPVVBUHBkwfdL4xVgL/Cuj9BAgTjxvssNSTFgyWxYGHj+/pWNxAKLeBUiKPIVI
5tTciVQDRuJKkNkbOvzLIFlkULjjYQvUx2jSGZBTAn91g40hjR0FDxs+maofUOfgVuGnJw7Cxhwv
A1odwHpRm3KQS/GcjHtSYoMoiKubk6CkRTYyUCAmBLMDjwZ+2lg470/pbVnRCb2+DeBAvbkutCUa
umcFoZ3Nx0EkDs3d2sLnV8KRq3FMJhHKstgqhrNrr8W0KDfshNBrCHn2oqb/Efocy+THi/klDg9f
aRDZtexnp0CcerSyx2v96v0GBVXiygnMbg1DiLAH4Qu6NgC6bnblCzzbz6N/J/BBohtuktmtxwwz
DwkxAO53KGicxb/vI0Em0yNxsEdRgNaplGpxxkKu+kh8s8vdr9Wi+s42I0+l62Py4/P8d+CDENKg
qjXwOhBG/xtBzwTRz5g69LNrO404Li+1de06D27bToX3qvUjgpTjI+y9TmfgROEgADN4kbxjxbFq
kyI+wj1n7Lz/9aXF7n5gLFfk/guvjm49i3fWrkiwyeoT1EDxz8eIu8x5Qq4rpGGhFFkLHtWQpzn8
bhWQh/phb6i/wL2jicA+hjBiYu/2RAmXhcRAIbN0xXn5H318ifRuEMlka5G3/MDZjbXErg02AzIA
lxsN2iX5LLyqFSx8GcTiFmYztVjVIJkWQcbtjayhos4YvftbVHbHrI7GIl3scbygZL6DOYcdnJvk
yCl0jjiQ3AydCEvXrmdbVU0l1h0ReYW3WJbdzarqJ80RvMvfeqG6qiSIQpSPJAvmLG9zK0guklRS
nzHdgMS4gv4e0MmLB1eadIbtt9XANGMhlUlkA9JkrzNtoFo7y9MC4FoCvwEleEq4CI3G3A/QCG4m
qSTe174+HzUw+4qRQu5qKIeJBDLmlUBph0iBltXXSGYMTkOEjbOp4Bkl/0+xdYJGwl1AwurmlAu6
AupLRm1NPlxIN5N1pWqetzj+/5FUHOMXS2+4GPHLS7cJUpFyvTGNK4i70Cm14l2YiquR/nuL4uG5
iKvgruGfVa11fH30AgBygHOXHWjyFhzvQRLdCyuGjkwidMUNk7f3k/in3BLW1HWxxXHxKJ1p5GAL
O+EBUvgWT1qFbKZJJasbpH9CcosXGX35YNtU5kwU4YeE07yZ8T0lbxQw1F4DbZ4aofJR3LDEykQc
Wfdbm9qV1quF3EBOeEaCcb6XPMlQI/83RllAHgqF+GPdIOLTw2JLdTCQE/vdBmJ8WUTtRaAqkLCW
wvRoiiGpb++SuMoDm4be5gVv6Z35pNlW6NrYQtg6g4F0MC6dyxcXb3sT4kvs21HkBwtoh+FWwsEv
jJKHx6bFW2/9aEDipzoNTViqg0hexfds+8bwrgu12M/uhDeyWuSIaXh68wZbXik9a7A82nCdeQWj
5xLyzhMaVcEVzUZYaxoBLkcSdvbkQZdrpomqqHzi4kaYXQPBeu9Nmj8vaqF+YKdqrK0z7VeOSCKr
ODdMbR60ie5pzzkvgJ2Avx3SG3h37DoxhWlgqO8CNJjHrv+Xu3SbJlA0No0TqmYne2N/gZzTAm0b
u3F2Dx31Ws7qkusfnqXG8Dy6Q4MgOj9LRCjbtEsBsmQkgMXpZ3kIuHx/PS6qCvBGT0HNZyhXQtI4
/Z8R3xL09yNAD9gStzjVgM7pSsVfoQAfUwF3QoRFz5tYdrbRb3478xEHNDCgI1AYhhqYwyVC4Nmz
ZxQL1DbKEXk4LwgrKAVDWoAqglEkuRvgYR7sJmN5OqyhAJWs/r1pb9TBI/JTESLEObGfcTmdWCHj
yeacTFg+TNhUOGrh0K2B+lrzZAq+Lbl8ggXI4NaKX7wDfqsmraRxCkJvgKUl+RKhN+pTO+ADmOar
Sepg4ZNtaDVx25owt6Fyj2zMb6bcw82YlAI4f9LzdQA2MzUwseQdDMY0Ctzsolpd3tGs3jg8dSq7
m06zG5YBQ+4z0oNh4BUi4CNwR7dKakbhgTcJzfpnrzY7DpNsC5zo16bd5ODeZUsSfXB83yKJVQMT
NlGwIhe9cQFHhdmmPY1TW2GgkKDvO3NpmmRql7+WfOX5QrHv0mE0jCTQXHueu/VO1ciVFKyh+LMk
hlsQA2qod9DCD42ic0iwJF7vB/H4y+NAuvGmMSi8M/HAvQbS2OACnCdSn98BPgPSv1ZAj7G/qrph
gJpi4VtY+oNSqre+q6V17FGPlPbaeKjYbcVlfM8yPKz8VV77PXyO6iQ19GEB51vlpZvlmRo+bi76
cD84Fkmmo+TolFvFi58zprp4+xlm2YzGb7lvhvD39ssEEb91XJwun8uUaN+R8M7ODfokGjGpbccb
qKaeVphk8ptr0HQiR1D2nRXzoEsJkAFZd5iBdIbVq5C5Tj+Hf/vJ7q8AFvkMoHMat6as9oGx9A52
D+7akoDejkFwDCpsDL4LJn6fa+KMFZYuhyd9baW0dnqa/OWM87St8Az2EtZK+N38cNhelc17j7M1
TnURim/znNuYEAjRfsfW1ObzcmFtSU2pf4OAjmQVCZYx2N3Yk+EutfJvjq5qI/EeaJhC9yYoO3ct
MJsMpk/IDLof3uJqHLuEydJPWR11R4LPPsv9TDEuV0lz/fZN4XbGd5FeXmToPqzNExtK8aEpUpVt
hDiN4v040ncXo/wkqzFwQEUpr0h8OaVZi65nJaIGtOYwNJqCvnO5P+zP7wsx8fovVUxkupq9mrfj
CjJoUJEHmonx5O4CSUx9WxAm7q5nYxqxeIsLRcRRre08B9qv7UdbpCvjJyxXA6D3XBhVuYfn9sM9
UKetn23hVae4KjojLjwqtKSFHrI4Y3rJmyJFRo5B/tamWFWJVy1xwMo7EFYKeSVxBdKOOT+w0Wta
4bPdXUMtuPazsUoopLhKuJPDfv8XqMlvwcSuq1hcP7r1emS+EXXH4vcPBH1p3VHGPVRY0y7ROzJN
dVMTf0L7mOTOPLxABVhz2aglijl03gz/kU5guBbn0ghmfusrLsKxC5My9dBjMUTwe60OHJTLEh6X
nMM+tNLG8xpQ1p2hj96ER/GCdqdNaDeyqGzKJgNj8tszD6yCpDB7qrB2wlldPtq4fqxLNhJBWr+t
5OgAae065E/tU6fGsDJ5fPAnBNxbfZVcTwyLzgRuau2Q2I3CdqNevs2KUam6D2J0qTvmpsV/7w57
hrns1J2KM6MVJC+sgYOxyfpgWSNlVowgnUUYYBzb1sxs6ajUNwQJHsELi9IeKWhs63F04RXEhT9d
p/s/SrkgLCNvMQxtbvk/UkDKhVEWRkaNssrQ5cFvUXLwykyo/G71bIer7ypKzo7OERj+bdggB+f8
lRoYo3TyqFu8ApO92RQJ/zz9BqfV4P16X601LEkcPihl9qLiYnhGU/UzCi5k8HBZ92vQ7IDo64Cz
mT0UQOc3bIojoU15rROViZEWlSp4nI69BpU+PrurhWQq28AktWs4i2lC+KuFlQAnC3bH8L8FlyMi
JhYJdhixs+Rp7UAuxHo+auAwyry0bmedHe/vdPGUrob3cpfDfaeA6dqOIAUKhqMGYmi2BWyuLa48
fWjsXI8fA6NmJLu2QRPpBt3V+MxulKegrLTqL/7bLBqYq0WYHGa6p2vbvwNjnLnelBgoXSDa90d8
hvaLQUTa4RLsPT+/bZJ2lkOu8RH0ukekvWRjET9AtNLh8isGCdKAolpuREVWpblTEGe9oi42U0IN
qcvFb90PGzzEyEjHNaaJ5Fn53uwntDId+L63JlZVSGoTynYkxyldX2wlpidZJX3EjXrGBV41HvPl
ervuI6iVY22H/r/AfD2/n3NewxLrNW94nfELfKnPLJ0CHQ17wSLIHsNRrFoMk4dsCkbZIOgs1pDX
GR8xws4daPP7kvID4AXHkxdk/To96dKr0HWa1J7Ku1g5a29EMTZzei8M6zD/hXMfmHb3Sur88dbv
lCDYY2VzMC49KvfP7iGi0sjIUg/P2j+yf7GbROzYOZETLpnkFqzdSnEaACe7iFH0ITPFCsR0gBQq
bgK9LoTsTNXN4TJ9j9TOKTz1OrPcIxZdD8XUeLidBi+8Zv4IZiI42Ftfocp6TYRwkxN92s02lXj5
gXqhubw2kkBsvlVbV6ScAJ0Lg4NDQ9p8PCbVwvEHXxeyjrUVrVETmhqTMq0QE7BLDiaYH3rzAUbF
mlPXRawjWrC5HTeaiCZMThHjfNJhuvdvEOOmezanTcFtogPaztUdAEyfdsaD3n9TQ26lDujGdrRN
LYRTo9vJ4a5dEbE7As31t4mkfcuW8TnYs7zpv9NSXpbH7Y5164H12dvnoLwJ+qfeirCEquOyMNSt
DjAMobHEV1Q7hZAdyFzCtm/lk2xkzZNR1GfxQZgHY3VgfTvViNqdiQUCobhCNmDE/xNy7ZNDJpCB
YYByO7JnPZNYT9tzgYhhtpPCRLtgpDRk77bNpUs4NdrbCaqPDJUL859Smm3y1UYbktTEUe80eTA6
WmvxZxgeO4GK+J2jArHDHBiTw/mz/GtuJOMMKFk0HY5S7bmD0FcNvFpJMJLOGUOmVFSuFWE0HHwA
IFOO7R8lTZx50/ZANGrV0AKvS96i28GOGDqVfRhMzaAiBuwlRo1j7EKXfzA/4ihfgYboBAqf4Rkf
EhJQP9B1He6dP9Y+oHekkQbUC5jHE43IHlL2CQRnQjk/vVxYyYR3VLT/wchZGA6pXGpB1iW3xBax
F9PwYAQsx/+//mfFkaxgX8zLSsny1nzPMXLPerymiZ/mvv2h+uTLuNQAyIFW43kXTZ/kv/N5ZVoh
WBICbCLDt1MQzdp0DpZjXwnRIP7bj6FL/rK49O+g+8OvD7nkKQ0yfVyDYlMF+i1p/h/K/LSaAEJK
a4MKvv/QFY1VlilX6so3o5VhFfUmY2WeYONNztgFsfyWzEB22iVf2nu3i0i8NS2Wfsk/oWdHdp7/
FMZRAilkd7HE4sS3uaW4+PmM3pQ9Sqnz6oTTX+la1grdDRV26j9WoIPQvK0ExH0pZPh4tOtwo9gh
sBb57Z/TBJGrTKAqWE5F1HfFOxKJRqLxnG+o66h6GVK5i1QeV4n5KSMCx827/QzfZoWunU7QDrDA
gUq0xU0Lf4gNEU3gh9Dg87UkVXxMYkU82AfUR/swmA7WwUja2i1edpqd/fJB8MaeoyhpZxr+ilvN
f6QEf877LADT0776LZwwE3f0RsQO5n49gAEaE2jHtgVYmdvxjZTQB/j5jL1JOhfdOtUcnLFhDz6A
vCfc9Pms2IHW0eHQytqxMuPtTnm6VIEJ7udw601a9BDJL/7EJIo2bddzlor/TShbU7rrMpgskmwV
fRmw7xo9KBW2fdrKF0laey+HmYG+8YBTcXCZP60qMEUcrVktcGY26D8NAp7YukX55KXVDK9s2ppB
o0k16ETTNBQ0Uxyq8s4z0XnNkE4XY/f9z/AmP7QXwCtnKnbE9PB9h6YkSRwKjazlXarNtlRHy94f
p1HxUDAzHLjOusfxKGAkWOgUBGkTj6CRDI3yvd9BkmQ+mSq87BZoJDRfhlDqLa6Krh3vDxwfwoAk
t4RSoXSxT7Ok0fsHp1mrC9DKaelF50Nsmr4y+Z5HGsLuKAB2DsTf6vKt76vR4xzft2zCWYEqJsJP
ltdoXg1Eo3DMr5SFF2ypNp0VqqS8uWfHuir7XfDvUT8FNf1N5FV+ba0FYucFoqgbUGZKmlTI72j8
BFZD8MyEzmpvKsUHWTEUigV7IKv6wTYcwiiPwnvFdajG4YCV0mtw7Tkf5ZslHkgxXYduPDJNLgCv
0ilctjwajXY2gFB7rqnHf4X3wqfPqX6BxBZd3K22ow5EdRajJx3IRvcdNSgXtTzNicH80cb/BXRv
2RQOQ+EbOfy7AjWpwctLS+sCjt/9Fnu7O4AFV+QrO2q3Fy1MVTrVaUmI41t1bQheMvGPxTYhTSgP
ciJzSsqdKEMf4Q69rZ51y6towgV76cRmqAKY/0hywFFgRpyxHSrmzw3RU+Czc/rumWvXSfMAaZWg
PO4tRG7Xnm7Qho0LzOzP6ctqDL71Qz/IyAfBeh6pTQrmhdKbJ/Deuy20ivZBHK51o1qZnmymFl6j
5ZHvI/TKEmuiWl8Mn1+Sevgqip9EEtNcJK4VDz7rJ1ihCoChjO1bfPSQaAiI4maqd+Gn8aDKgXd8
g8TIEqxUCc93fUOzmJxtiqybiaqVmRaj2zDctA6wbFK7kfZtDvgzGpfViSbFNCqjGLWBR5ANZhr4
XIhZ4jEPVFCgl8YzNcgI24bJZ2oPuO5HfOlBvjiJQWwsITXOWJQS50gnNNHy4zmX6nfAhGGmDsmt
z3ljdAflEng8r1UKEvyplu2at8siab0hCSsaQzQmYh52R41qcWM0TcxSP4LEyDgLx/47BfzcYhrp
h8vYUNjI45AtDS0vi5fLjwVGBsKq9zLe3HJL70hGqp8n8WgIuOA0+ei9iZO+PzXhfjgnwDoryGFg
ge5qk1+BpyNz59ZywMYWx83E0Wz/FwIbsuRzYysMd1+Z8+lWDHQ3+koji+lYaamZw8riRS0Bi2kg
EKd0b5QTMO3jdkuxjGLuxzOksZFONfPTazgbzI0BbLSDBCwfjfOfrEKMr7qrepQX2xBv/4xhdIBL
HFdyx1q31kqSyCMM0Ol/69Gi/0RWSToz5mmw147ej2nmuTdn8pui2mB3iyACBDpcg+Z85LuPgw+2
uxgy8/9uvKijWdtEK01GLx0B+LrxRGUM7pu2Sx1TEtw1jr0rO3D//rIDYzYlnH1Zu2z3VioIGiS2
7xdt/VrPW5Kg8624ZV0b9PwZ+CZIOWllU/2eGgNazjMYgs5YUEFOPRxfEGQFWv0hZ5+D1C3072z4
9oUeQikIsld6K3QGgHt5ie19ge8h/uaMVbHX2EJjT7aZO36jLDp4dIIEY1yM3fz/DFDkwlkg7S77
PmGBU3UfRHyTBhUBVDrIWwJgo9f79colo1Hqhemfl294QGZlxH5jr5ZjTzDSg7o5joSLEeXhgh73
5fhehUl41mz+aS+UjoZEU//qSxApBcAVgXiz8hecdANRcMxVnRZ/iljWM3ak1+Vn89kzWDrxIIkc
k/W86oemL5urCUMcP4Fw0AmeqV8aqr0drVzQzNC+yMpGij9YHUIYUPuOoma9Hb24GaBQrGlfNrKa
ntnIGHQVPvq/ctHLJwegW6VQzKlXTR6jzifNpiSATMm4jGy3INAD0pmRqegLEm4L88Dc3yX+vj+T
UObnKeKvDFbJvCdDTosKVtfbz+CwWtcWty2LuS79XXNme4Q9Xsb6NJmyKD5ZU70su4+Dx3WKSeyW
Dd0PsV8k3HlMOnUnVIl7qHOqk8tdjfbkZbp4kbf39z6NrGLJ8hCntxm8Egt66X0vQ1Ur1C3lnY/5
Lfz395x5Rdt2aae+FMV6xcOnT9KEx4nlXqENa8qXg0S54/EebRLI6OcCxeZO6d6uMUgz6FCblDKn
LgFaF+Gj5KMAxoTJmqgjfq4HdBF14evuMze0QR4VYgkqQk3MIjV9akKlpgm3VecG7YtBNqUVpfNa
m72tzdRvNns/n03egDLdqT5BFMAmbvc4CtboOw7+xcgBmlCibe8jUZePHlU4zR+9nQmOLvXpW8IW
4jem3AVbvCGeqZdsdR3KnSTcjsdGET3s3ykl4zVMLfH3WPhFOATB/wSbjnZCEU+yxjKKUCb9TidJ
f7g8g0AjxW5huuBxOhDysvtFwJ+p1CLluynCoXIBTmLgmki/DNO8yEXzScgnwwUhM2fGojIsv8wE
P/Nx7gj/r+8evwF6iqHz2XNURyAJyWozXSGMYALPBYHbClJyO2WMCUb/lKg+NEoJo1eJls4d+RZ+
61VAZfG/ZBkseKa96L7KyM9D80kogHCLwrWESK47dLD8uIeiYNFM33RO60S0ldF2wp91qJkZ4uCE
8cFGO/zC/HO6Ck8EEhd1MDfZDfSnqDUxdof+Xx5c8mmAhUxKOcGUgGSCJOpzY0Mz0gfEpZw93zcV
fmB4/a5NR7udpMYqDmHzXtQo6YAGgLcjRg0mdELa/32w4Jw4tLqhbnvt1QFwPWAZL7EoV1p4rgnV
67D1I94+WRlWEvb3GDRuFpXx1OO9YI7vGCKcC/Ef2vcSQp2gKYONEcrrDBfikNFfpBINUPve2g6v
qnkBzo7yk2c9n2ysFt6iuWDP43j6rdinhK6eElouGkO1lU3wnerHklUTlp3Lfm+wvbBjOrUpU+jY
I3BGb6xoEHI29bFZt/rumb2O8tOiBR/BhFBp7UblARNpSB+8+Ah6BU/m704A0FFHytKS7SWmG1OU
y9meykb2Bb7PsHIXqYv/CUh6P+w8hSulPq+Kn2RiVw9ceMowW9E4bfW9684npbSa8co9GVqx06fW
diiYXVA7LqjkHq6WlHCMHKv2W2xXUAjzZ4/Y3sCqssTusBeivq2HHM3CB3iHXmfAElWeNWLHS3yS
RK4hLPO6eQ9i3WHqSDCzi4I4RnXG1FOhRNqSy/E00IBBjYYuRNXrGDEwT8G/Teyt+OAn8LIqmUXk
Giqcw0E5i9KG+va9BarGH5EdYIkHkVxP8E5Solzck7fHp9QsTkoohr3d1z7AZchbSqPRt4XlasXM
rmKyD+bqRw9k/GZH7jI4GFvZJxF1NqdcwXWEMRfBBVBUxKAfbTYIoWGx0L/obFCRCZFZj83tcLwX
G1Toue0wedHDEnjXEKof9OVZVtsjV2X5SemAcVgjGj/25n9otU+I+1Qj9dEwH9ugj6BAqr60jyYr
w7e3TEJVMNBLvAEXn7b4I2bETQrH65i9XCZAmZ0kh/2L5yPiIyoZO6gnrmZ3wp+Po5lUu0WQcYZI
prPPSvKGRHoxSuf5lW1SiOdHYgMMjhDZCrF8YyRxWedOr8KeJArOJP5hXWrKTsj+OVqlZuJc5tWs
svQPnDaVuqy7fyixxJtVGaLrl+fcC8sCHbaMd3kQ12R28HtAjjPHicGDhwGj+S94zzyS8yowlvnu
CutBNSMf3eJ2iKhpsVboP/gxN71l62vkMVHFo9MquGBOFwbtbfxehB5KBPinvNAfnNddIowyTo4n
anm6JI0ojss9Dgw/BU0TCC2AnyaWriKeVV9B67eMsKgR/PXwRCroJ7i+8h+RL5QynBfTAU7TGdnh
5R6cqDtnYv3TDq/PqiunYXiZIoGpDJ4l8BA5Kr+VD0YGlt3f0ewRX7SbGDdqWDOsEe8gNrth6MFL
p8nsNszILhFKyt6hS+7J30YbrRQkjNZ74F4H1unBZimOquImsQdJQQ61ptIn2Kt4PexIzAhYyYWD
0ZPw2cR8hOV6WfFRfDU363Gll1f9BTvj/oVerJzgMAvav1GnQMUOm9s904ej2nanEWazN6RLKFr+
9ePvMryCAnowB5frtQhfwMsHiub+I5bt4QzSaLAnsHwJvvjkS1wTGklCqpxABEv3IVE6aMhY4mQI
eYR0LuBrSfE5t/iSErMzM4kOY2R2hruzbGD4VbsjxFcWIIhYoEB5lc9GEiYY3LolulHQ+eIk4ytI
oJOBeRUyM+kPvouSQnDCjtBvqjqJtafZ2908y/tmDcPAUS+gXqUKC9y08kt7ekiBBPlZfVxdnyrV
v3m+8axVhwgCo1bIsvF2SJhr+xRGcjiWQ/1UW9RIs/te+SlN1OMvKgUlmvSEHupmM9eVJfDPvSr0
n0CskJbZvkymeXmYnahh/nvbWo9BUeChk7axZAVsgQesrZnfX2peAl/MsMRGNyc6p16D092uOhJk
fOnT0LaZqnt/z/f8l9ogRCXSslMn323UOdFUI1VLWrXRAZLOszeTaoFAPDl9oyvwDIOx9sUWq/VE
1hvwAcMvuq4ZEPkBbdaVgwFlk1bwv+nnFyceWKGveFX9YlR7Zd7+wDg/RpxhEB4nuM4BVzuzMGOe
TH/Aa6E7Qx2Ud+EZibcZn8WawRM9dKE8wZwFpqFqC+AHWRMVE5xnWPMNcJd5wgIFak9nNVDJHYKF
fI5ixjFHx+l6BtrLOkBX1b06fdqtZMGgbGdH56A0Lazv3Eq6z4zUp4xB9R3vnD151f5KINnoEM3a
JSjt62wA7/SI2cdXiY3ZMX8urEVPkeNpdf+DnfImGJPTt2j0PC3hnG4OLIpFmozA6+bd618oNzrj
LmifDzpxmbLY2nX36qST27Mjr1BTT3pP9VCTIEj1ex1zccDKi/WcmpvmyrjQRjCsb7/0mwCawoy0
s/xBq8bjP1SLW/9T+tSDlXb5yFEhTI722cTFhA3NDhKcRgvZKkYXT2NTeN3T4v0C/cpX2FTQhE4a
rY+jFUEN6Bg4pb9w+OrcqaWfCI1GZi4fD/G1hBgzkAQ6CbZRw0OCcMuJmEHGxdP+//7M0VqOz9Pu
tXUGE3l/tCJ5LieShNet5ydbqWc1aB+GArnt81jAYe57sk5FetFS5g63WpVilTwlMeqtZSpgsEQK
PxXrGTGmD80y107wrEaLh433tllgqNZjLgLaSsOBOn/ICFX79I55RHi0vaf2X+wOiodYQ8sg05R9
NsQ80l/5LXXFA9HzGN8kT1UViVNzT+LPWBBFRehLsKbwuXNJF92n6vyBZFmNubBMAmjEE0T/m2KJ
VsC4CXQ3wPChx7eg63ekdHhukOIA8l5nqezr/a9oiC3tvg5syLdi4isIySLvj3nrv7aIqKsHy2xo
sJvUuzaWN0/BgbCEGbpc4p8QG+GYPPgcc3tbG3otQiOfK2fRs3k+L+o9wcvYGtxQGtiW/xpcL52H
dveQc+lhbjrFq5Qjvdte38PejcYMmjXTF+s3Oms+xOT74MpEy0sxbGFQdLGATthhR4sDug5ZYVm5
Uw4e2H2DfNE1q1weIEerur2aifXOrzc5vLhMZHDQD+yMItHlSy2deEGerP3i+m3NWUOQZLijlEtO
QyGMrvdbCEUSDZhRO5F87aiauiQW/gYerHqXz6ZkuJbAhYS5OMIz5lWed1XV6zX1Noz8gG4Yss57
95pxIEqrAyrkQ4FRwEreASG5I22UCrqBy6msO0DcCQpGBcdeYpu9j8pOy2CineEwtBShQO6zt+9M
8ueKuTCw2lcZObKlF6+e2xiNJDxgOkOtBuFPTiHLBFtLIayezFCeAwu82kbVFc21RKpPvs5REznY
ma4y4j6WcYa+1zlf1HUdAmrEJDxxsGszN3DxisBvMlJqVD4Sm9MyiN+Yrge7bYgo7VmxB6KxjUnf
OI3Pk2UO7NthaNNpfcXAzmZqQi+XhndBelHcOWHEym3y0c5FUs23KewAKSY8RujOOY/4cn3AUgMv
rHdOk1tm5ivPcw2eyi9O+1Xy6P+AwFcNVNADR5lKj9me2t1sSSsiYEy9jkHg9whbJUkoGiAN8xU5
ErD1qtJmjHmGCeDF1QOAfIk+Vr56bZKpT7dKLTVwxzrGLtsvQOyJ1nPAxSNFJUloXNNw2bPbsWOI
0L+JhPrVg1myD+AeyX8pjydGfi+fUd6QNyLQfTpdjC/SMmcVfyAXq9x71VvtY0d5x2DWhyE2/JvW
2bd9UOXp0Hoq2SqtmT4CqB0IDeT6A9QQhI+v8sn+x47sLmnbhoBfs/ieatH1JT9oyKHJy6oxsPws
WvH43UtYbaAcsPTqEAP/Acaha1ZMIk3HYYYLkcTatoryLjYbJotg4BOka0EiSg0Ql1eLcjfw7w7/
xJtrJKxlnugTMoangYWb5DPksGuSqXH4KGR9z6JFKG1CvPNnj2uuo5rleLXp6YT2kE1vAwY3QXu0
b4dLeExOJHclmgZ9JTGSZsQhjiz4+9KW1XIuXJymQfDXp0JPeeIuy1FdhYr7OzwJkE5C2D9QMCOQ
37nQGc2WPZU4SMjELsDN4P36EddJbmXZq711Mv7tMz+TGwdAeaposuqgfktoEkW47cGSGYopfhRr
1FXA9YkAHaZu/iHyMcfc4N7AT/RA1UFe4lKc0qVVmXElhtOWKCyo9B/g0FmwxjwPzVMFj/Zd88Xr
tY0CQY0aEEtgy1w8/b1y3z9dz9BslriGteDwEgJ3Zm7Ab/oFlyFE0S3BY3rhpanK+aY7PXtOCNB7
CO5fFqCpDLUfzvlzW47o34nxzcqMfoNMLi3yxoT6s060VNDMdlzBc5LMDAs+bXCp/98FMJokmInh
Y2nEXFHcht0AJkR52CVUmtYUj87As/HMB0rOdCiltdI1Fau19w9ig78GxMRTdzUb/YZTOR03X+RU
wrtpjOsqDKKTAK6+pS/Im3JLvg0zAAjkXBMYHlLEKpqnRuMg4pO8xUxb9LXGBYH0mGl9HTVCq8eZ
quQ6jydC1Ro5cnCrZfd3qUyo+zifTR3kQWqSjEwcH/Em6fkDTwmvNFxBVuNYZcVdnhzbPaZuwXrl
6mHMsnzKpBp490Z2+KMuwb3rpN+5oUg7vxYy6TaWsdF/emBk+hrHKRqLg9BTqgURXTkU2GwaBZ7X
4Ar3yUhVcJ7iMiIJohqfKtwTXdpOqRyvvDewxWH0hh1T1bW8M0WqJgK5mf+RtCQilgoTtuO7Evdh
gOscGgcW7YzOssCVww5lMk5kwRStYfuwOtZQomGj38ynq9myVc4s4/FPonq7HaJlrUyZ3lH/n6RP
DBODG1DsFiPljd0cyrXcouTntLMbAJbqzAqITSJb0QF9NtZSYHfED0dXysz3EFNHRj4xxeijzouw
ZSun/tYE4FwyRdGlzyhV82ClHtTC8xjybAZRGjWo5CcbnlI1e5Xy69tVDahIyBCPUKaTKzK/BCCN
o9HiF8dZXJW1lULVj7V7sigbUAuzQMMYO3rNESa5pA6RkoQ6dO8p9UOLORONfJPG+wQka7BA/WSD
Ik4RSAc6BuzXi/2YTqIzeGLtv+vSzxvpJFfEzt9hBSh6JMQrz8Yyxjfi/nM2dkmYuKJ51Jk3PqVl
zHPVFTHMGJY7FB1Sqajn2gvvdsmn5YCQCjIblTjnfffpFIcg6OkaJqfThKybCAnhSs/lFwnuHqSY
xrZwZTHzJ9o9mraNRSxC1QmpB25h98visKjizJJau+rZAyDB5ugh+UAbvjbHOcfIsD4xe+Iao1cP
AwghiD8C7rwNMFur640WF88Q0xsfV5HkWBuPVZFhhkU10nQYrtE157453Iti9lJHdHmz+N5koa77
iI+Fw67G5SY7jzSjfaLL5ZNkhxhgqfnGpteXX5tlOU7+C5HJ1K6ZxKPsrf/JI/vuHmbTiQuIwRzz
cn6ZL/CY9atfsH6iiBkaIKD+gm6XWFq4ACA5G54xvmPFU0QJJu7WUiKEb1cv3+3Q6UELt7aA4ZbD
cpVZt2gle6VamlsSO9Ter/zQ84He/iEVA8sNt2ttoGkGUutiySQLaN8JEvLPL+Zq6Z1wzjdoO59Q
+AkiDTfJkasqnbaV5iaIIP28cmAixDAEXVf7m1qnA3vI5x9rh3Aqrn5G5kZXCtqb6K4GdCmP6QOe
yLYcnaex0mpyOu9XN42fhMVaszk0FhNhw5aktyULLQ7MyYR3TC19D3ZnVcbYrxt8F0+soy6BkC8J
GboH5rHRoIDVRwnG1IGElx/4WtnDhB6cur2TY7muoWP5akowk5/XdsUc5MC3lbGEexQF4nB1CA3d
1UOWrUZ8XWsCYAKno3W4G/Y3wNSSi1wCCv5IpHgKG7WBRwq5IroezjmDvjkcTP0s2PkViWZ7I0Pq
g9w1sJsK6MRydEZSyLZETMu0zBB11VVc1sPo/ovQWS9hk3hEsHJpF6UmBIzlZhqahaenIpY6vuRM
WnPvlakLTxDdAgw7/561Y+4D5ak7Cmwyph8j/cGUPtYUB3Z5RMX+maBSBHNjRFtwlofU4KJ1Fw9r
NYthR4F9nApXD7fIIQ/88s43Re+JmzUJ82Tirn3mB2YCLz6V58ZRWTsjaCHeyRYL/+On35juwAdM
fg3NO2K5LUoLG7/UrdfY/O+r7eQG1E5rR+mA9D0zVqY5GNMLN5q7xkr4YaqUDDZFsvQ5jWD9bB6G
0dem9ZBDN/n/di+Bcb47zyl0NTo1M8/3PLMC54batclYlDI1lnkTdL2WyPOBlhJz4aechW3V5LJz
oqvYrNC+nYBBX/SkjsKmtvOw7kSEH/MxMMnsoGq3AtvdexJEcXIR00ZsEFtslFcLVlB1rfKglpGq
N7K1ShF/KrvMm49RCAWDbFqbMeIPFlLSRM/jVmuk9z2DrNDxmRmVMBq+OTJbeznJXo4eIJDqFyji
tVv+7Bj9T2o7zKcIzg0YSada39nuH2xae4MyFMBPaHpnOD9IspDyKAMpBShaxeMQzAeyVIQzpzIR
wsAMgA8Fs3RpGtibcxcP5xjLQp1//MheEISp743NOUCvXh4zihP//8YPAvgV3BHBd8gicGDW5aoK
0/f5NURZlpXy1OvOyoqZzkzs0K9f5VXORFJai+L1bv0OmtAnl2RYKFWv1xIuNGcNPJy0ES0tXtNk
VQoCPQ+++5nmhYHqema4Bu5Xvuck9pYxUAv2cHbNi8qC3KT8H+TpW2W3osE7Snp5uK36CKYxSMaa
Cx7gSFAR7r9xvt1Mvj+D8neQPJY9w+5VqOHmtUSYhXmva3R0wOvzTkGSQco+6zmh17CBT9wWQLHo
/4AiI4fQzNQQjc6+vkR93Fxy1im0mMwdI/4eVLw84i84ojv26s7D/kFehXTOU8A16rTje/BXKkgr
N4FSuw8xh0ESjksCcrbiWcGISD8rSDbB0zUl6HG/E6Z23SoTpXZdLQCssFt6ZyCsgdXUGjteWKwY
9UWNAGzwQWNhOkwS0wejxopEP4F0p10EKQ1T5Of9JxxXUXfc0lyYVDxfe+dryGOlBHgDIUu45xvP
ZilH6famxHstsUCgS237L50oBH9hmqHvp1icvFeUbcgbw4XT/ivrQjYsHd+P9IaGyueng/9oqf28
2oiub8mwir53jyY7DIgAgXjqywe5FtTPMLQeopfEfu3A33ZZT6WJ65M7G+smcqylh6hYlFEtCh1H
9pgVAgjT+oa/1v7sOkzvUi89y8jlgS2PELSjOCA3NsqkIxmuOOs0pxJORzMuLpVBtOoc6PnTn/Bv
uhGLOVXlMW8gknAMR9sbI7o9118W/wapnCEWbWqBaIH6MrkWxK4Jo2dkTGORhmL0r+8vuUefD26L
qBI7zwLn7nMFcu5+gfcqfX9bdSMof/2J6wNN8QNABnkDE0GY23GPqyiYysnMS5eJCK62MKy21xP/
swcgIpFxL5u8wdLconT1a90gO448NUAF3Ep1yULjkX41lXrQtbSLTmTWlh6Jwv6zg5rlq3k8zqHM
hCXT1zZgPp3IbOEfWZavocofAWoBBMC3m5GYBks0RBI9dTWbp6LWkl++sl6+9dLhK2zWZcJmhKA8
U4cArhfxagZzTqstmaYtGes/VCeG6l9gisJ7730jDWLiYpd50RHUi+4JD9PB82i3VlynZJ2L1w7J
l3xCxqKd+QDhNu+HwVOv/VIN3x1MkDgzZ6z9hZtjvWjIATiVtGSgZjOrM6AD7KuvI4e5+5LkaodD
yK8wMGTQ/TE2EhHseHTtl7uX9+8f5L3lkMrrf/9j+l3IwWEjcLqQhmwFjMYPXtBx7F0uHsNAia4m
TQlECeGfAaES8O+YOsvzo5D22IHi9QjhAPt4tBJUeri7/63scu12EwRaod3EenTiE8tfnrZaujyf
gI07l+jL0FPz/jvqxmObUc+Xfl957U4iLSjlOmNYquoF5y1tsQq9Lz9J20wgork3dFCzsCkVAW/t
kplCLgZiSEv8s3B+PXRdFIMbczQ/fNRRCGlToRNoEvNHE0SK7nscCsTGxYwaEHXaIHzmK3/2qc6f
XN1so5IscpXVMo+LkDjH6QFCFzw0VTs5qUKkc2bVGl0rTemQSbODvbIcYKP+ixDNnQDAGzMft7dx
Q8pDBfW2HUHgvCxYi35eM7dVdhMsIIIe4kSHXyGUG+Vs2uIu8gzSyE85pnoGtAUSbRmtNLuF5V4A
wqszIMsIkqq3KDH4qsXJ0MPqSLL3YiE7QbrX301HiYe6sPceEzW/6GOSQTU1atkYgIgUddPCtOiR
oooSn4OzAt5MdHK2IW/K5ertVOnrjDwFaIKa79z2DkxYy7WAkf+dGxn29cLZw1bfSXsNtYXDnPIW
DrTyJd0u8+BVLHbjKQfWhVX20ipadqNSqOiCxf8XrtM/2U/LjFFAQYKg3CvvhTyluCu7VQhBUJ/O
HD4cVsBLsuCo84CYlMSKDp4xCsnJttJe+f8QtkIhK5IcPeNW+gOfE8atDveqHOTpmb4M+hbxh0o0
zkFljMaB9yRE/ewOTO5uYvJ6gX+J8aZRBgnSL32nqELCFhAM9qN0rFjyqGHZkWuBxqL/0zBrDFf9
lA3NEJMM/CQIwbatcabQAclvXmnuWLAOSPQDCY2AkPpTUIC3HbLl//wniwlus5Cavd/YWhopHmze
6K6vC2TWEhJGP0GAfFzABt/e7dgVgmxfamhhcZ79Luv2UlfzufhlStQrpOwg4ggQLX8ap9WcQ2aR
Dn2pTGgxWfSaEzg9I3oI7kkRC40IBkjf8fuz6e6WWmBaFLO8xiVb7PoxBfs7fLxsyjolCekx6vLa
RXawMP7LF8p6KvFnI1WRNR9hzWtCRwjMmiIunusH3+jRe5rXREn+mAkLFpX50l1ZWb/Oxxoc0NYd
kmDcTABrpkRVqC4y2hCuSlp6ajBLF0aBFn0gsXD2dzC0F+t16notG+891ilPqwnuOLGILXhKCdtT
2NvTond1633cSDSsdNN/m652/NxhZWZHkKZbrVDQcetrzde4BjEdrb+7577VgWpSACY3mHXkNygF
Jrrh9oaLRw0Tymuw4uJQ4fDcmvmmZlTFYPCioUoXtXllLtBC8yWzAzGDwOg6FZ+8k8LS2HPgss7S
bZe00AUTPvH53f6O7R64RGGzM1r2JND0Oie7mZ+vMWWlJWPYQbuts06nZmG+th+YTIdbQmj9xaji
SlvIp9hNpr4WgA7bSvLzK5eO2KTFdRRp0KkJJx4wh8alFN61hQuY49ycBMjmiozICKihS4W5PSgI
tIsaP/QoWkSvMbkldoWQbeILqrpY+K2m5PzipMEAMd5kUgo6Y3C4z01rS+nzbnHO0iF6iF3W8QvY
4pkM2EXSebmN68w2uyhuf+22Kv0BZ4iNYER0gsYL+sMqaWw6I4csRRpdFlUUKbQNIVKOws4PvMjL
e/1RdG6pLOf74P4ZyEoVSjhBNyU5qs0HGoRVZ1T+g4YQsPGk4z+m/yM4K8+Km2Iljj8AP1iPFsl6
P24WOiSeUPcNMsWj5oawF0NnIWG9mJKFut6tBdP8PHmYQvWgDjrRs9imQohIj66qQe2bvUfdlWWr
s1pGjJet/Pggl7Hra0h8J+yZo1W5SmVM97TsHvc5Rf0SYAaI3/16L62cdvaO8ycXHmnGRUV8L4Er
aAns5z5XBznLnAb59kEOTyv0S575qn4QxpobkMIyXAZHXHFY85gThenL6h7CsBornk4U5JiJLpJ8
NDQXxlPmPRqzIDupZPg6BZcmreo8SYC0psbnRn1DDJG1D8rqxzSNQ9CD2e+Q2ikpKpPBOKLpeEPY
3jEsMAoszqJZILP2Jv6q8n++WRy1YSho0q6ZZzAwbJayCqhgBkhHociIAA0HX2QMESM1m7HzZ25c
6xmzJFz8IP/oCby3Wh7R9DX2W1zcdzZOoOCTkw14159A95xAz8HFrSvXvEYhPTgsVwMRlb0FUbwT
9+I68t5MxQY63tJT0M0ioeNGL7Y0zcZkoTJpY8lTyHgLDeopNRaF8+gqRSvmL8jn0inj/vRbSjjU
M3zyCphy0dA05IsaC3KBDLHoIyq8vdz914w4mHyvo1wY9ymzRvRw9XcBbOBPaM6XM68rt0+/vMqs
ueN75Oi9YgUEFZ2YJ65kPhFi0jY4WnDyoBPMoUD99BgApFmRIVBOOc/CNjHjsQ+xj7rHVbanVCK3
BWawP03T3oGmfEHFeb8AC+TxFcVgee3VwszMgZhkWL+2ciT85b6O01EKQ1M6Ck4azFvLYvid3jgp
eOMFuUPFaD+bnIBuqO/1fiuwDtEuUCimYfNlYEVU6+RPNdWm6+RDz5rOvCrQItEuIcJ2HvB3BlzX
2ZeVlYMGXbJQEBnPJjMy/UbNGEDJx1lpRGFupYmruV+GBi6jnHpPldWA23EW+A0cTo8LZRwQy9Q+
lUDqpzJGwZI0+jLrmcw5/DRUCda7Qc9CiFPdooSAVMAQpN3zt+m/lJ1/w3Sb86sTd2MnmUwO38J0
UWjCzQM7VMW5wvv/PtsL2CMOY8CaCmPBBDJGCOZf1YlVcQqNGEkpmrHLbIOuxuYk852bN6ZU4t/d
c+lAjTvTOqbVvg0dvTpMisE7Zb4XB0hEP8B9xlfyPXrJqxPk1m6+xlIg3tt0Xz5C/OIgIGWm9Bb9
2EDLMiiHQzZ1+CY/RTsXBT3bfOsAFJCFvsZ12vfKDAU6Zv2YjpXxhUe79NNk4KepfkfsHMVZudVA
7RseXU9W6pBUDnoXoLUA0LTKfT0NAnsfQLFSI1YCKSZkPOtZh4EzAjsCPcP3Jhh0V4yw4iKc0iIu
r38MTt4rEXjG6RBvVUtWYI1E86QT1sj5SF8YgR1iPcwhH+OEndYWxj2XD3A5We4y7tKnP6bNtlQN
DLD4PLONDcf8B8LRpoyn0RG0dDcz6Ilh9p8bLUBIlqU+VwuqXtNekozwAZSQZWYuSZFBBQ3sjMQ0
Nhn6lCzg68zLFqQkG5rCgg38u3R+UGvyuK8GQ2YRZ/2Bzcvsl9tdQWdGa6Igpz4AYhudkLROA/Ck
dfSQET/gaxx67mz2toXSQCrkm8dAx3COQXCFUeFpeMPINCaTF+4OJZsPlnh+LOfTA90rUQAKk20n
Na1flpAkJVW4GGScpAOxSXFK+A1ntyCqlfhpq/uVXyvivDrQZ9cXkjKB6DVDlIvI8gucBLNsLiOt
miUgx+Jka7HMfw9bor+A4z4smifELnwC9uHf+vVCaatgjO1sGkUHDWk5wehW0wbalO2yG8w6AK1x
nYdlplQ46+vP6NnCkMIEmp29uue0Cl6cb6/HCSdNAoM0tWTwO1fxMw33kINBGJiT444BJOALIZfA
OH2Wr/E86tLon3nh/XvOma8yOVXtONKGbyy6tB5NM0VUe6Mtnwr4ou50ReqpRpaECCw0hOe4iFT7
AQtlJPv8dmUfeSovkPgsB0hdEW5eqF+N1vWd5w45lPb26u8Jk/h/4iFyieoYG2N18QXq2X27MN2g
cqbO767goysJsf7Q8kXCbit3A9WrTXXJXmO00dPukWHGtH4iPskev1NZ9FbH7+YobAsUu4BECUh0
jwwQzSZ9cOedT1P4kjHhD2zRQ0He6bzYfR2oeTPcZzYYTUZFAjVfXiK6TXbjYVS6DB1rXlfCdvMQ
NX65wqEzvwKHqw91xD2E4PBynPJ4UVa0jAPTObinn5qIaOXatslHX6g30D8IeVszxfDZy9TvoEh8
L59pe6lQEMt/JQjVxeMx91CHD4AO9+ekZI+69gFMML6SnNI4myKR8qu9mY4FpiLvVHE1Nc7sURLc
lNpg91RivpYj7KAJ+DoI16k6FXRXYzDtbbc8pUBNS6EdN568N2QzfRMvX+VaJC0HOs9ixG+C0bGx
fKGVavHJ6WvYsF8qtMSnUATd2KKkdIEdNsRi1i/pFURAIP212MRgUlx/IRweFRaiSSGnaVcpSD2t
9CSYL05ZI5SlnAbCJjZTFlNYGCjhWCx+JbIC/7N4fEJdTRzXAeJfDdX4ZOj+DG2K4+yTUKYlJA+J
AHp6MfFJzRejFhK9eEzZ7nAGZi+rpgZeQquKDXBPhkjd5fL6spKsUe3zLU9LMncrvFzSBAvmLMUG
322qKKtkDeCdnz/3PsNtf0WKGXTPwZaLO/plc+YmJHXeqIuQInV3IU54RzO590/B5GzOEqUFiJ7O
W5gl4tw5eYnZZTJrEjvEjZhDL1lel741l7IazAEz3N/ic9Ff8u15tCOXs3EBEcbDYiyK+r+XTT5z
OUygGGtUU1NzfMOFRxw9xHFiJS82ihCR4fiSwag2C5nFOT42/Mm+3Wr8zynXVtr0Vj0iPaa+ofv9
P7YipqDoSjKFzcqbgvbPwGqvhUWa0cOe9tE7pJKdU61pALbUkJqkobaxk+1lWBJy5wtTH/BFKRUH
Q1e3kcTUTF0gTL86vZ15cfbYsB0MhjeltmZ8HoA6mBeEEbyyhk+6fbpgxotsmLG0UTya/mCq6pX1
eIydazU+dYhzJHGA+ny/OQTbdcrcfpCbglgsY8Ve9P6uHo/vOwDZao6byp0Xe7ToEJeWIOwZRuNy
0qhSABZJf+wQwLwIuA/7ppaGzWFu4RnEEm/gDLqut7FxNOAZU+0WtwfJe+ZQP25ko4ib20/RjJSl
4qtzAV2JTNvC3eIG3AdBEDvPwa8YSIxkkz7ich2JtkkaI83DthfMUNVNbSkogNLFsAigiL5b42Rn
A7KlNKny9sHzNTDWoCh98AzhzsQ/5x1494YD9a0+3q03zP9jMGL3DzqsZl5rZ6ycB5FfXfTimqCy
oRvkiLTFKDDWlbtvNJzrX9/8pRpLWFK0BGcpA3wA9hR5eFor+u4onLdEZL7ioGVLmiL0D9Q4rI1s
N20cPe3iyJ56sN8Goa/JDo5Eq1OiSzrZNaKF6sNxNOKf4HRla3X33cs90gAIDgjT5rLQydDBF6aj
T9BbNCAe4gz5xuCE6OhyMzMAqCjE060FuvP+UTdBX5gZI4H2Or7XnPw9hJrnrtwTrLpYkoJvyHPb
d49im9eGAAC2EJw2iGSTb3temtmoL4tss4k8jUstkmXUJZb533fyT0tF1I7BFPfvUNsDO+zsAw6d
fi8giiiDh55xIoC18WG71es2gtTynyhztOW1iXXB0/EqLytpyWNw/A+WYHP8Dr9+Zu6/QZe0Rxfj
t5LrOGiE7ZI4dqy0pUAjaBJuCV71+vCtf67EnpQz/4yeymhwfFTZiEWRf3p6P4VDj6aMo1PqMpCo
zXsNDR2LpW0xB6OgWBOssPktU7JcKHUbCAPXx5BcCfYt5Lmk1kfX4/dMqMJBAPx6PYsLRWSRR/ki
8Nq9tzOXsqgYQ/+I1XzMye1J4nusOI/GGyyCsyeci1k0c9ySdbDOj4SwOWsOq5s7fheHUxI1CgGz
Zi7ENBrXgoTv3AjV38gju5VSuMmkq4NO1c/wUM1NCHakAwVDi6hokIgYujq/iB6dGoNsUOoGCSe7
l5BOpjxVptvmuU8lJonuNR4ksiRemjKEsDh+rOlW88myZceRnGLIJSrfayTb1UqXTd4xxBiuJyCX
hrvzKF1zfewY9Z2eGVTiOSKZWpvw4dZCgbsI2OkdmYJ7EqHdPd/qDYAic7Y2CtBBJNX5W04gDqwr
qhuQQaH48pWi9q9KQt0nLRAnX2HhdRqZheYnOFHgtd5CwnFRcq0NH5zEXOVlUElkm2s+ZFHXOj70
D93mH+nxG1VZSythTB80yPUOiT1wR589mfeGFGWkuD9K6M7T/CBCpHKjG1IZREJaKa3qf9enLDUZ
Dl0RXipt5WexqDzhv9Z982BsZiFnYIcXorozTh052ivV6JTR2ec6gxAkCFwxwRZUq+5m4ny8AGsY
+9Z73qiMKSajB4EZWgVwnOg6EirQ5JZhxT5cVbS2krS8fBFj+fPHVIzDasJmlt85dKlGd2YBnIZO
yg3cP532jGo9vBYn1aKXlW40LMdrtXc4D6nsOfU8IkswyV8AddQVS08esWZSgGWGMnt/TgAeGf5l
xk4ldH6+AbfBXITtd1vr6mD2qEx0zws+mf532obUsZPE5X/PUPcImAK2DanShnoY1sijfJVEZkcL
KDOsdgjQaOMmiJtaXVD9CCH5D1rmqgz8dW34mA9ElbQML3jqQEb2jKQf0KQUDr+SB8cUYj2gk9sy
0fyUhP0MiISy8bQmNtRdwzu5Q2cA4PZZZHUQxYlMCNcXkUnOYgV86SzS/xZjpgFzl4wvPLM7g0iu
6ZnO2ZjE2EMEg8Cy6TFMnASu9jplboYYhiKu/BTIg077i5lmLmCZ0A2fyJQ0epoWLp/Mgt1UtJlD
ZYddpPCYZTAFOPHC+nffRVYCbTfKD5pFTuI0OMwjp8HGqETUaTK23Y6oloy3Ffx+hTBsLwB+Pz/U
kWSrOIYiW7Z27AikBAlBuXVSGXJ6HWs4O2LrLU5eXqL/Y3117mGiXrqBIg+EKjjBIk75RyoGiqRq
kJF4z9jeKeOtwdhNRxOS4WaKiy+HI+2q8uZANzc4ub9uWVIxrxQlNv6ZNy+Lwi6kEOtnfFgD5fZl
SKA0jVlQavWQ0Zv4AhCxbO1AuSAnd6CVFqaYlePRmXe12wjUf1Q1MODYA7o6xmza3lix2k558z22
AexrNJd3GcrVC8pb8B0Q4i3PrYLNX4MVrVZPjWwdocfk+OdaozXYVRUXJVTGSfRflM2LUYRFde9p
gOOd37MIA2PxcMPzaE3rdasXA8ViOfDla6rYyA4gxNdIMvnC9COJXUWUWGl5DIZd2FVBDovlzWFm
S5y8lMluiKva5wMykXAmX9wd60/0mdQEzGGm7+TkXwKvfW8OZ1nR+ZOSfg1dy8QfNQkjcwoZKnBv
Mwmc0GlTJ/imOU6oinAt+wZP5fidCPE+F+Uex395Ddje8E8cDIupLn9cf8YsICIAfYQ0g1L9SM1P
YNYY0mW6kYGL+8ltkC9ZUlUVeLvRyNuPMyzY1iIYB8h/Hr+X+OqAdBCt4+oC2lB6x9PbqEwXLDrp
OI1O00sBfZqUGmJBFv2MHj0dB67Kc1sbjPiYMGgl3JkYkF7/y7hE1VfVuuuImXKqVvmC7pz67e02
MSvo5sHRIW+/j3/wCKIdGGxazQEfrDbdF5pOODuR3K8Ad3hPinJb+PZJCrwng7/E3wg3i73czN0Z
Kt4mLxI2njoed9ItXeahUY5YJszt64wDOsNnkAbA4w09ogPr3/C9Mmgt3wWB42mmQiQmTaaz7jKK
6oBbBAlEv6SQr1xTJr/iZ1gugF+l0/wzxiVVi7n4UnnV/tGQA7WT6UAf6w/1pC9wcewrOyi+RuTc
ASuu7P6yGUOCAhAojU1SvKVOgLn887zGtpi4H/v7AUNlbkgDSD0jJtU7w1tye7lWh/NynRBXP6s5
jcUfGqTqwfp2deov4U9vM5AXlzkCvTBTl8QrMIsrv09pKKX58ALc+MEXkM1bJwG761qiNksYrsor
xBJqduMoehg61xCdxYlIpuwUK6PiIZKadpzVduzD9PKCSpfr7rwsSnwpe95Gm3BEGwSrJ3yuKL5L
P0r339dhl0dGv5sIbN3YH+3Ld+p4FiTaE9qvEN9zIGR4zxfmns6z1vaNPMe0+nsjqWgDDTQQix+u
fpVMpyd1/e6iaBEVN/qE4bddcEYQjtH3SwWAbJOVwOIZgn8HSB0b1ycSd1YCXS2BGYV9+27OtJpI
ce5+cJVNvhyyJ2fb3bNNctR8Hb+yIuPWyYI0h/AJLtnypE8gSitC7067f9rwTTlACj76OQn85h24
YS3EZ6egUsYJ0Dkpqe5GoaAmw3vtSUj1JK+s+9MRlx6F8G/OiNOOMvyMxp/zlI8R6llcuSUC6NEj
toVIjYOWQ7DjZXheLefFRb46yFJR2WVopeHKfrKIamRoTZTSBWclfZltacm2Z3/rKgal8qp+wTHp
7/Zgso/5MS6ZQVNv526SWVmKwIHdqp1Ef5BMQFpVeW4FsPbickR6KlyBdFlwKRdPgWQaBrvvOJlZ
RXvkeTYS3Xxqng19c3iWNJLeuLYUsFQhaRiZIA7ZtSyZGxDnQ5oBfATViwKgDeRFmUVTvdXzGLn5
65gqhRuWRlbHbdGzSEOsiBem6d56LdxJrz7hSiGQbmRlYe+j54z1Y/OyqIsn9G0wyDWArMJChzSA
+PpGmX9WQoip94/PTsDkiL7N2fB9zUezclNdDJRAm1iKGhDagoPDmOvITlasI+UeH+Qw8/6a/i6B
9cjjvwzBNR6D0G7UNdx/GI8G9/25UuyoAe8Wa+7D7GFjmVTVOvcDp3pnZZ9HSEec0DVQcouu3TL1
hpz8u93fgbYzl0Q3kQRJeUB0dF6JT2gLay6sJdqf95fdsDWk0LJFCi3RViB9PKxs2sAihQcZWE6O
x00fbqlDONngnO/ZyvYEN5LYxk2FcTR/7wPG7k/tmDYW1tb+lgX7APwFpiLV8emXPQvzC6PwICJM
eP7Hc+lgNCfL9NR3bXjBh4XiIYSnHr2dAVErCf3AB0ATrBPln/ZeCKXyg8G83s0K02i+o5mX3L/E
1FLbQI4/X2sRJJqxfuftG8T2pDmjEgRMuAdl5B0cqrYh7nzueoQcZtESGy8W+VI7ZewHe3GtpGEh
H/4QHhTCB4M96djc62YDTQKsnMBxg0AJJ3CgOWgmtwCR+lluQvPkROv2Gscj+Pge5AlhUR7mGDDR
AtiGDTrBlZIaMhJqwFaWRoQRNcwxZNvoOyjgBLUPdVeDX7FxolAOESblu4u2cG2pLzVJkruCiNB+
MJPgXvhHyBrxX9o3ITWOp+1fbnvtD1Y+te1Rz7oot25/qbWpsPIvoMbs8jD1NsedP64OyeAebQ8b
7VsL6MT5yK55dP0elcqMHA0b+0OSQNi87MeEgJt3djkSG8XLeGHsKgc35GOiQBvrXAjA/UHbUdPX
DTVi1bsZ3wUAJCibRJUVhtcjHMyyeCXoEY5FHH2Gdvb7VQwWkJSwwLePzFXdBjBJbuZW1gnFlcFi
ku+Vygx9PupJSRa7jzW4i0PScKkNpuBm3zBSCOzHINRvPCnNqfLnkHRpdYNv76gz55fooEbSOSM/
I3g6uVn549odIkifm3Kq0r6sAikGejgQ/MawtVHde7TpFi+jLHvd9Jf6fGBluYZYNF9KtP4Re2r3
CO4IaNEUdMpNJsBBJjIYLlq5RNWCs2aI6JqAcJa+06LzVcg8EEZZ+ylS6HIcNZJsaPFBMuGNG855
pEGI/PKbu0yRHNX2efTzN1Bg/KqyoGXk8yB7qUnyCY18jnEueIx9bMumDTlE8XRMXCEIQeOXVCB1
7o6rzWhFC/T23A2q8FBuHi6VjocCJ9Y1cNwWfWT7r4SrvMhfuyyDVaY0tngNJvtfAEDNAEGNLUu7
MtL6qb9z0kMM+3mvyh9va2n2+1SGwOs7hFvUSo6Q1ln5BAkit3R5wtgGWEBadC1G6Ox4/kOaci0j
WQCJgYEl/VnCqIUMA/l4Rvd2Ukyra+eE7jLLJQT4cfIoywjfj3qqjvBUgnuijUOoYQwJYsmxjrVa
YFSknQsxDzi07jGqsWJ0jXMG2Q6krJrmOkzp4t43jwT+LaWb3oujiK2PghJs8igGdRianznsOkOH
hWNNle3ZnvWi7+P5bVR2lx+loSn5kNR7dX0d0cJnRH7RTZKI1/WKX1Rz80phPxUq68rxwce7WCYv
c9Qt7l1QWtJAOJJdfcrB+6yR4TAb2VWo8nOz5WIvzVVDJ5iYQxe7lh/+54oN/fAOLaEla2HLBG08
0VtwhNRuq71nt5VyQbNobcc81IaQuOGAllu3mz8wZvM4CiWD2x1zvx5IbYTZjpyTyd7pSiI5oX42
hL1ld/s7iJl64e00DCgYDsCPuFJf4HOs7+RxgvBlDtpU5ST1o53sTXoNNzeT61Q/8Hr5Nsxh8S/U
V1rve4eR26D3zEeDRrjQTA6Hfn8WIYeso6QbPawyntBxC8Q71dI+yR3SbfC0Nh3jnWc6SgTms3YO
VUtzIaJynj3I5vQeYzThEA1cbn/NSyru/AWVIo1/HxFWbJ/szCCivHGrchFgBOmxuyWl4SWkzyU/
GrAC5U57eLYwfHfsbR6XHZr8V2VXUM1mtVpRku0XN7vIG24FE94ZlBFm7DWXAfjSmnjQUY0uPwkB
zNXj/vpUGn9Y9BZI2raKUObjEUBl9qu8h703H8fqIsQ9DXpiEu7SHCGgiHvk0OBXiZRELQMLIoG8
9PeWP+qLfd0JYKsJwMJAKSL9WCUCqV4r4CfWtbVc84YHoLAQZL88b2WPUcYree2Lnzjrhjzcx/Hd
A0kUDrGDco5wmUBmD88HQtbU8IM84tqRqu6JV5UQ5vM/KpPkXQBUaK/nH+997ofqg8TIVHECZh2V
FUeiTVEiO0DZ7jrK57SsMcKXcPPRe3L0LylxQU5vb2fAwEuOw9Z1IYiOslYFFr9j/ouN1rKTI6F+
xkpm26Ecta1MgM2jY2kty/5y/g6YKtfExknRMRqFEuTzhE/I3EG0WFzkTjM+vP76jSuTNkguCxVl
6LnuZKkw9Cn2s/7TLbqC0m2RYW+Ni1pJjqdk6azJ1RZQzTgIxyOl8XRJehLKlGz6rzDfy9xw5aMK
bpKmoj0XBhrs5AXBiLVs7gwNcDUY5katHPpUche9EEx71e2eQ8lbhjGSIlOKC0s0Mmp6cqMHsqgv
sbPENq4yzZJygnGeZjPEKgQC4+eEaXik8O4VZ6zusQzRwVlsf8Mmk5Bq8Hjvvw3W6fIoZD1cs3D4
nzyCOc4G1qwzV7V+OxBDaRrnX/93Ts5GWS+M+AWGmZcx/uEpGyJJEWvHx2sXtmy6lSOmzBCq6wK8
eJ5JPaiUpko6vMBY08hCMCkOQh2wAwuXc3YKNS56mlUfeZurhje7H7ktBGrf+OBENyHjq00NvlVh
5JR6DlVUq69kmuNl2EoR7HoTtHYR+j8XXU3vzGPgMtN0CYuS2WoHvq1FAU8CXoeh3TW6Eibmxf4d
NOTvCb2KovuAhi5Db6JBY1K/KXL2oZFpW2i2XXgglQiBnbv9FigVW4hW6qANf2yOvfgKu/6wOogh
qa5pm8pwXVkKS1qYpSVd6V6YiLa2khCY6hloNjrLHHzwr3orTWM7IXjgC5EpwysBYEZSuBH8ZowW
ImSY5aaDvoGgmHbNnsO2UewzmP3C9rMvRbO6wMuDOpdcgZWNwhueaAliF5MNnH7cU0xwii+de3iL
qAMlGEDvuVsp+xzZ64VvpVr+XLEAQ2oRN2+ISYKFm1myzKVqOQwwI3wct2qv5imH5wiGtLWm5Sbx
NbYksMRb9WgY+xHmyXRrdecPPles4kaT5IlA4jXQ/hSEIkZHfaF1gaIB5OLtUTZifpjUXeg6OYzD
4rOvMVBcZGClxdx0dUrE/mrF4QiBrFYykglHX9caan4ro2yRS0hgftjFgvsRZ9ahF0IyAdu188EH
duBcgAhWcesgIaAGrtfYqRYH8kB2YbgE3Jx4mjtni+R19NtuVwlIDyU6l4REWcPVDmTlmKrbvXcS
OUGdXhDGdsafOJbfrGQtsMYirKFyd8MMZfQ4XF2aXm64jsJTfGGdLTHlpiPOpRztr6bdppJ1IQQ0
rRseJNPhb7Ds5ygEWoOSNuhb12bBxmH8nk4xsdwS1uhKffBCVpDdhnTN6zX5a7QaRykUozwI3DlT
/gghOXWQ/EpA8629GtGCPkn7nyTPhzMvIKJzPpwSjrWEKZ6msJUFmXBkXmNCnjoZyFFtoT2DZmgT
MVSDvQfC6Kat6rLjXihfX7urE9COD86gP1ZE72kHyrwQULDrLlvLYcqUo1ngzFAp0IsQ9uKcCm2P
/yO4lNBy6p17rGz5WKM5KtD/KrvFGiG/XU6EkhJVFqXegLFEc72aDMFqsjXTBxRuCUeAih9yFbz3
z+h4dMudHo3BNYvhY5ycs0akBb0MHyKSkj7zbfI9SKEixH2fi1Sm+oCPTw3WLAIKK8556D2wchOb
iLF3x/Sk9LrxmggC3oXrsjXugs7SD372XVwOwAuDYRJ76kCM65fn/agOGALs4E+Pkb78+gwe0cXo
Ed2fafr1ChjLjoNkzBke61YmKFNeKpEwVC52de4Ku7qgASsMG8yuvUmO7KnswgNLub10O+VnINFx
VAIDVtmSNOYBaBsRqAfpOky66CH+jyTBIeEn5JJGWIRgkqUXp2WmFZbi69CztB1Irl4C6AA79mH4
Top9LcGLIxN4w7yRXvcOSB1NTV21XIFyNFFhlXvYgYfnVt4VVYkTrXXWRhbRCU6NzX9lbOSJOjUm
wGDWWw6OPcVJsX4dl1ojnASHLDpF5jSGLBIELt9ai/ZTBOnexhdSjXcGgWxg0VcTNPlhVLU1+WkA
rGRG0D60/2Np1rIfE+U43bpEdqRzOYYDNZYcQuoXjf4bJLGyLP9FGdC0h0K7Me7du5k6Th7z5+3T
YlnChcySMrr7vM67KisO8Uno8iygSuxygCGnHBTw7Lmfd6NQX40V5cjKF9HhtafWkTzjP7mlyjmQ
q07fat3I7V3nRw85h3vCHtWj96sZ12QMyXy9KFoCpSB9stwl80+f/i9zthq0frS3keMZ4f4k+YQB
8rx86n+DgpiUDQ/VvalJm4LxUvyflC0m/2npobMgvx5EcbzU+fDoXT+M7APlIfe/UIJJF9/mi7E3
c3+OLxaw9dXg1Nb14WqrtkuApTKWYR0QoESdO5Tcr3cvGJw9A+wiCqlXuGc2ksRsGgeukJxRWmSC
eGhei9O2GIYt6It5lJyOkHt2CFjaDx4iLHN+SwfwUiV0jdtiEeM7sh5NsgFYQm1WaZVGN0yyvL0O
tcFlsts9p66+N90yPI1Tscb2RqzXCSy5nEX7m7R0qakHJmv5JEQAWXOXEoKw+XvZjsCTGt0lwANn
jWqvPfYMa+K2UZRAkQCtftHeNpe0jV1DJW921IAXg3tG7Eq2YsSTpwyj2S+ufOjui7eNPVAWjHwV
CLuywV9f9L9JV0HI2DklD3l189tirvxIgT24K9FkEbeDFjN4lfboY/m1Xonn4XKkHiGieIUXuPXG
3EaskW0V1HOu1tHCaSF9A/hNndF6kFUnRJ2eD+MqLiEFqMcYRQkb20AUB+kRrCP24QKRN3mHaD8o
7IflP+8majfBXGoI1bSMvX0OljJalGPBj/q8KvGCUEyD/GzhrYdsqGLN9KRa3uRsYCMlaPYES9sP
lTujMNFipsgervQDpukh8bKLA2/nxjUDBb+fZqCvgl10ZL6jAKhOo9xQcMExcYezlvUjWd8maECc
A9r5cpbxt4YvNdx+sgqlu22AKT8JjyEGGsmcN0gJu4mFhVJxj63Gxf695EgweMPnlsx2ExEHM0Qq
SGsVtIVU1OFmByOTrxdziaT8ugSzyPcZ8daNj45MKImOX/GZOTNa4xxGx7Pg6NGeV6XehrqQHN8K
kYg+Ab9eR2I6EWZelIRJlfYK1ew9RNeTh8oJo25Tqvs+5Jt30PR6E2vnwVPhoM7PWR9PVcv7/GA/
Jq0ge5RGSDyIoYGrv4RqYBbwtsJoYYjQVLXu5/f0cX3UOKnw/Mi7cmWXSVtz1u8Xv8s/D3yBE+R3
XL0kWpI3eEpSrJGEIoF+OzkVadxqIBc+EQdiUg+ilILs7ov2ovwo7Vybn5KzjVePgviN2fJIT1j2
sQLjYwJrrT4evqF58Qbw8bptfXZAKl5SrJYXZx1MB3m2yuRrTd7+bJEYZmml3/9ZvrbozDyjzgaQ
dRMcTYys35kfVn8Dc22oXk9XEH6+Mcvb8nDltnd26eiv4OhoaW3WzrS2OAUAIVGNmlJcgmU8QIkn
9SsxTwkHF+fAgKU9653a7KqUJGe3PCbEYZaWH5ieGz1M6khO7y7O4yvhbNJO4zGiIjkW+fJxd7gl
upmvKseZt/ORvd1KQ2RF6mLrbj6F1FtbUU3DlsAI9gnWXBkZpHA81DrszHO25dKkVqoKL5bbiUnp
VkyeyPDdwZeueKNuvc74cor4pjyV3kP+5DO7TjnTCk81A8DidX0WbniBjB9xDO5LcmjOprMrsvIC
h01IXmJJIPHbunMwGt5lCirh4pa1FjIjV/CMvidtxg+YAc0hv+lDbyFJ92M20uks+Ax86PkU/UfA
MM5sWyIvy2994jadKkACWkCTLBMf5UNSeQPnJDDy9D0SOBujG3eOjjpufdCQ4eRszQXP3jfwzKk9
VtZnMLi3Xs474qDlIC2P7drhGkwBFycV6h/JmuoNvSAV3bQQ5P4HBsXnSeSRmBPZSjIztBk5QL07
ZmMbtOKiTgHWQCVX0Z+/rluRTgKJifqOnHknmg56KSZ1L3SqbcC0EcZ1+Oz7MdFcXbn1KoAW175L
Mya0jA6gvA+pUMUMYfYns+9nhDCrFoIpGLd+5AB2jkKf1P+o6a86xKSvipVgBXo4GK2dLxVd9+ay
8twCqLaGCycX8OzEMNnY1sf3QRlHMj7TqqGFX08xmhZzIVAti/4mauC3TMMcM/gIm5JwkxofSMny
5GeLyH0DOy2upiUVyT4MIwC9ngzK2SaLHoU0Wo6e0RXqs8mjmbSEWt7Lx/nayK2Bf7xlXcHiNXvQ
1BHxzeS+G7qJi/YqmCs8Km1UF9WkVB5msE+oy34GgQ6FOfivBE7KKWjuMPZ3Whws0F0mUnLNeSq4
V12/S8BSRBAfii2AOadlfwd+eLE4w14PtQxACcUaXdFwKinDWNo0rndHArEQb866N1orCeI1H0lo
2sci08Jr++9Z4K13FLh4nxfqDMSruzoHSO5sGKsWuljO4E7YfKI4pMKFwiTxub/JDt7xISx/ZiZ/
6lGS7oqGaJKOWrffxYZU6RqeidzfbzkaemTKyMSuJnblclWAx7md70OqUapjjOLegmPxGgPbjQhd
Awr3ntW5m/+ep7IHN5GxjJbZtm32mS/7VFzWcfG21inayEKTVAqzm7PXwLOrP2hRD24R0Gtuf5G4
24/J7xQzoKnq6i4UN6AeEKqB3O6BjbLHPnns+MWcbxSTjOxq44+TjlEbYemkrT9mqBScDZRrOU1g
MheTHzhmHmTrscHNFvZbZC4tqHfcIB6ZKQj5bMs9JplRBMXHCk79LBfl6k3DAqnaGotPnbS0mT30
RSoa7IdtBI92ndQn2g3/nBIcRdBaK7Za2o0StUz8gHXT3X5tPtpi58kycvKyJIyAas4J/PVmt5FA
C5ZTVyWkWbJdoABXQZH1Y6g3TR1q7+Lm7/cLV9kiLdUV1d6Ghxkyxhwoje4I2FjEscasEZHVBIeL
fDp+0ck8IIwlOaiUc/jsjgv2gwUOe1D5J0hsX0WsA49bQ21nmfcpvFC2C7/vesjLqfxfmTLqfegS
SqAG6MHTwsSIuIT5RplN1vc+EnS0FIRHWDDo/l4Ll1QNAxFWAQIuFuyHPzeVA/ldfUTv7Ii/MWnG
wOV3bO7P0Mi2X2MZByX17L6d7hqvcLU5QeBp23qeDFwXz4sWKNBUu1+vAP+HpDlsm/cGB730bG9H
v5bPsztKY37hc9cG/KqPG5CXwR/8vMhclU635PXEY/ggbOStKKUhiZJE69zql38A4KaAOWdabF9+
G+Izt6fx8ivUu2kTJLFKxF02Rfguv2Fyz0ZK2yMt34B2KuLouG85GR5JBX7h986UwCDGNW+IPC4p
spP3uU1ZciNByzgxqHjapuAhOydqh1NjYW8xy1k7mOoABIpXiRG5BOVue78T1+PmGrspqfA1x6G1
KEgV303NwR8Nohp5xLz/3EwvdWZhJcEZZ33KsJTm3ehj+3rf/4TTyk5wNhfitWaqCAbV1cE7VD78
pj5GpcOhmk9RzRUayjs3tSqtcRSbqYUD7mLnMmHyl3sHy8pGrtEMHqjz3m1ZjG06ZfwuouwQWPaP
dkpubiSRKhsixiTEpjyihClZ7xNhDvwo3sx6xomc1UfXCC9YsC9Eh92r4Qh/BrDrtZPC/l14l7ZD
4/pbZ6na60In0OOWTasRjJEKe5CL4pRL7fu1MFqbBp5NuZLCjjRke3OWCFPtD66rU8I6GHWz1CR4
4gb3ZTkbbrMNdr+Mdtab7tvkiNODRBwgfXtMNrKkuKduyf3mjMgTOQVMOpXnxPuOYv0VLfRL55FQ
oNH+5gXQqz5Y4GDKAloMyXz6kwpzcJPxq9X5olUdTlsHfTSLuOY1ayY5lJHZOa0FvYGwcZQ6KojR
seGtjbygHUjnjUMnEOj5eqY3rbmZMXamdyV2BUfK6SyE3Jgaw15W/yKKfFLXmTre07TraMtOgNvt
UrlCi+eVRQVLCuRrEOggb14HWJUsdP1MG5mNRCiXZT73Jjf56zr+IYQ50YLuSrlo1ctOxSD03sUR
k+rORbVyev8liSXPoX9fWzTHJm+8nutXJf1eXmucpLORo6R0NIW53ftQzqLajb+N6srY78yd7YpT
SL010aqT+i002GDL+8KhPiAxhGFrRpID4xmDPq9IGh60xJgIC9J2htYsqmVYrKmwAjETaSNzpn3I
ecUuVsR8C8sRG4K0lm8EYP6jnr5r6wypRUkBD5QoU765jJAjAXVyFG0Ej2jBhH5qugDTjWlRGb12
Fc8Z6vdScHM98WB8ufTH12Q5mrd0dueKpaUOkf4zofZCygb00tScYhXBRedTpCrz4liCiYJPNeWq
HrzthzlXCt1+24eaSd094Pelt0qVCNOHXy1PIY2O4nMTjIQh3nTMnVjfBrSxjs9DRaZRR6oRdm7I
u+S6YJM4n2bpLy1u45IEP0oWO1GduMg3PQ9x2Z8GrPDbURA51yX9t/Y8H9viixn7XF+N7Qk844lT
wn7RdHqLdmNCGuzIgqRThHrJ/z7KzNIcKKKLREQdHxiaja7Dhc3De7gh8epB5fPodwokV4yAgLVQ
wXXGyAJ7DeXPnHeklhP9X8BaE39I7wg/DF0p3H/7mIkIeDEiMMaDJkT/PcW6Q17W/adpp/51++vQ
SI5UfDpU3aLT/q5LyMo9ch2bXOyZg8p0Y5ihseQUIxb8/Siz1D1j3KrDy667f3PbgG+b9jW5hey+
Zs4ZDO2eE/Vw4RtbDz081BFaZvmJDzghL8s0MhKm62OFv1ET5oKuUFSIjqzuCfrsLM6xKXKMqmy7
rQu/IERuZSFgPjOT/TpC6QVoxyycBYE3aBQ8Yzu7FeBugNzt14qD9dCGgM8s19f91EQgVxo5uqcw
/qKsYYMA3X6/rJUrb5AMf5pyX4YCCr0ZK82Z1oZtGAvVLZN+/hrHW4mSjdQRsIqgxmlUz3TfbSnm
qWlJ18AEvLL17Lda+bVTA5YKp8mNks/7fZQWl34ttAuvuEe2UVIZCRiWTwarLwyvm2p2ln11pf/j
+LDQLNvIQAQfNvvp6pDsBqO/pgymQv0oZQ+V0BRwC890gKm+D9/a6MLojubH6T7ycUw1lhZChHoQ
KfIFS0A40RYsjYPt7aP5D4uP4UHCqWB2q5+p+IBbNQdaAk0HLmJKkctI4WhqfaXfkfDOjYdUT4DR
ZZ9Wwgs63DDT7AC4hT+tpE6Fh0dmx3hnRTayvxJeZQpKBQ4kKf0HVMcLFKl5MXP0HelX/JDS4FuS
og7Iir1hWj6dI2keKzydxWR9VeNCdCzEXcSDBZwrY78B/5n9EatNoXCs4LBH7Grw5wywDmJMhQEC
1px1c39B32TgTHTVHgiVE1l46PinBHsEkChdyzCUTcbC/MdsFg4GbjFZNhJ7CYpwdVZ9ffLEjuJF
QNH2GCvWsPZwkzb0yVsk/X/ITe/8QLr0tbgKFcPFAD04v3YBfCiPg0C6p2kiybVTgjCjdrGj4MkU
ch1iLzJtmxsFehfmZfOhwZ8lsCwG4rsEjRH1ru8CBhdLsI+ZmrH/KWpRDPxcKdOJDPhval62DxwQ
lVTRsTR2dVFVX2shUwF26oQ5OzZdjwwBYPA3cRrcuv1IGc6cCd8s2wAcsZJiGOoJI3eCvLUn4h+I
PNBdyaNSica5IjCFO3bnPWrZsuSjYLq9Fv87JR+Zo255ErsEmEmU/aHOMs3fxLGRcEMedBykP0Vv
AKinC+46sa7Y7GaKKVQYtj3/S8BLj7AqwMJIlqhyjRLTp6BWDBe0yTjbsYun1osH3Iw57TrDCrY3
kAI0rHG7aTSlHKO6TftMFOV2l7XFe9ojwtxeh0SkkAGrEKB/a1CzniTdv1+c1mpbPCZTlB4iP8GG
3cZVpPuaJBnuyD3sY5ikmECnVdIbO1DkCdUu0yWatuOZRbHc6egnxtegKO48hrwuzkQ+oREM5G7M
KiUAGvXKmm849CSfOFt2t55+gPNcvKljQtchErJLTjtZUiq+CoqrH4nQqVVTRPGqb30/J3GhQ+WR
0lqBzSd9SaG0XZeyAcT+rIWYujSv79GnWV/hm1NxTyXfnwvyQTOrC/Zd3aREof5JzKu2eFp3T5nQ
JQHLWbJnl13j0bTmRPgZr9HP0S99nZhQ23BByOamX0ZLsVbfnUl4VXLxmCECRkJdlDPY50vlLJO2
d6HAxGsR7+9qT1cnVfOKJDY1zEN5VpC3udEuFyGst/ml737pue2wQElwkxg6uNK6C379YKyf5l3g
bGc5j8FoJ4iPzcytxuNOG1ivkFJZ4YiKMLULd0Xzta5MnpNAwW0WnFHjzfAbRgX/Ou/ba3Evcgdd
rnDfJVqq+C8/509/R/f7cWm5JmVSfxtUM3DJm0EEcK+EI+6BiuuqqOTUNb2mUrFy/IpMJ54a4tkY
q/krZFnuWntTFXRSKWoYByYJ6YRzCCiDN2x4ZeN8c2AklwFfDOZfAF4zG2/xyaISuoBYyA9tVvXq
0dFI+hgEf0DpZmQsWKR6VWuEEErgu4kuyjK3Q+pq51jpNjYMis8EsKoRrEvk1pzpnlnH1VjX4FP9
X+/7vr0a6g0aH0EAhRS1IAm2BGBXAId6sGNaL6VMPHeZ+rEmYdAq5Qty8nY8yDqLMDgMQ3XmEnWt
S7xFzNbU76Xvpfi/Uywwzhli7RIX2VgV3SNuDEBNTgxwJZHY7awaHI4tdwCRSMKaXmAQeoxBex5b
ITUEy4HY683S5qE1RaYkfKFCUeyp2WQgBe8p9puLv2JNvpVfgsrjusoWPUlzuWWiE5MehYMYphMX
qevsnUPOFlOM/3unMR2nydPLpO0mLI6TCaBTZHrWcnXNfaqDNTCYpIalS6wu1Q8emaACRnoECoIF
Hw8vda+rNjjg2KZvkFHS6LLD7JpKnPx2wsDlH1EMxNfHMun88NRez6jIV8vVYhLKmnpGWLa7+leo
FF5yOu3HkPWsAw8qXQdPs8u5Gk81wCM58TCpw2bk8pGCfVWGMhFzG+8YcraUNPyJ129N6ns/ygx+
r9EW3gYDJjKCM1bE+3bOEbIJfDWJMqEj+jS6dibgjbYtGkUy+qwILfzubR8U2hj9zozhWoS/K92O
uQXB3dDEoUPdUugddPSX0EU906Gh9fD3ZCeC9cjTssFrwqH4gDiTQRkEjTWrqJk1tHPLGeyJZqXF
R0CIn59JkF4NkI9Mw5aWtuV0aNHBzHzTvYRks956IloBRi+0sfXBFnssdNiHGg0lBRArkXQztGu1
oQ5VXgVDi/eLkX0/k21g3lcA+4M1zkkz1wqJk1a50rUX1c3HdP5eOkzTx1zVfVSp457wmsh0hcYP
8ka0fwcl8aBkuiE6lKofLYDiMlERl4ZlrIXqM6a4OUpx3A2iQtYPg4WU9GFsE8/OuzJKzJcDFvjk
q+TFBLDllFdh6tc2iwNAkD3IXXDULEuHIET+TXt31ONkvC2ax3nY68mwkErOF23HowALPJ/3yQ0J
b/14v93mJw7xYfe52qOlw5Um20mFxrXI4fiMZ2FhL91NmyY4uAtp3W+TVjTU7V0axTYpXFKYyHP1
dWUfetUtyC0gRgxSCktgyCl2S4Rg+PyC1DGaK4J3H4fJD0/UVWuHySHhWJUDGiVVDwIoqCDUD8SZ
GgwqA5yMrQPm+//hjADRc2KPlXGgjzdMCFqmjMB6zf3LrTJmjHcCen1NIQjViqSoG+CVO5kwPoI9
GFibOE6vEWFFpvQsD2SiWzcnWb2Od4TZQG6HbovumREt5D28TKfNV0n1VPwv0lq5A+RX3NAK0eUS
y4LOpwn75wymTUpsazqlFpmgpm7i6Ot2VmrPFCvJG3a9b7QsYgQZypnam7L8XUbxitgUxrHFw4oC
rG1lKIMUZ1jdKbT2d/C7R3ADuqaJcd1uf1UObE+giDzMwVinEi1xsH9lClKTZCvY7WnnNktqL2fK
xJdQNTxcbewfAQ/Xpkpnzv9fojLqwfhjL/+ZRmGqHA995JpttCCRlDKVgw3OA9cwbS8qRhAusVmq
XBuZ+BhCOWfQDWsACNbMAm3b4qmGYsODtamvcXbZTW0lwur6PTzkQuL71IFrW+9K6DjJRs4hOMzT
uzgLFtnR7dAf0ExxwY2Q5kZxSnvM5A2zBadAtWbleWYuXoZ22Jb82Ob1y7O5HhGi7BCdC98SqWC4
B3bzgJN+mUzy0sM5CUuMqCNC8o+Cmf+nvXb3fBFvFzhb9VubCBtBb0J78O4yVOqqBWaW2/P+UiON
ExJenHH7IHuShUvGgdjKhYNF57CKF4c+ifG8FcaHdlxcvNzgDU6aD7er+I9uQjeU2msit/6mUxEe
zco5aiAY4JLxm7snYvEiiUKtXjV012G2R0R0a//BKqDcsjmcWh6KqjF9wXZ/CEs79WZ55tbw035g
hxmQJG4UN7fwC6e9ujmk88u27m+3FhEyV9xom92xG+4OcCwHQFpc3cEUxip3VjBYam1lzZpkm1b9
s1CaTbcXUfFp2y4y8hEnD+9AgYwJPekjusE5ajO17vDoJDsUiY2X5fBnVsMAN+SI8psjhuRDaTFc
I2j963NnrpYUwz2vpMlT+iQuWW9cK/LzQpvv9TVob4YUa0tfmwMUU2Rr0v+CeqwBB4YxEynoITrT
YTsP2eNYiZRYbks73PbW3B/PItFh0zAU6Uw3o1go75A3BQPtz9s4Xsubpf/A6J+r0yJmvq8Ihudf
iugRVGMQhZhHsx8OsA9w57VLxYw/4Zktt7DfJUqIQiZ5joE4W7UVk3Aga+MB5YfrQuQsUz8L9WoZ
ZkAjvxhMbRwDidI4zou2ZmwcCFacjJ+e3uBhMrTN04WdUzbKl0Uv+rUCP10OAV/V1Vs5P5UYdpq/
ZgRzcqr2/uNDDA7s0+N9qs3xqoGumAXDVVS0Vwz6s9ooZHcki2DBYFOwuj3qX7oGfgbTW7gwF0tj
3K+xc1yNHM88VNl73SQ46okVSiNP0fHMXFtCPfQKxzpq4HtVuAohBAHHNu6xUWPTSiZDuJ4hzcB7
I6ToH4d/xf5zGvDl2DcEw+LW3iEtFLvjxAAI69LRv0Pmq5maZYVH8Ayy2MabWWubOoO0ZM7L7v+d
qacl6p/3NFcdbVZ4JBNjgE87ZhIzWmPBzdp0u9DSMLo5Y7zBkKyOXnQO04QCr2QOAKLhr7no4GWz
sDLZcAn73N+X1oLAiFMVUtWrj2PGBk+KgcPPgkbmMQWy0zit9xN597FDELSFh6nuR2acLLCnQda+
MIuELgtGgr6lo4qHrBh3eIhakWn+sW5ISOQpEauPw88Sno9V1pQ4DpdIH8RjFJ5wroYIEnAW6gp0
P/YWs0eHRGGl1+AqThwsQxyX3RsNQh71fROZuB421Korz2we6SWYqZ5SE/2ywLcptw2J73fU+ed7
H62mfG+qZHDPAapvWYOUdaJsxuCYHUN2y0gpkg+Lc2kqXUbKM4Q62GtegDNsgYiyA8Md/Za3k8mW
KHrJfPHMxDOMvKhRHoxGo8i7aLIJLkJ+gKrTIwv+DqF+Rm02BJPiPAyWKhR3jhnvYg9Feki3jusy
UNu/92fvUmxbyHaWGXajiBpYpq7eVzsbqP3bxLteK52owBQ97Lp0oi7IymwYFC7LxfVgAzsmtP/b
1IrhCm1VIXhzgPV11sgJRiB6fipaPcnBFZm5Cqylyn1c0tnsWSI1nqvaHb/BgmbUzSTTcLcy7Yge
eOPrCIib6nAOla8D3spdv505bsxmQ/CZtQ2vRsbSzS9xYYJWq8qistS/mRTIqW0vBdcNnY/SOJsh
reiirojmklisilpa4t8B6jB8NV7R7zqa6im+3eY+XmC7PhUGo7F9sCOZCIxKKRuW2JaIvxF/3G9w
Rj4MrBqG4xHYto3su+e18iczzLCrDWCz5umx/idIvdhoPR3SOst+UGS2F79GlfK/9P8OEjiiEWvQ
1+LpomK19Ic6fgvuoYY+gLtL2P2wN2sBNN+h0PzW8p4iXRc6dIKbxhaOVcBqnHO/LZtCTlAh78fy
xkDYE7zCd1DB7Bsq4dt/ShOk4nutd7GhHehHPSZPNB6WBDTKWAbRJpeTjjplWyeguC/K86y47qBJ
475TgtCo5VhBrx91tCowjdLylYsbvubkga/mxpK7ctEzPHFGNSHq9F7NgoA5FliWX97/3O3ui0oa
tzngBCVz/fiqavbY5efSOa5uGcnlQ0TNzEwL1X8vDsvp8bLns+4o0dRhkcncBFqQwfoN5kxSngvf
yN/WcexhaqUbsunOTtrCQTzUysZFjAeukl2YbTrkYSt45MII/aZ+Z7Ikm3ghylbu4R0IbRuCFTxP
048z/eWw3CsiNsYjkesu/GUPmPzmLZbvG86h4DNbuTYusSYgG2BUhPcRZji+3hAvMjqW/ourLxeB
s58s5kgjRyjMDY09jnowmZXkfW6nlciNA+BCYJwWhal/UeFyEtrJXMOPq5ZTcMdnkeR+R5R4BA7g
OE7DgN74Z3cLMREiIsjgC4JKf9l8REmh9JoVs+K2I4TQYJNN2BaHd3exJO8fAD7Sfu3sHBCh0Iil
/7HrCTfG/UwXupaReuaxk6yUaKO6NZGKRpfGpuYS19zlpfS/WBqvKhSs+lSA3e8E7AG+6wQ7x2JX
qOvApU7DukEq8o9OETHrFyHdJ80UxQqO6L+k0NOTYHb44lcnWRDfDkUymvTuS+XyvevGAt1NRW7E
VhMQKTpkODytJSVhudPv2mrGviLSThoO+al/oR4IeO6PtwMhN1195bcUv0CRQGy9VzHYvOeRHT4x
4FrE9yMg+Wn/4v0QGo8gH2Rcxcj5Dpbc60g8ZUNB69/NQWt3Be6BKsOFYNAfyGdMoTweg4NJWEKl
2o4vOFoEpwjUpDjHfZHDyBsdjj7YZLfORojqlkr2pA5obki8+NtvL593tJsioPOR+JYXUActOPLF
n/j73F05yqvfIV6wD0LMYbD8o3dl4XYSFlt3/iVzYt8UVGuG/ahtHYKxDKXVnvunbSRO4+PULZWb
72uc6X94ksTSLohTUaiiANM4R1d6yP2NakM7xl+fdR3Pdh1sSAFinzO2qTx76EL1cVm4k9QGayhM
L6fwouA4+stS82MZy/uOI4YouuwVGJ4iQLFp0dnwb8SXC2jc05E/3FFMAO4+zg4Lg9deuKg4mk5p
dF8VuHf45TI7p84KvbQ7ugb+L3CNqkzw4CJrKy595/Myy8VXD16UWr6c9MLZvD63Rdj2UQHLmQmZ
DVEOvpKWQycR4hEsR30LKqk9z50Qb6RKXiWC5vfxsdZ2lVJUz3fLFUUMQTU5gMesAMnpKx6ZbHPk
qytLFm4SeFofrv8WXFWITChV3Llbyd1R9yVlaD4o2teRoaZMyMaUOMwKCX0Pys72hQPeK59fKj0e
3ITf/QKizNnlT6vWZYh6Ww/mpg9fjiwSev+wPA/wohAlb8wR8fk8CqoOJwwe9fVVd5+yc5XcVknk
77Oo8qYZ2OTTtkWWEkoNewk7gWt6KMK+kz/HR9mXDbbcS8igy1k9d0T09HGg8M+guEyxI+TBC9Ll
qrNUFk3tgK6zOOgdIGRvoUA+1FLKQhhEvMEDIANEw03jKz/VFqZYe55PPISg6pvgUwsDnEZLYnbp
Q0YNDTErb5zPhT3iGgxxNPveRYu1k77JYsNoWosCOknFfYfmIU+o66ixUXSc1Go+RWT8HQ/WXfoK
vZ1+QjWjg3uUbihqbabasqkbAnSmoucFw1R4YuCJYMsbsRWuPdfX5KmMARlA0v03maLjJmOY7Ey3
ydzMsbzyH5Ev3I1QKfuoirsyUlY6huCbzJhpbj82rQBnq3AI2g+Ylvdz9BRpshDX0Fp42KcVpn7w
4C+Yc2pLhfeMmGAag6cJ7hzeUBK4sfsuVAA7zePU2o6lNrXio9/1d4Ox48pNjYsn1cgMAcU7xwkP
jaUZBPp4fjuMQccjhvFUyUJ7sO/8q6q2Z4EKCGtS9wb3GDd6VfY4ycIWPArbjXVN3klhEndSDnqZ
ehU6oabzsoaVZ94tYq4HKJwv4U14+KgrElpJwfC+UzA9VBlgf22Z5YlMT/Ptz4q898669QYBMFSM
eREvCEhQ92kwY8sTV67o0paPDJRim5iXDjfA3t5+Ir87oZKigoUPkglzrGoS9umTZzayFqEcW36K
he876/WKv50nh+fiC5Nbm1qB2Uo0TG0+4fXEPKFpcHENoHItLcE8RzSeA/McuFG7ZCK0iQQPEznx
X6+9LfejwbumnnBcingZnClXAhdsgdCe211HKF1vf7ujNIlmSb79B8UkqHRe/h9s647YsO9wfl94
cfe0Byum0KIZ5vYt/ND8VGPBap7Wu5fW0+aHZaQn0Psnr+6XysK0qxUCxB+0f0bd2x3r5VWeESS4
U+ul+JkoId/lLVdgQ4dEBncoDfClToAMLBTG3UbViEOyNGamM2LSFl05lg0q+bBGGnAFc1+WYhqC
PVCIqQx/fE6pt6CO51h+hoUJ3yKC0O/oVuZQS9I8EQNGIeguPWoqeFeoQTica9+056p3qU5ZLWK6
LInC2KeY6fuWINX8+eKiwn9+23hkvolFaPsQU3lij6JvWJxZh7NcmOqTQelRv4YtfwQrKOkDTvH+
TVFby9iwYRYO5VEJCimhVjKJvt6c7JBAX/iZsbeX3FNdlVvt7RoaJyPRvTruxk0Bzl13uUWRdTlp
gKYGxEOp6LgF7dKG4pDQnC45FEixFJP0/pDqZW7OAguHIiaTzDDjdzAwtew1TR5ibF9+aipamSF3
+rdGTTIeWu9DTir+AgbexL/I2LlfHDRu0keSYevH7c2i3OWJNyhBnqAUQt+KuHKeUPnhZt7gdAgK
RENsnBUUtQ7uHPZYOQ8q5IqY0/vQvlVTYFiJw4gTdZONoKMXjywdQV9G6bQ0QlzHQ2GCJ8ccKlub
5m4AHmImMHKMfaTFKs5F/PcEjLTG3tPPRmqLeElsay+jbJNSs1R9EIraMAzlcqoYTBGjP8hI34VD
wB6mmsRb4XhAAmcBf1I2WJPEhQHj/CG/U1XhFD6oZMpXvErceiOw8iDiPODWyrmUi3OTMSRRr3xR
3hr04OqWJjXrzN4BQxvuaR7L6ZMSXC8+2HP6fepFUdGlX1fkpA+umb2kQ1p9E80Thhl7lFTtEkvU
5aLtZ4G1PruwH1oPeKyR6CyOBw0MHocvFp2umQgZqs5QeX9EB0dhL02wR6QdkwroLkT5G5cynQM4
BXlA44Wwr0C3KN0Beh+ClQEht/6Ip2w4r8Wu1qZc7spXNW2jEIR6nvK/sxnzlmMkENt3CzFupRca
z/MEFZA9cw6Zv2XdF3f+coaZkjrXNGp3fHhWeQHQG0ewKXOCSNdXIVSiA3dG/ZWUf7nocozpiOOo
A/ciLyWMOZ60J4pXUhwb3lIS2EmCpcbuYCOLa8odqjWmWmAcWFhFgDQ2Msacd4G/F6MYLYCMRya8
bUqPvPkuMpv63MSLQjoWb09+FQ/qu7z5ACATEvKIKvq0UU0kxv7S3Tp2vElnhCCeuEwADoKsHvUS
EGgt4QRWhQZhzjIVL9WCxB6fjaLeVQL/GNylWWeb8JJvIyVAX/asMall8CY0IdgUY3DI3L/lmpZW
OCejrmK2l+T5+zFDaWnD0EFN32Wa8/Gb0SbFmxR1Is2j1IxIxTgEK9OLfWBiK3v4YY2lfpCXpcb2
QhiRKLavqpadbz90wMWG9VXWlol4L5QvVNB5M7TCyhdoU6v439s3RsqcoCCdXBqyo7LDOYKQjJDX
hGdhXlUqWXu3RHYQA4Lu/dHWor6Dp53C/v69fUTzdVJGLhCQ9pJKVbw9YzIdJSIIdzYajT/abBdy
d00AWLsRc97C9q1wO0IRnQOgvex4DdnTGTLwEwGlwfSI+sLqenRgAilkCRgHohcvZHSDCv0UF9kN
wfCJxi5/aEmkmAQNtcWxYACtJ8hNBahx2mKpQzE4OqjXpwB3MtAVWoKfp8mjeirNaNFwQzscMb8q
QCEd3vhkTZit1cfTUkuhXiQu2xY+w5K6E99W4Zlc8ooJKTjwX+vsczyhvIwHwdCmDSHiAiuyp0rB
KJqchv0RDtrdiD3dcRzxOEZHxkzfklVQe7cV4CEeYezSoeSWbLnKu+RNZ/pjD4Vnjlm2vnpEQmTe
DjeZ9Um6tctHEcQhizfb+OO0TDTr1A9vXy4fNrOPjfXXzpsnFFsKztEGxRVaWcrzAeUWJvlZHPb+
5v6W56qlB1y+XXGFb2NEPGtvxitrrvwuP4qCp/QKlOgSze7xYYy/VU1bnZDKA2OuPpI8UEz6E4Xr
em/WhY3GaPyGlXpn6ILAysj849/ffMQ+pramKzxO0ym5Ut9/qkTQIdiG2fzFaX+Qag6zF9Dddp9w
XbemwFl4a5uhLuTHBVEeRoHqZxkFbUW9N4cnIAcRq9h+oTDK2r47gTTwEq9NQfx5yiDyYcnX9uvx
Z7MCxi+phhve4ZxMkAcJ4tighuKdO7WZ/FRnk9x1k/XmscOIC7tVLgaUQiR6WVHgiqO4mrI/1+G0
K5qUKnH24v/o4yvB+1vb/uzSzqO6c149M0RGj59yOno1txQ+Z0TEPrqHczPLwHrM/tVIrmw93WjG
iPvivfJ1QT5If8/3Np2JL1UiBWHp/dvL+yMfGe0/g4MqqZxm2x+H2Vo+SoO3sL/zco+oPf1Cpla7
qmc1IYa7LvMVJ/qhQW3vqaGPFiebCriXKs8aDvhLk+A6tYneoKQkLWYfGcyBKdei+Qmqga5wQdI5
GRnLZCvzkjNTUSppcTuibh/Rda6PRbY11oqY0Mv8ZZkkgiCAoTiqy2x6EPQrF6fzclX2CCzSbm/E
E/UTEdgynaZjfsGy3kUBO9OhtWF1lsrDVUkGIGc1klPL7XjQIsDdO9svLmlr1UT0a8I4wGXOaTmD
Vu2LI+aLQpkVpmGkkRlMsWD3Kw7Zd0LBSetISwjNnNY4ulXGHLIhBRcHBl1ipUK+xlIUi1tsyomt
4XH6OhUVe4e/QTmBJQM2vg7a8SmAonmaRV0J4hA/we0VF89iH4GgCrZRqJajQkb88QS07cg85wYg
eEhAXuH0b+6rtXss6H1aZKZFcncUttsdw1DQV+Rs/pJzL++QAeg7SLt9o4twAss7gMbRWj1GCJ/P
suBJteYJN9l3kMoYBAnaTh2GYpTtZzzTSIFnI4Si8gX7Vz/49dHEWd0wm3NegL4o9ZoTi1NpHL1e
EbhdXcnwBks/WLucywdVAjvnJO5FJMhIIPK3uVgStibI9oNPtB0ZUy5TQx7ly21p35NHvq39Afyd
/cJ0jndSIGc5ITTtvkfN9cTvdTOfGt3Vfm567+4JwRNGHg1Yt9B1Qg7XOSqPvQiJG6bwoaTl03tg
8EiZiLf+I0QdIT/tyDrIHYUiriZblZXhs2YajaKiYvtHJiQAQm8H+O+qFRE4B/IROAPHh42wTQmb
KlRBfmlww0RbV8/RVHFTlSN6+lyYzeI+a9N83lbqBA2Q3DvJBmtcLIRiXQsoPQFkUKcK/9L3qR6i
wq3+0hcp27+QK9bM/Tvnood10aExOnOiWqJ594WHurUo2L9MOq9qgaKsPYt/wmoq6oPxiPyi8QbZ
slgaKC1oIDoHRxclLY8PEqlTiD4ij+vDdW1xN1hyUUbQFC21aWmIQJInD11j7humYsyoHZQsOwMP
9p8CYykfoUnNhdWM9vHL4FF6t1xVq2YpVfc0LCmpZ3qfTFprRtVFukVnNCq44VPjw4ovQT1jPiHQ
FAYLqLSEnWHZ3SfE3LLILtOhho7bC/XL+0W4mZ9zS53U6fWokCOIpqzxTeKJAVveZ948WUjQUbHg
pgZG/wlNhKidDAR3l6RDi5G5nLNEPDIt2Edbkm1zmHgFY3YrvP9Gky2BK6bvuyG2ZMjVSuggzKz+
UgWtL76kai0Hh19FXHhdSRFpL9gliANTxmDg5zQgT270Ueb9OrYqdDppbzrWV8s12GLE2h8NCAU6
lVbYqL8ySTmhuwtJHMdq/hC/v4Obgawy74nmBj7lwJUa+/z932LZodHDJ23ASf3znyM5Q3f+5Jdu
yVoNTT5/3k01iMQkuHgEVHIySYfJpHmP9kbCjwcnDRNmFwEjMxoLF5YGCUN67NnYd6blqAWpPA9q
VCHzbItUTTWndNbKaT5r/lnCB5/6G3n4xvsDleIx37OwaKe9gouygeJYtBAlwa03dCej0iI7xQcL
dBdTPOUs7IwEMktHNuuIb4P8M44KSf1AlKYpIVl0CyA+sxIZzTpdM1b/7VFEOxXJ21cr/LksYluj
vIU567sBs0/uXYCrQme5vFvfPeV/7RJOtHfqXi1ijV3W7hWDJazy/MNZARbIwfPhXEFaXMiBHwYS
MSk7Xc/jC5tpljJwpUPTZFwl7Qv/0gISDPlHRScYTgzIj49I26k+zQTUjFyV3Po6qOzBEYFPanAq
I0Y30GX/eP5qU75bnuRNUC2yaQ3anaZLj/E6SaWfwOw51dszDbOK0zhcKg3QlHG3UMDItmgWF4u2
eOSleGNpV9//RAvEPMI2W35d1Gzq8bu+LRmNUurIlap/7W37f7i6Jqs8H6PyFUuqWLXPdwVyoHls
NUqQxKQyFZnFk554uE8S5q4Dz+aaIysjRTo2Od5YeZJ64uDZlXdb1L4bJ205m2NdHYDADGKqlLFt
N90TFNBbrLEcJxMZAs97RZus5+ts0VkDlqZdxzks5oSC79TZCPiwdnCXMpKWTOZ1sX6NzsiQhxkG
3DZK0Nml20ZSgGmi8mNFKNkpW6DxnQzMuf89nTqsfEqipypYFrphmwzypix3V3DVwhVik8LkpDBh
KNwiavEHRArXmPPp6oJBF7dfmwS24Y4MSzwm8o24v3FEZ11z2quj0usFxLyPomO3Y1hGlJSm5xU1
e6xnxtRt0zc8RKhhEaM1HkGtVdXR0otw9319ZOphMkcgk0FunQWJ8RmVr3woviKxYOHs/zY0+0Vw
pMKTL+hgi7g2K5c6RM7v4QuJUyIy+QmDXwtcEDpsOb673I1iLq8zR/8V7mj3Ljaxn38x9UFXxMxq
ImBndTMsbd11NrwX4uKhDFRcGX4J0u2lRkM5ZnzFh1oo/1qTEoElJmhn50CPGgy8xBlzLq15LhdV
RRKu3z/uiGkXeCS6UOgZDRV/mh/FgSqqNuxz743CvuT/KegRYoTZ2WGp58UHF/1tO2pFH6pswmwl
F4FT0BX+hbOc0+KcKAy1Miq2dFMsxv3QbJAEGxZEj46jtwr5jILhiWOmb6z3Pcq8GLWNDVSFFK5P
GlIsQt7UDWqwIPTVL0GZt9rVMUaOLxvk9HkQnynLjt5A41ahc21E0OajpLgpo0MIRnn3APVzNx1e
g2NonMdG+0I7XJPAQpSIv4eXn5UxAQ+TVM+gIzNIrrdWn2ug7qFeiRiZyq7F2fotSvx3yOW0ZRXX
HAhGUQFSoXjAmBBVYiPTWJsHcaemSw8nIexiQ1PXzwLAI/HXyn7X2EBNE+HsLJeXdOPss3LxHud1
31YZjv90SLwHc4aMDA+XIFvxTQ1A8gcUYn6NAk1ikTDCYyEQf4ajc1Tan2kBWfQICrTxSgRN6ZZu
KU/UGm6GXKUL2SM1Vc0CSEHbP4liJ/I/F1tQTBeu0sCuz3VfVB/+uF6gByCGt8Gys8ipk/XRpjO2
7sFumnNf2DkgN7jPbrl5Vjr1aFwyxQtHhAyxr1Jr6rRBnGVWtGpP4L4rca6hm3YvVZbM6inLLKCB
0m0QjEkdJytV8jEt0Va+LNRv+6UhjeLP/QymAmEIjHhevyPMAys6uiQhh5T0089INAgjyLJUj7OK
W562X0l9Avvx4YjVp2P/VMss8FhTclgdOTpCvW6QilZ0pYhUSINIF2aVCGVKewzW6RL5xjH/5eue
zqY0bubtwTu0mESKxa+Moqdb+3xhitPcNs//isdLsRAxsrN9CH+qSA6vh/pTwB8UtM19pIo2Rzmj
mmtqvsQSmsCbcbho41kehxBiwfnVklS4ccgYnNK8Jxv7eCyCu6FvHciYNEmWBQNgz8JI7nzjrfnD
2Ecbru5tyL+tWlh3ZpSApXNBcNs2dcp27b3AWVzFA3Ac+tqJvgU1ch3qVC5UXsJQAu5j9cCqXD1L
fxIHqoXV6KwEX8a0fady6D+VzAH2aR8ceV6y9m9CMOG9s7pNvFNppbJn5Ps8QRjESIlgYvnPzPmE
wjvHnb1/RyMatl5mSdOy2raGHtv727htmlMqMl5uozU6e/mTOQMUequt+aZ6K5IOztc1V8l5JoI7
AjgCN7DkyCJxQW3wovkuxe5JuqrDl9uXVftN+c/8PfgnlAf/SIHGGP2Onu3WQg0l8U7okgw5u1fN
KJ8tybqAvd4LahSkMMEJFbVipnQFE+gSlxIxvRdpRTK+Ccjz7w1BRljebJSZ4KOUhmTZbpiyszmv
jKj0STCPKaaZqV0aRKDV00dm2ShqHAGEAfHen2AW2YFcaW+S9uv+cbeEF8tIVNfbX23SFV9UFRGb
qNTtoyzE5AhncyGB0e+xWafyvJ5rpJCvTWvUdLFIotK8L3mdF9Vj3pt3W2bcMOsbmxggMReh9GI/
Ghy1DBsJUYxiVr7lma9Ehg4oscRKCZZkBScwh01IXuI1caXXQd1raa8qmX8eq6xQ5ndZGUjXOs/g
92EAGQaU9AHbiy9/LtUXXCyjHK20soTIZ4rGviCgaNa3IOx6MAHCh6MN3uQZ8FHBTf9hakFMs6hH
gNvBIFAGdU5Ec4LKOdM0pxv8QEP20fBSHREUjR5uqUU6qRQhZgzY3o639+2yYQzaoa3WNClQ8TIy
GGhNsdiaF43mA68g08BuZ3C6nATX2kiHJxTrAEYnp/mc/RpujITb1DR0i7sUGMTy/ug+u5j/IU5d
hZMp3EyVy4iyhrgA+FnLQdIBP3nhF0k5M38rduPzLNNWGjNXLCMk3tMUIAVTOd9OW8xQFRxBuisV
faFi5yqMt55i6wrZ8pvfQoJn7q7PzC2skK+j7VQvU5F7Us097hGo4GNlxN1A69jOLQ6v50YXlyHR
pdznfV+X174w97ATcqhno+VPoRPB+NlTa3Iat/5Wc48F73dNGQDE3MdKHw3+Hnss2Ghpx2qjXuNJ
f9KfKwb4NN6Aw82tLV7yroXABJtpuIwdvhsYrL8c31ox9Q50caffq9rWSPoKMBqjPJeku0hsQedg
sIKsnWIYAYU2+YljSXUJCJnJvzXLqkZ5C/iPDkcPOzVGCTcHFtDtGYmma6bURP11DuazgMy+blhe
a8wJRuvtQRAyIuxH0LInLtSMcVhT+XraHaLA270FMLOlZ94N1JmDp1zzLCI/b4+xyHDO+JPafwAf
MhJ49xqM0+w29m7A0gUgeZGJkZk+v6DedcON/ZgP6LeD8rXCr5PGbIN/h/pSA4d/UGyIh3D0BY1M
hjRr/nW0ZgV4EeNnnNFWz8VP4Z6zuFz9P/U8TlOJQpNrbGMAHqDvniJwzvTeg9l66GS7//kGxXud
XUt/ar4xogyP3TXVM7EkR8zJVA5z328+haqu3YSWBB/58+a8rdhMDo7z9calAk8ADa2slkTqHAyH
OaedJXOYH8UOPpMFq5i4ZQGVQ24+SuIRO9UgdOYWftspoxvVwfL7UVXJQiUGxMPbrc+KICM/rW+k
M4GD8DespcuFevcG17CDEqHslCm5pT17K2DUNtYCitB2ohDifKd+HQkT++3BKAehI8UR76U1n689
NtYAXdo7PbiMvXCq4Sg1qrF+fbUPyVnkbQ9gaGqDj1IztSnl/CQdcIF1PZxKpjKco5vmvhPQfEQt
gfhOxXR6X5SCLRqiIbnLSzRzP/fUbNJ40LJXdsx0cfbwmGRM40P5R7fwEBOTQtRVPXd/fY0K528a
ctbcHaWYAwYjp1S9StaUEao/027d81Oy61mSJEVV9E16p9sZkGbnL0tLBZydjA/02d235pD1DS/F
hlpzyzPRAjIrl7madz4QTQO2EZJiNMP9gRU3QgSpwRt/fjVYKbn8/ykf6yIZaVl0p/FEYkGzrxso
kN/h/mP7U7WKVQ85HFxipakwk+uXxZTs9xjk1LtmqKQGdnRP5Bu8E3FBNL78Fb6kkILcQS54JOTA
AJTf2OhdimmVsENuRCU16Haj1Z+pcLDRwVFefskoKWvmKPnMXWWB+CaxE6zdcoPacEYo+8DT2e4S
GkzmBZ9E5PAQsi3+LKrk0I5k9pkZvYZi4/XnAwHkaWyRMrsRBAT2niiYxSzc0qm4DlZEEWtOxuW9
+1hJPf0q91YmT43yVOTPbM2B822RHMp23XXxZvRJcUXYXxbijUmRG51ziFBkSyGBb+UvNbLrYK4m
1Q/F9CRh0+EiAVZaJRH9GI5q4PCH/TBbziaR0hrdnB9Sqy6A7PaTz3OXMshT3i0+KOgrbCue8bwe
sIMmGWOwZuFYYnTAko8xx6Z/vX3DGHcMwxsXFouc5dGp5EUcV10Gn5Jfv0e/LFbDLZJRnBP7efhq
u6y45B6d78XWB8KcxVae4YRY7fiPCyn9Y824RYJFqvJs2DW0TM4GzNm1z0sV7UPZogq51sF/B633
RTsF1Ar3UrBZjl2LO4mMQzPoXpXkxVVG1mPq/fx5HCYuCPXVrE4ZvrnfZRDKovprwKHltLxT6Jgh
dj1HHyzhJqBOLUiKAiEOIGnrsPMLdajAMs3NXO+XShSZ+nit2DVJfi57o0mSUoVMlNapYFg+qH9S
0udL8UoEMeqAPYoz31JsmOQ4jlQicLeWrSKR3JJrIRleqydFPgEbKqNSf2B0LHGASpn62NX4KV2y
KgCRW/z23ff39lwOy6Z7PuqhWH0R9lL5/Ftqz1e8fIM1FChLcB5A73/QjQ/cfj93Akc9T1dynX+w
2V2lJA0cUvbFN734syZr0RnnmvkCRjNcjK/mgjRLKkspBs51mDNLDuNCsZHAlZ7v8HEpwXO+yWo/
Nvsb7S+ZDCLRBZ5lisTAq/qKToXJeAwe6y0AXqGjXrLl/W4cDjei6lttRhYgiOPJbswPVCWEp0j8
zFvX4fT3DuO/k5I4gXlSs/h/imXwSCvT8Z4TBFDshxn6mFJCNU9v0PGwIf6BoWvpiNMiYsjSE37p
l8huJQKlwddk696ztPtpK4TZEIs5K8gKIIQUEgSgynV6pGvPBlFcCQBHuCbsAJpwHoAGc8GL2mrJ
jnkONzSyN1EBSv/M3iCOPUzMszHfTy7SpFwjlBeWcshKRt5j7EXbDir9bGTERjrVp8cu8I6t7/uP
lEWedhEY0qYyqabOMUQ7AblBOszAdyuX0u68VSI326GI8Sd5PWjGfr6p2hItYhPhAkzgP6viQiOJ
/D+Rr6n3/zpupoy+GvuwZlShZ9fuCaQovx5M3x9npzCRpVf2oij99Jqy0jVzZu/2FnS5FC2k6gtM
GnRlVrPRsHHEcyefkBdYqH6PLPYerW3Toq9EmI5v9nkn6/s6gmyJlwdNuLBmZOP/va4cZombVddd
P771X/i00dAAM0pXTOxp7g2g12wjPoX5KkSQqu8o6E4j5Jca2H1aiv5PeVxafuXg4WndVyEU1tE2
J0u7pk5ogRFjhtYCMt1QADrjN8wjW7NIM+O4M7XX8ZLGj3dqRhb8ckH/Ln80nFFp7mBT6V5iqzsS
sWr+/o5lw1I7+664LxK/dFizX7YvgoDqyWtm32w4ULl9xYk5xbtXN3RaPFjWyrRCb1Lguqpww1Pl
2l9n1gickhmxwsq8dVVzuuAJCWAzZC75wYva+9PRlBk/DLiWXHUjaILwJIGlu43wZB5/7uM+6hVB
E3fQi17NLbou4iknT+CW8WPhxBi+aNis8Yxo5cRmwq/ng4BoBb6M9f45mTlVvOhs95i2m2BdrxQR
5niaXyBZQT6jWzywk2iy6VgzMWg/Edev3piJu3xXXZO9P6tNPWaa8EENvJiPgNuBU9EvGWR5lxjO
BGRSqFJrDsiBwAoZZndIrR6xEtX6ULXiQXjh1XfVNEZaYxiSMbYy/LDgRC/8DLW24dhVXRT2OZF2
HgxBvNvPnyZEKc7SpPhubP6Jb2GvH5FQYq1n6Aue4y/7EpT28dUJHt3APU0FYgSgCRg/nGIB8pl3
1jB7kVuMBwCW+plPmK/iemfJrJiXZut3VQvmOi3GY4eSXXVMDY5GWjaU96ovFwXD3o2a5Cavh3Gl
HnHsGIZSdPTuKgQ2rF74x0uEp6jlmJwLBw2q0omiQRVS/oEWEcBwaMLE/35Sncv8gc1bdKe9Bx5p
M0JSllgVoKLaXZpwuB0VXmFB/5oNWb27RZb8duDPYqt3OcSPGLCPfiwihdal3ymbv7edWMrLCnJI
Kikhse8cidxH/62pMXx+mdAm/XdV9ED/vvcjU8QHAkeB8kJ6igDklCvwVx7e3aRwjRVYiNy/bkWk
9cTfsnDapZehscx4S3GI5/0+OdjlS39pu2gyDcB1MTVeL/1JdkktgSKnIxWUuMh8esHzeYYnvTep
pSWiS5FT9FmaaCwoJerLDi/KbzZIx1UFnkA431zrV2bgCCeXXwdEaxDrEe47SWbjGv4pr2ZnoTml
TbWupB0cbZZFNkqkydT3gbUA+or9xJGVcJRlhksyLW6NYw2xVop7EPakqYpUMky6x+x03jiFM0WJ
u0OiXC6EXk6DNaXaH9RvlGK6baNc/S4uKJdcMqYSMW7KW6TjbhTjy3O2SNuX2jy6NQPy6XiVDbzs
OFR7iLW0naI/Bbc5oiFAtkRT2xl6+fLaEUOgsDhKkQ9Yk8F6IL6PQubupxBFoBXxFo+EGjynquYS
ayuP6sNFgXUPej9RUknQkDKWfRrA3v/WTe0FaHKca3U2Xf9XCQY22m4geYzjTjHb0zzUFdCaXPdp
3lbqHP4xaetbHQo0NVFe4f94I0xLG8MRQ/IM4S7tR8RiKdvhd80H33GgJw61gaV7KONewBKP3Hyt
nsV/wQKxFb9n3jIlqsoGQ2zwQofforgiSSb6y5uZfrA7rfYBUW7/3egZpDvpirb92rjJkG9e3JnA
Zv/QYvc5+VZnlSWHZRE2t0ZssAfpQ/lCGDw16j6aNHFuZ8p4l6PeeFu9UmqGmGkgEMZsrTCk73FE
Yooi2nF2XLTHgsEu/stQgC89uI8cxQGT5RNkCyJ5ZIQpoLRMw5j/8Nbn/j05hu6cJBCOqrNsjG6s
kETlpTCD1aXU+iZvP5nV1MTD6oGDAX8KGRavlBa9wJoORJPaWQZGSTMWXvKn3klQRc42EB6IwiOk
tjbrDv8myH91AAHhMKTamRyKNimLAX/7s+54mOzu4kmnXGei0vzyuUVUSaEWcMuNFAY9I00R5o9T
oEfD25SY7eX5DQE1faTGO+tnwuRAfwoqhtu6o4u4geIUharSvinLSOS8epBu0xNzRUnEIDBoJ8rN
kN098sL0jd7/OBfp2dS4os7olyDP/AoPxnUdojsm5g0XWa9zT93VyJFitf0YCf41q52DFw6Kvm5r
6korVkbFCaHGhcPsqfZgz5QmgPD1491GBV4gciJ8uX4/Sq/GP6Bh4UbawZm2mjg2U9w870gzmLui
lBDKFl4AvBCxXGN/nQbgA3G3TYYW8xrRxfDWH/RdT9WvSJO7cXX0Gu6YSSPPwWwxdfK7cTpYwCT2
0nlNXQGOMUCnzZ4Yh5N3ujFGP0h086abGyBZETrgFFiyeboNuA58pq6/NB1NVU4DAUjABxPPFUoE
90TGgTrwJ0amw8ipNaLSFpubKumoAm9ipM3154AnG33PgX69baTss6CWp0Q81IL54HaQj2Bho6xo
d+u4Ne/aDitTwvMOg65obM6L4cYw38qwXpnzzHWDbGBF++QQsMlU8CKoWVBKUDDGVYq1Xj1vgFAe
4vKYZDbcfIZK0tjbyUj5/q4yiSNRswpwxoQl9lGflKjTXMn36LjIzsevZjxe5SNAPuLmzlhfKfab
j80cdJpzL9U41YOqlQyyEsB2PK67ls0u5O4NTJ7hc3Rdm0XiuS0b+zlBilyqUrStXX/WkmyQ0aJM
/4rd0nj6m8fm+4O8OWwsYDKGKf854EoFAPaBJUaCHT8kuNo8eqbdFe+tdoUQTHwOl6w8UdCuey6y
rr8b6Nl/exbFr0ULEJcnXpQ8z34M9PNqYXlymqCLatjjMnY52GV2eQk1ovrCJyiFj/Qbp0zswkTI
lXrGTmPZWZM9vMSO32xwbYHCwrJQQotGp0AF1gD96FkaG7LUskCyIC1yywrqn4rBVgIdTD2Mueen
cx2lMmoZsRQ7ItlBwaDlaIrLedor2vLq/gSxSP666iCgG8uJLcrIU28rbFAxAaMz/E7dGs0IHmxf
dRjitmylyocaqZSCe5aYd+RzovfsoMf1WFbY1TFF6rK4F7essjORhNStz4+jz3HOe3BXis/+/CB5
hQdHV1oT0Yk5izTiEcQspFGD7zTwvr0a2WyntmKl+WXFg3qK/BzCcbwaFCJRwIZvHWX3HFONiaxP
mRsDMx6PyUECnUJpHEIvPHjsJGglUlIVzijeKXHofnjMhUHLXkaQiPO6AJwctiX6f51CQOjbuOFl
c+N+VLFUcedZDDkxenbMcYvzozYifBzECEyWz/SkGd7XE2Z+32WNFwbONoHZxeju2hxcBxDMT3b6
eTSYdsiOyW/JpsrTqm9IiJJzRtR0QvKcoRJenaKPMb4pLgscR6Jjq+/kTD9n5K/FzyVY82ulggUZ
TmB7ESAs7HBecSSpuz7bgoOwrloN4qlA0xws34N9gVZVFDPJY2dq5qR0DT2J5a0N92dwGvMzZfgO
7H1JQb/TYE6ol4HIjVzncr/4DDlLiUUuwfogWCRLjMRhaGzZlpwSBjUyJSJUrtXjVeL+eJ+1TI/p
abkdITEDMr9QzKkthxAlm3iXim5gEpe9UfNbDLt71GbZPP6SYJgOIUI5EBnNAbeb2fPCDy4oP6/8
5xrSnhkuVQCDu6ajaABKqs1oS95MU0S0p/28O0OSlIdae160ii+ul+hpwNK0esbGoS/byAfwmM+H
CQxxLQK/xoxGVfi1EXET+8+FzTZy8Y7VTIdgMd0y0CxkbDncW3F8BxWppAbNjI10jkQ19Hb93jhd
eB4KjSVhL/4c4vm5irv1fiNIFNlaBibMPoc3jRlOFUan3eaF79G/eCUR0wXDzCxYBHEYRMYpD0rV
DDGwSDI3uLHrDNrBKUDML48FygpDVkV7vxG//cyVYLswTjMPjupiq/HDkSUnR10mz6EJ4zTreOkw
VvrGSptVBLjRHTqh0HxuWqplC2p5YcnR11vSbiPbGO3XRwu8G+g53mRWGqZ5jt1MFntee+Z91iRl
jWVA5Zb25ZMVeCpW/jT40xA1nmRLhNQVa3cYYREmeWwiXaH8jJmW/4wJFChIQ2U/NmryDaQTYSh4
VAsHwQcXfWxJ7qfiSdbZyE/ulNQZjQ2OI9xkIQSm8I9SBCxtp1U94U2aq9hjawZhSwahqVoCAafm
PxvuI0qNgIInB4jVyJeGWrUObk9fttTh/iu7FG2s+ll7tjDO7EjcleLu900pasYyBRYMtrer9Erz
UgeAejyiPxcdOhYdPVKEcJm8QbNsLItZVWQYYKWjqEbL80xvQjQCq1W8kxWo/WgiemfM9eeW7EMc
WtbNhU7el9j/fwXjWqtqlhoNPFJeiSEyhqgORgXgWwof5q49hgqGNjCx6bSod0MhL7kE3CtOyIJt
E1b30wKsNUoqGGYKp96S5AV50XtO4y3YKBgLswQOWJc20A+NbbERB3N1k784FTFuoAB/VWaTqlm8
kCvlxMG829TAZaZsOl6zm38K8aBCOdTfWOgRHb4KcWbbxR8kb6ISOYclA4bwtWCAMvMwjDOT3RKZ
+BEJx+AfOmvszqzIAGtMKdceoU1fNypiB6ZonWK/Zd/i5YjUmlOGOu0MJCQTgI028dbO5EcwAjDp
XvbgXdbXxMP9eUy71reF9miqdJrASN2FFEd8sNDAAXb/6SFX8VrwdH0JVB81KA4KnekolHAIttJH
uSK3f9yc06Gk0QeQ9H9YpP/HR+exLl8dOtJvVugirTfNK25juFCCjeTeeyNAmYwuvRfSS+rxIQY+
CDKu3vlw+DylC+7gVFEjYv71wSj1H8FiEqwJXsgCEvlBGsBlUBX7fy2mnCPQ3udRDgaBxaV6L1Zu
dbqt84lCw7sL7eReKEu51zxBJ1eG1GfuS1B44miLkcq4eTdOHSphqvvX0dGMXoDN6Bl360aNQf+j
t8qk8x32qlp1U2+2dl272yXcsh5Oc4i7Rv/v0yFB6OgcE2mEpnIeP8RAe9Jsk2ab9LK6jAVoTyxm
H7VwBfGTcYt8s1JuIfsX2hGvLuPjB/rVsfPCj/OVX5f/CgBGqoMy5w5jYgfBKKXefxZIUkG+gJAL
Xl2QcGfvShjGiY+3A6uM+yLCmecCLhKfSRologblYV+tTA3obJpSt3mV9yzcFOu5aeD5/fSlyZi9
ZwY440yeeeacYYgNRXVMAN44CcCrfjU0glUsxNV951OqRsVGhkFW/pq6LJfpq03MZn4b1bQNNXTS
hOXs37yM6Y0SUoDIaNjKamEpBkt5ZEVnZ7g8fZh1AL2CN+aI02stU6Zx5ldZgnzBoJHjPQkL/+t4
SyHhIeX58eSaFU3GhDKarNJRdzWYO5YPDjTbN0A2fCKTtXkrzcid2g8HOobtDKFlj2iN2MElMY5b
2sOvw7EgnojkzSV4hAn+EcYT0KuH2nmwJSxHNhNVTI9sHm91EsxHNHItiXrR7m3kcoro9Fxy7rt3
0+CqeGg61DdNpok8IKaYoi1kObJbxywZ+yrMhm48I/SuDNSvIey7MM+cGGxh4hZ2kHsl/dFW6/T5
6k7Rg4XzH+SPA4MjJccVXg4aUNeiwOc8k8cMhQwWRix4q4VATq+635ow4ufdFrWxKNUvq7uYWmuE
BwJasaOkBAF7E+vFiXSpe4427hNUQGP/oHZa1N4rUyrpt/rV5I3q2/ISxrkgRmq6qArvPy9y2jHk
xkWyyXJ3Mhw+vYx3cvIs23z1Cgdc9Y7RsCs1+TlkUa4Hu5SLJ62kd19tQfdNqaPBqP46+RXQd5IQ
tx+dRYFDxJb57IB7jmS6prpUOaFjOHVmv1bIX+26fbeab02ePAiCuLjOsrypmGaSGNDYpVxf28Rc
RMRdgy9Fd0maWhvA2jHapbljwnJKvonMfWIsns5hLd0E1SHydOOw/pTSHYqtzUB6VtoWWEJMMSyA
x6yBJymuFQYXrbqY0S3GzSDdI/OCikszylPu/vuVoWm5fRR3MddgE327TJfiHYK+ZrX6/lvAY72d
t7suW3bHAdtieKAl5mPiCQakkO/hjUDLTXF3uWDno3h3m3bjcs6RCbey7GqhGMtCxrQ7VHloxro7
xEE9BgSZAyTLmA+xcZHpKxnBBkXtRX5OkGOshB2n7htXJWS92mziydqlbMN+WkaPtxjdyf+CLaPt
Xsh9dWKexFgcH6cmTJKyTNoFyntu3WA8cU+KpWNowc//xwDzu/iPiHnmT7uSjPcjg/mVguuiz+/q
2wFkdeZ0XHYKGNp+l7+PkpO8WVptj2LQbO7WVDDEc25KhwRNXbViAszvH/vAteUMDYq/vPsHu1EF
s1nu0g6cvSsy8Wf/OsY2/ayQ2f46rPCVbsJCD77++cm6a9foHg67qqTDe4T9bhZZiL28BahMucpI
nZG6mRNIhhrxUzMSZ9QAkF/rtEq8mbuP74LkpoAnwJR5cSa6VeXGHQ46njANi2XZG4HtTJXomZ5j
7kKi8Og/uCWRaso1oae7pkaKwQavSQjD8JR0q+9RKWWTFPhdBSE+Nvt2tbGbvkHl1v1da6z48gKO
xVkny9mGunRSLPxvoDDwPGKFuw6ikYh7IQxzbfFzRJu9JSujPlJzIcSjjSaMhUlsakjnJwXBCNOI
uFvX+Prg7fmNNNkBQ+s7zjVlQ9Yq29mfbSK8osSmQ3swH/trDuMk7cQP9ifXztBwMUqAx04lI4nd
lfixlPSeTdvXnT/63Ag5OgF9UOPPejklg/rTchZ9kC01tH92GWK3AJm4ijTpJFtaheUMaExxtQ6y
L6pybgJE46n3kKTAwYv3ZuSpU591EYiIXHcFd4riQZdej1PbknYUtfymeInfwuMgg2K94eT+roBH
ivl0aLdGnDhRTkjYtPhK/PAO6ufnB360uHB43pw1o9Ty39a2hseZbgMihpF5y1KHU4RJHfhovUkt
M0rGepiZMC3BrUMxcE6y2cEXnU9UNd3FNgxqd4+B8OeUaNVC3S857Iq/rXH6Fy2DNs9hqEgPe8WC
PTr1BLo0cwrCvoV0OpLqTeGoucDWBhKvkZ2NU9qN0/KbVMqgF2zOsTNy9h5MiKx8dmSHbAmBweKX
4un0ybZkSgU2W2/V/gmwCDU10t8GcLGFpqLq61a9pyPa2N7YJwMBUPKSGzIY3vLk+5mhEWKBz209
f576wWDssOudWluPVZhqb1OAbKmD1rz+E9bMJjWV8kA3Fui7iiqF3lH95wpNo+1KPwaDwQF3+zon
jwcDRZLHJ4nWggUbHuxiwIugdhz4MxB3jHaKTCNO3h6lrY0cRkYl6pCETGJc3YjXsRUY6abeWFCQ
i9vIv2Vnh3ZVRjUl1kswXzlLkYunmGP5ZymK2i05HalehTGM13aGsbkhKsnkdBQvEDpdlkgNbxN9
L9VIiWX1fohzEcg4Ynib7Q9GvWRZ8Gm0AwCgMyeSq3UKUR76npv8p5x37IbJvxXuvD/lErD9mAwL
xB4JFArdNH+JHBB90y8h2J/Aekxvlt7qk7+SHznaLgb7l7Nzs90/fThQI2fPpuNay/rk+oQQIAqW
0Odwu9JJ5AcuYvMhZvXFy+roTanplycMnsOUOGQwEGM/EIQwLMjl26tKCFeOCbNMVPjVeMAxTZAf
1wLAcz9c8X3UrearOCeLrH+LISh8j/5cZJ0fH9e9wNcuWQSQNNiYqNKYRW3RlhSW4nKE48DRCDSd
4GH+el0CT/0nt6nJEty814gZ1esG5rdvSgj0ka15fwT9XN+5APP0ungklHB9suk7f/0WawNYH5Vb
gCLiFjawdYNI0iMQdvZfQcZ5gTmjR8yfspsha5wDziAxOUkL8iHgML3Bjn+Te7bcBy3RJTlRNWps
TrO19heQAAzB7kaB/PBXN/oEcFVRLZhPq/S+ipHHOrUcUgixgQz/7Ch97M3y8M+IhuF+lQuk772T
oFeSxiSGhG+RiBXOhcbE88XxNFo32va6DCYpUpb+HJFIkdokwmvAiHQ6uVX1PfvGDZ/l2TwyWwe2
rXdiU6H8KNBJ9fpwfHQZvsOWC0jRyvnWWZ+w7JrvyT0RNUMNi1nXOm8FWiJr9BNjv/REfmKL9W1z
wsadX6jtlYN9Bmsg9iETK4sOZOobVQkEgeUIAd/OdF1skkhvBq29u+rd1i47Lp8xLgpM3Ba3LrBb
OKfUjzwHVSaxCGUrm/eLD/NCvTq/wBNrrD0Yn3Cy/MFToQpTxHqi0i5OFhrcFRTSVFf1u/le74gz
gFQ3VOlFf4ePS1OxqMl2oDUc7vKNZb4vBv4s80lXcJJomNr+HXmQQdhdN0bNERB+Ap28GzhOkVDj
bE6qzCxzXX7W/wvawvXrQ3JqSaMkVCcK+HJ/5m3TkGOHMu6vSA1iqV9+AyP3irETtjscgQgQavaa
PUQ2YFieGYHOFdRsJOO3n5Z8eZRTzZXbpKwtViZto1Eet8QZMfIj99ZnbJQ4fxlafpXIPYUoqmIP
eaL2Y5embb6z4GVdOUa96nxhtWZzXvNvP+XqPqkrWvnKiW10/EXjgTc9i1c0VSuF5luorkyzQNL9
ri2TsL2Vf8RuWSpQVnL13ZTwnItZAn45CURREznH3GL+PBp0vxDpjdB1fFB0k0yIq6FHskWWDHRL
kQgRJBQ+cZdyp6Kc8QCYeXjl4EOaNNMfDbaOEPnjwNMja5cBRtPbb2jInI9c6V/XUI5vtIbOOT9J
Tp61xNE6kqU4U4v0+UFSEsGdUrvoxa1RKLhJhGuAnzOtPDQZVtvGydGoHOzSjgN0SZhUMtt7UlSV
2vrN3bl7qDkAfINErF2sakpb4cp3d/9i8p+s/99Nry8ztHzHUY1H8yri0XAE9u2AINHOaCbPkcjy
dcD2VdeF6NSve6DZfzoIQGSEkhj+296+xMzShXwCclB6eLz7M9DIrKbAfg86aB4kbeRSxhsZMuTs
83p2uCBsEjWtA0tOAVYssTERG4wWXeQLMnHl7Xo5uxKT6SXYlR25pe2ncnORjjeaRjU3I6i3ppjl
5NL3wD+Y39rKKLgWaEhgSrBNpniwJSeSvsxeD8AKGhAszyxQHPOAmefG/BsKLZXUy40SGaXJyp3B
96A3flw4c3gasWLRXQstInMGvHEm/wwamjT4KNed73H9eHcdtWMmEToh6FqmENbfg01OnHkPO365
ITEr/87b5GrUZxEWnSZPoCWSMaZgzFza0ckOOv91LhyN8WSni+sRLBGmQvmGfrBC16Lol+IpAx8+
Y77CIR+bCKofv0jtAp6W/S9oU9rzNxFGpaP3s2Kfli/PoVmumatAC5w/2wANBCPu6p+wvJ1/JwQq
F+R900OXErJ1BH1vG1M6mFgj26qJ+AmI8Z1kmQ/wGYsoTf/Y4bH0x8DLPjqhzJxJP2e7gxVvnVow
Fb4TYTCR02dYLo2S+/j3Rc1461gC2qSUUgL6fOT9iZjpPikqeNfySZ2Zw2BVEvm2EhyJZmlhB/lQ
2La+Qxa6cnxx5GI3mda/7gKJAuzdsHl5YNAEVY0zyp95aKKmm8CcVP6G+wtW0rKXNZxiNgLUoA0B
y11SJSHWlygnuPfqpSHgCVR9cQfbrbJbEM2737EDxzKZ5/Wtx4+YcRQimCD2NuqbFCZDSRUi6tkn
l9coGINRntgrY0tmv+k5p9m4b6Yujmyvte9FaMZoFWsqtt2Q9prmRtIWX6671KD0bO1NNinMX4jO
WaQ4fixrOkUjtmIraxVqUTY1cR58d6r4ap7su6dKxV92uPXTQ0WJ12AlH0ARWRT2VmOzAgGb0gf9
anoW7t5WJmpH7rkVqNl3yzz+f3VJK1//qvVNlUcYpWf2MZcVCBQohnjIKzoptXbFTY5TjfmbOhsl
n4oJyDjmzTCkr8XWuGDnwYv2Vll3GZPCMMZAt5PR31GpRRYbAKxy3Tk5mpfeSmnCa6mu3p5RlqNC
5HiFTd84y5kwBEkaNSA8db2GbDp9z5LLazCOAytGssxm4HzVA6mHO2uEV44UeBape2RYp/9xWs/q
b6uvQKXHPY9DUCewXXQtwArVtDKAueXIgWML3rTTY0lX/JqyOwBuBK/cSBxWmGcYlTeWirjW08Ld
9mK76dDBfX7CcGiYyvpCtaEqG7V4sFYv23FDP2q8qCH95JCrz3MU3718BI14rZKkFP9C9aotgokc
xiH5PxG0IG9ntqSgRBWXrQd/BYjC1mJsTccwhcZvLX9TuuFVdx4icBZHSWxmnk9XKkk65OvFJ9Er
e6XKXYeLToDMf25QzQkmTvjlrN46S6wIgYjYkE+/ywD8xuwCsJdeecJSJvRDMPXMavkA8FsWFCP0
/UXmIox7vJ7C2KoOE77e9Sc/tz/vQI5/0JS8N194yEZ0bxtrYWLrKgSfh/F82I8pfkzHDNs5HsNI
Cul3wQ6fLQMd107BTQUC0nlNnOJh2hUVbSRCNSg8lUZaRIuOYS4cl4BTwpujKAw0Sg50YGCyzQxR
5U9O9oqXJrzWU9umkMOuke2I8YqICaL4FRdasiwUJrVFLelruA4D7Kx4Fa4C9c4qIAjxWtfjIGWO
ZCKbvzzrsy5Qx9njtxo/ceEYfJukWmCmUuuPlauQG9j61gZvScDPrG0vOmakYRFaaln0yptGTV91
Z+7f+lxU/KxtzUjBHcEYhM25zcWt+r6Rs/WefCjaHiAU2UsJzchtkj6ImWLalkM150YdSu1+B0TO
EwO56Y8oxkA7sKz4J7BpEX4MKmg8YkKCF3hAvpv0stq8Bg5Oseq3l4+FyCabQo6pNtopRW5ZlJxO
FCQrWtLlsk5lZO2KOrM+flJrAA6paM71WWwdoq6IlhbENFD9kQoJMU0lTQv3lk5iLhTBv04V+Qnm
e3uO9gp8qDqA+RZhW2oH+kkzXUVmPqrWPQo0uF4EBE3ZNLD2NL+SXtapLdRNAWuCVxmnX27eT9qw
g5FsKIf5aDLK9B5kUHV7ZndR9tYN90U55BM5ulns29Up+F1oQ+7mstzAq5aseJSq3fvCgfdHUjce
Jg6EODo9P5qSOb0ROTrOzznnE4xRPhUtxpPHy5DnDzNRCr39gFoI710ZsGf6bFenMN6HkqE9T/AZ
imn7jLaZnZxivGvvnkWsDuuZ82u2cmxvj65nWuACc7xMF734SL6I2n4uuNzrNNFeK2RabHn17Gvy
HrhIVSTngC7jTydNFXciMNkZv1wqbfZMdCl7DXs/JGaE/bdZm4w1hWf+NM8qZzwuDkBn1srVtDU8
Hf8/n2+ip57ni+38cg2YeZP+QokuJ5q9UVDV7W4qNm6fcJnllxI3D0cEuQ+H3gDucGS9Qji2zkm1
jxdUTW7Bq92Fq2xG3gR7vZMYyz39973AcScycepidoEyRxT0YI0MmwFtMZDhzzkadmvg0dnVFOWs
XbioQh1v7CVPDH0CRuOdUChSaD74xttCrR4bm7bKvQCtIrN5ryyojm7MTXg1CIvFzQkrZxYi6DIl
/bq+/wL3cf3RQ3kIJccyATYcVGYC8k7kS6EdFQ15zpcn1FJ8M5sKqUaFdbokcFYRFzWsjB6yYXor
iGxgUZCsD9y/prXXV33GyyKs5EJuifZI+8DbkNPCAM5V2w7JFlgoamPK//QMnIY4osys+tnMll2Z
VZzl+7+JU2ooDZG4ILiVmExqQFZVnCrpad49thmXdDNn9hix5WENWQTUxrGt93OH1m6BFDFZLRpO
Hqe4/voJpESgbhugs0iyg0uJgS1UDxLCh++LkdmdDU/ClRsDtVlUBy1TGo92TP/lOGwJ2A8CkNdf
z0lGgLaGza+2yoLL1trTeQ19pfgWDXeoFqssOEJOzUKlXOf5vShL7a+JFtDkx8G4B5/f+P7X1NM8
YRCP01BSH/0MJCG0Mi1lHw+i2VbvEcQtWSrtITJ/6sGTk2qWfU0BX6Cvp0NYaJLjV1c4ieFNwcvM
y8ed/spYYyTuBc8AwOlkrj1G/7KFP/+JSnJ5D8kZHPXVo2Sw3Y7ubceCvMpA3gzdkzgP1Gm29+Te
bLw1B7abTkzI1UBAt2lUNAxvOi/wI2b2qDCPWc3vDTZR/+vUfXqye1hzamhLNYbfnmQQWqPdgeDC
v4lOIDblUICxyiYCeWeRhONtogUQXI5EMMraK2rr5aOP+AiDORSDYKkxieZBKL2pW90CfAUALLzb
NcQy1wzN9VdG/KWVD22shmiN2UrEJX/kFo0qBzOSAVam57yiwWEX+wZQABOzNX5wqdrbr6d6Sf+1
uW7bsmZ9g7XJAxMzp66ZBy/x1pgZHexOxx90/r9QngmtTpQ6qQ9k+NnTqGkb+GYwxWsqn+/0mab7
6frN6HSwA0s0hp10YpjBHRlV9aAc/kI5axzR3Sj6wTmUh8xCVhWrnn0f9dFR08rm7+uMSdQjL/aO
xfp3+6LFedqRzclpfvZ1DwwuQTC5krEno7oqkCGoiWG6RksGPrfT3wq8JLAM/9R0XEEPx/r/Fo9T
SDt8NkBSaJ//F5UtpBAsJV0Y1kj2eHJVqOF7Y7hJ5/TS0WY7Hg3Tz+MwZTett5ESEbTRa/pxMAwN
4EJsUynxIFj7px88dK0u8emgIsV108VQOjQA38ZxlSX/n0BwmiRfJWeIS3Xn/wYXMzkj8pAuZLgk
Dcm5IVgQ25M+Cjmzq0EGhNTiULw8+B2ppZeH8fZN8zteGCLw9FUiFh/DS9kdZj7MxbcbLT3JD6nr
l1I8o4bKsILRFjvdoa2F2TqqgdsI4HTrjerGcq1M8W2ono8GpH/zdHjClOMECa6BQvXGFfDxX6Nd
6doSa6NizBs5z9MuZA+94aD86Ip21faRvQBe07ebdotkFQvFgFAuBXhigNENgA3D3qleZ1+X9sW4
+IYqtiiuM/AbaSpA8sT8pRbhnQws70l9UUOaxjaUZdZYmGWJ3NKajbJJOnPXycyjT9awWKI3gxVL
YYZhPhcKgSEPGxHW0zcbBgTQaNUKDg1fx//10Upp2Ija72WwVs5sEet3no5GeF1xbP3Pna7bsJWM
Toyw3ZphMG9gmFnLRztenimEivNwDuLDKnB8kLk119pSCHL8QEK3DPKeBIN9mnvdX7jz235aNhqK
R8G41fkic9Oy31DD6y5jjHZzPaJnG6mQOu22TVXdpD5ccHZv3J4ABHXz+lbDABiM24p3cWvmyQTN
G1zeeIHck/h03Lha9HK0rNlvT7nTJy1oD+oK0s0cz3Z5/98cez4kpg2P/z1EzHpTl++11Ab7ASME
a1V9Cw1YQ7Ew2eClbBz43e8aGp3QjhIdPvKtzseFiHue9fnAGaU0q50ZpfQVlbkkk7wcvISHzPXO
KrPCk46eKs93x7lQYZQd3zaGlzaQjSQMNyNXnna2rvSjaFaNgcSRjfnClIu8PULlOdrqsQDalZvh
WdtkFYzUE5pE9ovtEoETFr/poUaSKRwcOHXYDdjSwZrjh7f7vkNHDUmgj9w/fCmotq18saF4E2AJ
HGFb7MmE7bv3A0kvLm0uImgqxsYBBqBa+D4TJ9p/LpeCdEVzD4hkqquYJuVvqIKf1zYMi4Txg5Ms
rcmbOwuL4s+JCI75MTQVo7crJyGiZoV9F4NclLLynyDE8UhhT/Ir6u6ei42f+xhQZf/6KP0l1R+l
tfQ6ALoz2h9c57Lpp7wESBFVZg+Fb/KKQRuQ5S2iKsxS6XaZWJJcBcPBCmxhq8l9rYrxH90YfMvj
zYVTb89fWNjokbWpPwdJuD3Xks/1XquSFZ9Llay/dbmwFLR/+7SobaVncvD0V3gH6tjBcxUUC6x3
pfp4R+A2R/0FaHsRcb3jyP96oNajnbrVpUjTGJg3Ka3c80e5qILHkBLj8EBd/iYZDaDC9Oa6e1/1
hvOHVW7NmDN4v2Y2nizsR+Z+eb1e6XOKusnUMbKpskh5YeH3vi7mUBUMrs3w0d4nSoyaIMRytCqj
5fokjg+4d9SJL5b3nvMY909qQQ6RqEXNlstE53UHEqWt6+XHZ7bPq1w0n1kV8b6KLKpMPSLqnhxh
KvF1I7pnqc1atts0YVNVwMehJ7G9awJSr5X/qPpwPMv5Zo2g4uHQcGCk11U3c/Y2n+8dGcY6P2BG
Mm19e1JKnmI77/xtuKxh0LITRpl+4wn+AkiYFqemKoOFwgpGUyNNhhFbdhgixhJVqJGNxP40kdPi
Aq1lI1d0tgD4ASQmGCCpfqtl0xLxUs60NkgqcrVjAfo7rq0RU/GkQs3R192dAdvzNY22RYNh9+jD
B/Rnh3urE7A6uFOiCn3ZpHdudCSUxiRkif1tr2VbYYIAp/1mq86u1QnbU94WbZGGxSXUj/nmeySX
jxPEy270ABJPXdZEq3F54u1r4Tf5vfYGgmfaaK+8UtCPg3RqL/r7FBn6lP3M23CUWdRzKQ/Vrmry
0oxfAwnELvTK9olT+vlB346uPnIA/qBm+2gmqyGTzRWBgqcVcJ+A/IqbqBNqKLhwsqCjP8txyhnV
cpc/VnL0TzPkKEklqwZ9aVmNEFH3cjjYnpRi1JDuX7Ap12tecJEnHEIrWVnlHQ5WERHHGNKU44lV
XFeAct2tuHIy55ydfTH5OWVmEO0Ewz/FCobMyiC4TREvUi1qo87LcdnpQmVUT0xnoKoX7ua3hDc0
1l37TOrhpjd66ybIn5uh8SHfM64H0P1PlDr28uSlfJVv9OpdlC7ihaeJT6QCzsEJxHMMKF7pYDMZ
jIWswi+hQnvv92HxIR8c6YzCXxBgDQ/IheL4mekcqJ5LOTc8hTPMFju2wFeIMVNd4xv4BhaDP3UH
5E9fXPcRbKwwQYAwAAXGeN1cwcYapjIg+P8f6HtysE31jwRj5b0EpT7vUHBg2mAr+8iYiYSyAtuG
MlrxJjRSSFJqvOqjas41xYWKoGNmceffSAKVi1v5TMnrmcwzxLsPQOPPjN27GbTjpr9mxc62fVT3
nsswd0Eqh2cVlb7FuZsLbettb97gdYmbZsF+wb8eb3QUcrLEBL09IKJv4OD9No3nc5r6EDbiuk68
kkEU9KfkVBcxkE7e9RRFrXtlu2fJB0C7HV3NJnliaNeQQm9sCLgV8rIROgyVzqmnwus6+7LDnfpE
sZs/8VpMm/y6XVdWlXJnqesVaSohHNtgcO9/EWagjFCaAS4ucUP/+RW6zc1tW1uBFaKWqVDFL99t
AjWA5WZN4ZUJsjek/APWw71uh/nldQCsI0ZJYQWDyA8xCHLjSqTQtmhrndUknlUTNBowKQvCdcUW
9Kg2PNxSig2bnqgp5q7ATG0fYNyxmIG0jLx40+uO7Ir6HRWUwPmSltXjdg+YEtvKYVD37k93zqbG
zWjeCsSKwv0J7qSMTWZrkKRfGmCOjOPBV4Y2Wv0uISEIQ5gSobSUEqgaZs70Ka30S6JzSfB8xOf7
gwQNUm4JZBX0CDBd7lIOdcQgRwB+h/BZEecLStDB6NQTwM+xoWn8C+JqQlwK9W6Nef3l7YUUUsNz
7vCe2KaMPyVEQGBgcvHJG4zQ3KzjOvZbam9tzwrlEX39mLi6VnhnS6U4CrH75czniqv02KRM8TWj
UzgCsTnNTbl3yDZS/0yBM5cLxZ+7iVdJEEP/SVAiRf9RDe9P36Kj0slbHOLsbR7CQ9kODIrtVic0
AkUHeE8eo6mrwEVAqHqM8elwgtAtf/Yum/EFzxhKWNI2noesZwyblXpu0ZjZeDaT9J7Binnsv9Vt
ES8ggAuzcSbk2LWJex+xZQNRTJNwEcqR7l8KO5q7iT7YWos+4fwcpGZAdRRpRglIR0wH6eRyMBYj
IuvUFyqQouTPz8FRW+UaSZWCR+MOfL1P9RLhJfA1qHZeP1oG8ilxBX5/nFuY/fo1eZLi7EZSXfqr
gbkjRw8+Z/QjOddT0N4WH2nrQwvyCI/Lf99wfcGLOCucWw8FI/Oh4icMev28F+bWGdsKmUVS3Rlq
hPSHb4VSLGnjUE8tdMITWZRIOLAcSxPL558/bUueuifh+cfEvPwXQLT9Ft2Q0ebm9XPthhGPYfbP
LL9eG5maMhYA5NhUK9fiiWlMxnyfYZalbz/Jt1eWGhhNiaHtAM2sr1Ut8sc/BcxI7EUE6maGPMC/
j/J2KaxXamkM7deLaNWVtakRSqE2If4bm4GbZdWe8FMRpctFkPno/TeMQtMKzHAIqC0ds9wzJUWg
FxKH2V+EjuDnZ4AsJaouJoliuOgiIELremutythLfRTWgdGSkL6ZuJ/2nGdowEUpDrjtJJQYxj9j
OAgOujH1rPoCHZrFMhXoLjfK88Xsk5IqXSBt5M4u6H0M2z1j3vUNP4GhoCNst+YsL5f9Wk3NF+hd
aRMcN1mB/9Z2+i4e1ZV5YgCJ9ODmVNES6pJm84xt1xDuWt0eN3jGiavblPPTrEgioaj7hXhnIkAk
qVnrchTvfrAY7f7cU3nf0qQVCJ0MI90X11Ulgz+BRc0c/9UaUxPBAKhaprUDe9d1O2JrzCcYJuY3
HwqNZNOXyNpxwztFtk8pHBll+zAHvaYgxfPUr/ZJ4tzce+31vF1NRR+Fm7mbjj3GnhDzigZopt2F
GE3/pIC9VehZr3b66yTs4wofYiaXrW1We+jZb0kTyNYeG66sUI4d9+/N/EeuCOxvEvzoLiYWcPGR
uwfVyqDpWKSrB2uriSmQdmlvXZlmTHdydUfTmXa0V13JeCG6nhpRuaTxN8ZJh1jsy2lJvK3rGFq3
o3P5FA+xSxW+CqB8h9P+yESI4vkXVtmPSA4VCFU5E9qDwhKyzc0KmAdkQxO8HcyMOTpLNCeSDhoN
/2oHUuLJiIg4bw9ndSkZiZC2UFzM5iLTsI3gcDCBfRe7MjMr1XFzunMvewlhvlBuELBNg9ChOOwR
ZtFxkedghFcIqxrMTlImTtSe5QCfqCjqGscAa0GUy0sCzncZ7dk9L0slI5aEv6VgWDLDpPxtla7J
9bzl4nY1jhr7lRAtG0gUOjJS+dIIqtqWHrIsA2rot7cev0GkKcjTPG1L+bXTT0VuamdU6aczXB7k
2hkbAprClXQXgoX7/VtCl8wdnBfEJf3M6YySzhiUOeZb4MmB5knPDEHtA16OTSeKtMKXHoLGoMEj
jhk5uiu+7ofJ/kud6LWsbMZOtFLHTSYlX7R68/eFUkoP9mTdef1WUhmj2TnJcUItvhWd+yeOlJWW
ybdOwx5l6wIcD/ozMLU8VWxqJir4kz4sIiufNGqjayUBLwMDJae3UAahKR4RokPuq1BWIPKwjwkZ
JpmPOD+0EqAIO5xgVSy5XGpiWkwLYPHBlmO+wnH1n5NNoOmGE31qrRrHQn7gfduBttBDpC/keGMg
hiaDGdraQ/TRoGFSF/r/+VUeoZehl56ICb+EZEfBNoYDUnablOJ+xDA3Wg/7+PR9cotXOX0epaaq
m+xKHfgqQLKl/mB2U4BXdl5qfNtLKlxNjZNQxOY2E6DaYGah/2if4q9veJ0Y73tw4Nk04TWtLiTw
ayz+f06nYiI0VxQ/nBPEmpIHzfmrbnWqkArTqlONSuyEjmUT/DfBjLZ2i7mYkp1jRUJbmftdppHF
+LBUVKY3Xu+TTUHZzdb3WAKEuaR9MwlrkdQ6IZPOJ+h7FrnnDUIOIgolhg16J2vttectkWLXpMZU
sDJ9iHttAdXInHWA1mjrHBNp/BUt0ISCBMrO9yqCuMBWuDgSt0XNs2qKzYU4Mw9AHhZ54vl/hvkQ
GmB6tbYfvRmqi1ZGiW7hMulsDa7FFWAW00OUcIy4E569vkSqBfo6jAdmeZeyfUUGPqXxDTO6u/L4
L5Cs0+JRFox2EoFWoEcealR4YRSj+inZoPNkKJwyi/LOxVG5Q+wtmIn8qFIFtbn912s+AO0niQ3/
CAS+nuSsO8EZhOixeYD4gIqZM8WjMRTAzgR7vvh/sdShwnYmGqyHT6h3EAWoaY6JpyUs8fYS4C/V
Y2ufd7UAMU95WX6ollzW94S3yhT4JrLAKry4W+02zcYI0kpKGvQ8uZLQrVAMVXk/z9YpfenmzTQG
jKP2RGu3Wg8vG4uRpBIUjxY1m8ixoPZn5CFq5iU+1k5hPjzuTnWj2YduCgmcepCKaOtOyFljC/za
OODMgK8eIPMp2WSQBYurIXyEozJhzUCvij/xDsblUuXCSw+fCOIeJkTVGfkHGYH5U1FUR6U2xXCk
DQWDH+YVct5iN0bpZayLtM9Wyj8KhkSWmHXmD+3uxBm7nici14pu+fgxv6I5PeunqVYir47lUfcA
3NfGuLX5u4G4+nJhPRzos7AUlpoiAzLpvoJYihD35R5izfKNDX/PlQWYZ+J9qGGU35yNeGEDnrnq
hYSi7BFp4Gka1yamyx0Ef8drIEGiVwcd3vKhKvUi09z5rgtYjHxZBY74cBJ8GK56drK4IajTUYTN
3bAOIRtrgAdil2033ICTko5snNp5Bln2pD78DQYmLx1V+EAvGhiStiZBs4PHtRWLw+LDSQ7uDEM8
xXZxhRS7vCfdSYZWWJMCxyQimRK5JAhkFEhB7Z4qbq0/N+ESA5LlAkkWLCte6xpajWkVHBLpWuRT
fWEnkxEFYBJJWyRvZLKF1O+nW/oQnGUwMvjW2MSU/h3Rmd5muaLzaCbZ8jJtiJ+03mVU2eVphm1y
ukgeDKvNNyBVAXJkKhmZBby9cMhAqwAOHk7lqt6rnAd1k6SAZqKA6Gf59/z5L0hxdeMaRL08QDfJ
TvRlLRfh0Fn/QjhhECtc67W4Qv+vgCkoYkO+Kz5aNoE+WQmKet/eC6uG1WhxaAGg06n3IbnlPB6O
k+5hjfGdhyrrS++uv4QoJBEytS4YyRJfpVeeVJ5w3tanHpqIobqM3jAr880FMMJ2l8Cdp9eYW0p3
jgpF4rJH/9IVc8GFfu5+6ASPKnq3FtqC9isbGHFzQU2QomGd5beAHda7P0+QAoz23VgrwSNNYwgN
UNkaCVYeHq8D0K98WrNKA19XdayG7lZnov97+98Bw3Z46FwR2WCIK+yBu4gxSGxkFEdEVZ5fBtyw
GBsEESz5B82Cq5yP2c1RSDA7jqaRkR0bDu+6Fq3D+iiHYLl1H0u+r2UJWfzy9xWHJxkWJqms2GZb
dV4FwvX/+xmw9mmrHEXgATpAmzx0LkEWYuoJdcEQfIe9JaaoaEFWtctbyzZmOW4qEmCmsltjG+sZ
BqxbJM1mykXZdDTS3yo5FOqt1tyDth5I6TXWSILb9f3kokZkVstG4bLNbNIx7B6rC2sGng0ROmre
8TpUM2WXnSAc/HYRmSy9UY1eQfG1xMNafGwDHeyOPbl5Rd6/1Bav0uqbAibjKBeAX4fFtoKhPira
vL1H9YTfxqZcK+U0eAuxn8DqJwD1HvO9QgEn8pMElAMypIW/ZLGYeZg6Y0Of+uPKUczr63nspn1r
eFVGXsW+aDwiHh1pgS2GZlnSnPQKG4mG91M9Pe3+7f0c81RMoE8mAy5ATKrq2rba1sZ+nQpF47A6
OI+0R5/HuH/bM2dcwOfOPvbI3PsD3aAUIiLMYcEz7SoSXfIRDcLWCDhIFiyG7OCLiKGy2Es7OeHF
5M2okUvEMrSi4velfLFSDBa+bFpjmQnR2aICCU4XH5NwEcCTgtsGi94ieWfPBAFJ3aM3hkTmTYPb
Kwh025glr9Lk6+xknVA9q8Hbyi9el7xYISlDQ4/nUepPyhXMOtbJ0fJupjZsOHyf7jCcPFfRxJGw
cD7+ZjxiKdniohP6PcAy2EN89f0OexzBL1GKftzs6J4AKavMolbgXxwHcaTeF6n6LdV38Zp+Yj0q
6q5Z2mN6GO3Let05kGPRVBvA007YWk+WHRwPF+/2hBxTXfBG/ROTs1BiAMQgHLwGEm5O4aSTd0M6
UWkt9luqGfXbKisvNJiIenDj5urIjMCksADvBfqv6LDJtqORJ9zA5o9oupcYf4VYZ7PgIV7s+oH0
PD7/chkIkbrhrnenkbHI0QKdXECffuRRJSImN5d0VnlQcDe+eyLtpdpSqGKxOD2NEnONhSYvlXSC
M2xYEvil6QT01rjw7HRkB/4nJad1XGRVo8kpgcAimhM/CCX4bErhh4elkV6xX5+yvW4VG+JBsOwS
27uHvC+z+n3yYuR2x4hnKVz2OgKr1liTrba3edb5/UBmYH+wMR0Hwxrz2W819XaBsVVsoxHXoOSW
saoKgNkypd1ChIdmnWzDuzN49gvlm8qpQbgiJpYQN1U6adTOsilxH0sc6UTTmmSMsg4Qr7YjoEl7
pYVvrSqC71Y7GO8X6xC9LxyyDV05MDaWz8itNkeiXs8EA4nGgFS+a7G3RZfmf+LoJpXoDSNfF6WC
xGJF/7GDU4L+xPlhfSr0CX4TWT09J/jTmYWXNF29lBbU9xL+/AqNewm/U80UUp8BHTIUb1DQ8Y3K
JlY8Q9PH9JzISJtpbhn9SBjw6ZkPwgK5LoYqItxXpL9L6mu5SMFNZt3tA9hV9bfySceQAV/kBzQi
+9SnN/JPt4XId3U7DpxV/L9kUM8v9hb5S1F6e8dReM2pB0JGkSX1JiYUk5wpwgz2BofTDOqUSl2e
Uk2hMC/KnfeH19VqlU3zz+d9JKBNa9yaJJ+Vj/9RxBXYFPumuy71fugt7DsJS+sMzTuiRf+oeFQO
JnLjpDoroDu3oEoncT1pFHbKizfwcwLBfoOlEwtN/IXigpMUPMLVMm3VgDg8KvKHSTQsgOYK07ZZ
28kL518dggl8rURWbCuFM0Kf9E9Ry4gNTwqyVEXOFTAMZu6Rhm/cAnJBXz6kodedPqge9I4Q1Meh
qig3cusSGtboQJRJUUey6dg3AbNuYn9+/5tPdWer2ujTnSg9pYIeBzgNqbnzN7dpEwhTSF5sTJsb
0gukztL7nWWYLPArqO2Z7W5Ni3YA2kBafPzRva0njwocckskTm7vSdf54c4bkWfYAuhShA8/z6LC
YJgVx4/VVfFGrbY70covC6uEe+EintqtIfIQt6EckfprLb580XmyNrWBoHRl0uMzjNkze7NVqo3B
LKXO3ZA+NK+2F1k4HmSx5UMTCxcXU2j0b8qfVMK98aSTTLD8Fo/71eid5mRBQtJCXYdS5KP+Skuq
i6vg8IzW+gKTshNMAV9UgUIf+3OXYQjwsptDUOW+OOSPcb0weA5BdFgouZKV2YaiWDo9+S+rvNYU
hBVJYe8WKaqSeb9tTuTOANDCSYdLjfWIoEr6yjs/IqG77tUuDcJxH6Q2qpu2hB+Z0aZGbSKffyxd
JnPAt2E8E0WIfgN8shcy2uzX7utTvcTYSnMwJSNXxfP0X5raSWjYW3kBIzQB0cNulTDVjW7EjNQJ
2wjf1SWjoROOvPXjq0Nh/FxysSce0E9tbti8sypjLu8JAm5/gTExRYgVeqagl0HyZANrsdokMFD5
ACAxRsopX6hb8uF05J7fjkTgb0O8aP2ga/JIbLqZ1qujaTLDJXeFVchflY3la7kX1JOgr6zqOuN/
DHD2aYx0qTGWVI4fH8e50c4XqXLT0kYFJheLCj+Vj1oDfnKXkJc+l2AdCF4dDwa+IpRwVDP3h2V5
gOyuatfNMONfJmPQz97oFNev33HOJ92MLonp6uHlnmly2oVGdIAhTJcabKWeXOWr95c1dEeDJye1
3ezPtr7sn0qT01rxDWwecAFl6P0CFJe0GthSfcfZ1wCxwHrNOIlXNVPGMiyYRa0t4Fw5p4/VBOck
H0JfORk+g899CN9kHnWZRO68iUdrmkJoIFR1VqI6Vfp7ATPWMimlGtls2UBlhHVH5xmX/xKYoGxo
AQ0HWeb3/ggNobkVgaWu5suzhqXbwjtabzYfW0U0YbxACdahBjfkgGSPxwDxcZJu75ZjRdwf1UjS
CGRE1DyEeawiX5hdAsmq98TeZSs4s3VBjQY5izvNIhR+wKSnSwLq7aBxuOs+Psm87VZ94LPDkrn6
zQZ/hpNJoUB9NTVp8z3ZkXYuAMD5BHazzVQCTTLB6pM0cM+Jn0F9h5kPKWTjH/2R0H5opkXJvi3p
mso3hBYfAi10w/BlooBRyWl5UoQCRxmbimODYSe2zfc1Jik7LniVyQ+vNYEZBceTNeMiDEc1ld+u
FCZE/r1fQgoP/F/2WE5dlWSgqJPlYQsC44Ug0E013QewHStz8Igs4to3MAe8IdJgYg84PLLahc6f
pzZ/ZB4yQvLuxB/oxqM/He2100hvw+W9AsTnqlDNPsQvnVAia2Otckv84RQ7fnJiIWEOFUz8/XM+
zQff4L9uEt1CI836DpcizoWvNlGSpJUMaYylk1feJuLB0qdVXaVtaVNi971X1MzPm/QntVk7t6hR
4nWQGZ/luertQpJEHpL1lJz08N7slwVygtoh7241ZagoitzjR5v80bPgWCYe13y+etjQG9oR0dZU
Uj8S1xRTc/aZZh3x12avETHqVzfFIo7S45FTW5FDxA/LFH35iSVbBVDwk8yZU580IWKUTPsLpvM+
sN/Lm9jRyeUGOc6X1LWsFklnPZUegcJApx9J0Bcxvk25aSA05UFYPc7mZ/eKtNY8eeZSnhDNNQRC
UqnHgRxw51kfGEZnU62dgCu8g+8AEmKGYP32JQB24myzTBgBIHRq8HomPSO5b4BSsMaSVJFOiLSs
lz6/zCQcPw2qzG5bAl1U26Tti9Xe0NmCCIYEAa/vBEbsjd1cTSM7nx+rfsV/zRGYyYSp2J/yC2wu
bvWJ1BVfGdZusaFfgbPQVc1L5znFq5PTVeF7Iq3mhstw8yau6qVyquSMUfj0HJTEo9DGJJdzb4O3
8hurMxatQAIcaehH7iloPmEI1LFeUvzpw0ogiqM/TN/O/wX5lT75WN53vAoM1fxhvBRZnoQDNnMY
hSSnnGuYTTkODJOp6pTA57PmCHxh2aSPfzC7xbXsI5Po9ua4epokRQ3L+nzgXEw6N1vhw3hZEGze
JHE42yFQuAvBwIwwHGGBOTDDfwnQ3oFQxDQvHq9HHQWRPaXzlwicgCk6F/GnMzrRnpLJI08cJNu3
9wHR+WTqbdwKhVt0Vt0iC45eeNgIYar2tJcD+U0C0no4IPN5NhJPRHI+KP9F1rbS1Jqm9RSvSQbf
+PnHqjLb7PoUkoeK5G3wu19VoWs0PIEosfOaxgcQkURYwxALGZYPrPVVSBIdu6xGXuaNaRzYNfX6
YxxcZ1sMtXSdyBVLTq/Ug21CkbNnptXYVTFJQkLRyJrDt1YhFWnSIaJHbzWTvc9hV/qchUQggXqf
Rt7W5e3S/HaDCAHoZ8yQrqubF7RFRW/gkX97pEjoAo7j8jvAnA9TvDBAfVCGY6iaIUNjbCXUN2VX
UBW3nXtkumnonoodOPSiJR9Pipj89e3airwOLAT7qUn6x554UmOQsbD1ZrtKQp3OQk7TEDyZH8sV
eu+BVwTOk7LJTB13QQcjcMCbZ3whSKUo1xK1eZE/YvUAAenIgOgJwIVD+ojNWRIuY+Zjb4LRiMH/
Zb8oJwqqDvQuNczaEWwzqMgq2hiBAJnhD0IbkWgwHwkj8q9ErVoCMQQ9i8PpQTPN6JuKZAYbHdwF
B14L1q9ZAA5P+uh5U8LTW4/qqidNPORUZ5XSxk1OTqLnUSO0rpKdsJrTIcoD5SUFx/X/hf8gCi6b
yqg3inQxyH+FaBJRJKS8eINuO1yf0eZwVj5f5TZv/M6QmM/EzBR354pspicaK/kiUF4pkcPPWr0G
4/UptoSkT0O1E39buCAhCfb8pdn6mnT4Z0DjF1Oy1WoqyyUppOoGhr/DbITYa9F/UFKejdhfmvt7
LQC3ooWP8tfqFovusTE82tH5U1xglOClYV1pKlsFn4f84QzQjG1aLBUvbNB2s0fVvf+CkSu4zy0q
qvmLM12Zx4q4kdv3dUKJlletpVJ7XLPr1wyM9SDPzkrw3cx7Mlx5AVcg5TT1St5eLt6ftmkE1AzM
B/jeljrFAubTr3y4EyMn5K93yLxVvopTqf8Agj3fD+GP/zdo2icx+aEf8/BKL6rlxqU9QRX82MJr
Hf/Nfp1YNOYWsW4u9zVbAasRkaoYgUsv15by8mT1IvEE0OyQwRgr1Y37BeTKPdWeHIEnxrthWFDG
poei8z/+FBCxstTUtnRDYrZuBFYLGCZvJaTd3IHn8bvxvnBtRqaBaTOlcjoqRmeQr6BgjSKQ/eyp
3O4CH4Fjlfxq3bkyCXrzB1QNwSTe8ESzAONONyhKKt8HE9Tqy9mNCoyyDV3DGvmtf3yPZ02jyum4
X40+7+HfwlOBOurbpA3bjKEqTB/lF73aduBy9ZUe3pthppe4M6woroZxX3kdiTuYrgTRJuUT2YCe
/8ArKV/rlslh8u7MlxHBZ2EiF2aFURl4zuuklcOffa/S6UB+hZGE9xbNWrgvxqmQceVf0zbWdbNy
9PPLca9IDS2mXVp+p2LyBWxTNwsfu7v+UK3rtzFE5F07MHIAbl265q2jDeh88eJAOd7OncLE5N5d
18mtieNuMTZo/ZjnZW58AYTkUOy4juDiGgfmUueE+3JooLau8IjFLKb2Qm9iB40EB/Eem+qVoXzB
ZlBbNPrG/uDXfEiJW8gzEYt8oprwKyWOAJgASpwl1pfkqHCSSe+6Krjlb4oOgAT5hdb3WrZD+ZCE
YFPdSp4aqjvMUDlLieUtt8Q8yhqQW3W810zfdTTU1xYw+3700ublvGlW0lyg0DxEwQ4dx8vnVvUL
FV0jjtOcqFG0apIt8m7wJT9GWcGSez0Spsex0Nfy2zGEWrKY6EWzmaRfKQe+ZMnCqyNXPeNeFkjN
CyIKcaaafwOZ7E6hMQXkeY+2mLeuhWDaTTFws0S5k4M5o4n8c6E6tbqfw7udA7zbfDiLZ/OBnj3O
w2yRECAdnl+GRT/UvfKqB8qGlNViKYmL07X4Js01YoiOOMk7qhbwj+FKHnH6h4D5AIinnLx2GfdJ
Sx33I0V3OXo62W1EtKWQ2wK5GK1rPNnNS4wSkqVidpGdoRpSMqCJffLopuRtl+MpZkrMTPTHAggP
1vUcjbBLR6qKTyRRMRLUOeSXiN9ThZW5BAhi8V862XC8MPr+zeTOhk2tzIRKElnp2nmnBOs5J6q9
lk3KD7jEJggxsybfWYNCZcF8w/cWllIiOBNHqaQXkTj37+pGGd8uRnEAnx6InKS+PVmI5Tx5gwlD
FkIPb39kDktZMuPCadhjIAzp+5y6AuNHL/EnxS+KUhGTvKpWGQuObBl8Xdlsoa6jw3VBRAyXu/DD
cz4ZbFrUbxikJISLbTa3FNKD8qOaLa+hN2mc16+TulTY5fBiCIlZuUjJZIlaj9dBhjANplG8Fr7z
urTWDeQMz5VD+d32pIT3gBng8COobnCwafhtx25FS13wo/uZim6AXg0iSEiZDKqTxcf3pG5qBFh5
3QWCTEqTivn05bHDJDc22RPdR2e0azG6PSaBNrNySBEFZS0ek6rhg+IFz5i5mJLte6DSZQlQbq+g
aEp2T+Go1cCWSchcWL2QciHTHVThPYhwumklGstvSJgtyq4qbJqQHAJRrnZMP9du6tFgC/3jrbWn
sGKCbdx9daOQeFsUFhl1SPZtLOos1JQdtKmHN8sAwatD6+CXFOq4V71D+TDHhWQO48uyLOqB6Ofy
vn4xUehVurZ67hPy9nP05qgvUDkWtzEZsy7vN8N32hvvVA0Bi4KVrNc3zjbA1ZDJlWoZRfbWNsOn
gqStmdyQKOHYY+MlzZlq+fwExnaIJXuDQ+EFRh+FgurwqXdx2f/tdCpHafnXPMzP+b65RvKx97MF
L34c0Ap0AXSMLbJ4wspYv5FWZxyXm56ju2QfPh+M69Hof19glKsxYBuA9mIPrey2WPeXAimFM6wB
nE1WGmLbsD+TJyFrZWDL294OU4aod6/1hyqyVQvOrxHtHv8Ol/eHrUNt9qZocXC+m9HltYIKNoYW
zQWxsbBOv/e7i7xRsmzRSEvBRVgeJxalsPvF3yApUMGkGsK2WmQpoKCY80LEPEi2ZNtNhc5nwqNc
OzPfAcWWMcEQOIt1L/lr4I32+nwG8KSRFwd3piCxipcRKlI5MzGkTaKNeMiw1fq9NdhCvLZsE0i/
g155FLEHb8d/nWAnDCR51vBaxn19vuBP8BSHXrGIk48GNdSngf5SjMXMxLrU28GEuguEzDBkB8ot
B3iXtFiFxBXQSYiuKtsvAvXi0KzE7GsNJX5Duu3KfzwC97B08xqQWr8JB7APVGbPUMsVANWfNqgF
YuONOLSbPu7y+YUTKVGD5rgvLyBd0zBKfdhlVXKvz73Hbwdg4An/gJEJdsB0+Gru5ZX0q0AqBMtT
a6VQYhwF5vermY7WwA8g6ctlL0qpFVDvrRmUzEgIHRlKo9A0SQ9Hr9UKiScQ8b4yQoalEi6SlMms
cxp6pdFRVcPf6yfFX176Ll/mmnu7DUiodSaCLrEZGdWeShK/lVW2J+OOSupHV/PizwJnQ3gmPDXE
BaaA02lItBdhoY46aVlgoNeSjnU/8rWK6+jLu694SELt6YQho1upPY3TlOUREyhZBqL0AG7aPr2c
tKI0auPI6/ozKETK2ey8bgz9BC41kYangfmM9aAl+3XBCWye3mbJ2zQqy3pUbw85gg4xVNKRR3v/
mzZjcmDq+/bi0wZiVmCA1QDmx5ZHUHOgoPNEEj96Bx5HfMu3VWgrtn2tNandU1UVw3cjPsxLFPBb
6dxglTZBYmkq8pWbiNhEMULA8/776z9l59OxSU4RHcfz+7M21pG8rICq1kCU08uJR7NiCWPMBfa3
eeSxcbKUX7d2mliBzEPhT1Qbdat2Hswb/KOBiqtV4+L1fN3sfqFmRxW65L8TpWp4xIKyoLD9ce0U
QxaOauCF6SCpaQfBHkESX+xxcUASSivhC452Oqs3B8wNqBLtO4pzaYxhGXMvLrxNfFObLmxuOizJ
LI2evT9oyNCJgZLdr1ixyfzasIi6zaQUFapU3WKMu2Jo6Cuf1hOguVHs6liCVcvuPeDFMkPc06fl
laGDC3Se4tLC38nhGUdtSHa/rh3oNfrPmCayeNSgPLpBqLUAvzYqgwJ7CKBpkkQRWfPMVy7Awsfc
+r6ijOvuKseq6g8e+y0Qt1UXMAy9hh+9A97bPf6YHs/PdMwjBLw/JhUHUYa6aePDGdnXSZLPjcG2
L040JFvvMVoWhFFdvaT6FsWYlbd8uxYArFJF0Qmm0K6Xmkj5tWZ5P5ySR0ZF7iEABQBqyAHPYXPI
4mNIkAX/gLuJkS3z3tEMBueyLAqqRhovIbrFsggKpOK/ZK6nL4gKhhu4xN3juUEaZlNPJnz/qzUJ
Wiiyb3kKicuk8CbID/LGRrWBSagbhtS3lepPcrb7PLL4jn4Puiiw4Tzj2PJKv4frGcZJVaR6usly
2WSBCuvEhpLvUQDbTFhEl6FNW6YJGHyQ37wlBdZRurDQASFriXw136RKypkBN0ojWMu7b42CUXyg
zIeCqs/DpeWaeH4m/S9z8IeSX87M94AJ02q+oO6JpS+D2TZ3jqmoz7r2K1gApM0/BD5jwG/L4Hof
L6YtJYrCGGCs0opoHa1OfTGCsb09wGIXhXUPxQs/3MHmSEjLPiCh1ro7BBldRd6aijBrrjvsMqdI
QshorYePvB31qHsKPYztfh3SrxM34Wa5kGxQ4po53YPZa+hYaB1Zha4F95HGxF/Xpe8AEuv9lfB7
h9h3AUVaJGM5Xr0FvAkPzCZkoFesWKu32uAiTcTYPIvcCUon+kB9SS4b80nNVbqVZGK5s8+5GzvN
JbYqNERLh0KoPlVplM1QfG8jvfjLwQvRVextY7gMLZ4IgG2gnLRj3NzfE3kjTk3Zdbaw7wdq19V+
0c7o8P+LC9M7wMyQSQa+rv/bhyE1j+W6JRGhcoZyJbWHBSl+7kjPlu45y/sIyt17u4rdG2WRmcuP
kiAYxiM9b6HhrgmI/jZOHfVmNCASHJVDtSV6/mMwXXR9WFtHvQ8cQXdFMnSNk5u2I0SKNELwaWmB
GNIDsHxbqfyWMbITODUG1hHOI/6PnrMdnYwCOyDejOctJO+FU2iO+oGJsPAdJg5BXU0U2rGC58DT
N9C2DGaamV5R81h/yoReQ5/rQX+R+y1Vxo0jUsyT/ttj1T4qr0pDbczFCC6S7XxbfFWRfxZT0n9a
Qp4S+dAmCms1nUGEi4n8kNUeFwQ21VYnpd8DBAVVKzU3lyrIzURkzhgHyfW+NtVuIQQsrkL20ZbI
gjhMlnLKPQLnI257bbWjO6AfBIH4GyTZMT+RtEGyrPJIJfmWnuTjOEXfPHgW9zLgFEs8ph4BH+lU
wAvP72D/vAnBYvJaAmx969yMzWGLXnGaJkPVdc/Hw9tzk2CHw1NkyCLS6amEjLFXoYdj0407cL91
JQeye25fiZwaRIRQp+2tNARzxIjoYDI9Y93vDBXf2cTp3B3ywWo+ZMMgqGqGAyvszU7fhQsvew0i
ZYHBuvEu74EsLuZuotocE1B5X/2sui18AcNsM0cqxUyH1nzcO6DhfdLI43fz80RGkshLHbVvIbU4
Uh5PPaiUWwLhNmo8vhorM8TDYY9dhUk/cdWY7VueWhTugjvQLx0PwztWPbGxtFTGBEjh8FiZw+Nu
eD03ovEQdMwClBd49MATFYwCYyDN3NCjn3VM5O9miZRJusWkzGc/t0FNUJoNyLl9VmbAmalviT2U
lmjWbJzrtfuu1hkiwikfLEcMjilTCmdBwLV3oGZBrgwp0ZKYYA2eHv/kqqrW6nRxBK3Viq4Og5Z+
plfBWwGffjl0vDaFFHZc+o//jv9vJhtDMu5D+zqdXZGYdxKDlllgiXQv3ngCb8k9gTe1ha4iz1KB
yDMviqU/JHDkQ8UiyQ6C/xwC0lrON0MmzEHGbQYcsFlVqzgJBjwTjv1ZjYm6xpGhgPhUlUUHBOzO
AcSd1orUrr6j2IQqSJKc6jNCsd5L11DXR15OxkEIrC9yWJMY9bLK0tWLLs59UIJHHpKcAqftH0XO
QgrnvSn+G/UsiF+w4rTsLfWOh3ydcN2Yx7eFd64p+CeUUPWq51veL94yOVDkLsvVMhOA6uzTx7Ue
tbkMDky0M3qEDK1JzSp0OlHNgFjDsh5w/37VqhOJfNIpDRhx68JXMIwE+bpszUPhvXyvnRq8/9mR
HAbndoM3Eq7sPoKkSNGfvVt+627CL1fWFs2ITlf/Arow1gUQkzaWRMs0JkVqcXh6S5ClhFgtTSv3
L55JLZPtZcuL2jQZq91kMfnuLI+qTmvP76BPU8DWB97k8uw9G/6NDK5+994Ykw+rHCkLbbo6OTji
VLLbRea51fr382i3bgCcQAPQV3zp1lFjWZZE2FODFOn5ybHzEBmooiRtIZgZ9onk+2SYyUEBw0XK
KqVLGYt/FRxSTR3PEgFtjLnzuZIvu0KPmdR7cr6gzSK7dyJU7tUkmBcsUJ+OpmeQudvI6ycHwpCL
HLdjkuH6Xg30bmHk5GyVOGIt6AMmFgrDbB/8dns8r/j/RsXrwRVjYp/PlfOQFV/VHXtObr3CZdl/
c5fYiqOUOTwtUns1/Pi4HxxW2djS6JP9splymMeUfCyJKF9H7tcjtqlRHaSMNCazQziTrmGndoDw
+EzNvH6Y1LxdWt6+y1LLZkUaZV+XYMfYPGX6vZdHMf23u4pWEqVcTk/pvoxkMrbFEeYCJfFpNkjo
KuFb9eiDrAUPoHyWkjZ3BtPW4vPc474/xVdd4xfijRSUe850Sa4KPmuoB+2ZoypuSc/2EU/cwZnD
0o4maNIf3Vv0CFVxjcClxrIBHPBCba+sNsihKYRukH+fR/U79XijUx06alcgjGu5t7xAYHzhjDwu
NxyAeNTxqpT8cM3tZlRcXz/Sj+TdmREVDaDT7tRHdDCYqWadPIpSkkK6twGq20UKtCpjf70WCIk7
HGRqXv1oBZDR4jT3KNi2nneDJs60y6vBNjsQ5wBZVTLb5HYnFRf2/ZP1WKqV9FPsYZPybuCE0fx8
mkcJW4CQfOtG09eW6BfowWGaLBjFwEKvwUE/2MpH7WO5lZVGohEZkScbQqoh3BmAXc4HCb/J14t0
yBgBomDlJRYIK+hWmBtgtWpi7jf+fYi/XSstoQnFVZNJZccGmQFcLQXWDkAyszzJis9a0fVpr/s2
2KHJjpQnZAdEF3g4XfDim1hl6k0zp4vb7L6DWy/KrGa5VeCZiG2dD+uV4Es1CUBhWWJOJXbtHfvc
3lEqt5g0L+OEcZY8aZfyc4vBVpvhMnVU4J/PIBeyOzuIw3Th/q4TZbxrlAq88KTVa9fYGAHNyyh2
uBM8/Jt1BqJXiU0K5sbsDRUkG2DC99DtJ7qCd30PB+Gxz/T9+niySkhbHobynrjMbqF366aXWZO2
6ehYMdM/oCZZUYlfC/oszYFr8VoT2W3IJe64BjICWbGg0/bNHg530xyg1+H51G7DiwLPc5t2tw7N
dQx88SIqA9ILfBORUQwPMFzTJT6lwjUMqJ8s+Kf1iMAmcc0Il4S4Nlj6rrFoI4iYAzvowJtVBREf
uAgq4o4sBi3gx3zqjlQE47hxmmH6w3WhA4XWaUQB+xZDHIqQ1cl+rsLqngc22BJBAFSk8IgBFnWt
9UhFHpn7vVuYv457r8SSNrG+WE7AIJKkogcvwzI1fKmcvQ3U2M5ZgKQADeDrvi0BivFdStlH3ZHe
DUpJIUb6uZRr1+Bj0x3k2fc8WhoH3+N6MoVbgaWsCS3Vi9Leix/BnrnfNbWhsx6XcIEyqimm4jhO
kM9wTGSGPO6/zcimvrehNmFUWt8Cf9rk6S9LGnDP+RT7GzCisyir76SzP3vOtNxp7bsHLgFa1Ye6
MoiwTIgYEVIEDfzhw8rZKGKyT/dmSbLdoz8nV0L0fzkItfvCnxDQ+qZZinCXIq+UrVVoA2Mo3VKM
Ff9LPCUoKOa0R/+JzZAtXPYr19ql+6BpA5b03n0BcyhysBdBmi/Mb8nkX8ykrGwWCZ9AwhOS/nDI
pgcmKk2kK9kyTcvdMdcG3ZhKEk/PAUfl69R83zCWfzysjQ6cyT5jZJoJPvfhF98dOUqk6vWcjR5B
jihMVlSuDofMY0E2MDIdoPTil4HNsPefWgDSx6+5dM5q20MRJjd5QRy1oxO8WzvQaZOfu8cEyErM
D5HU+gHbcT3dkQEuSQpjrNqk6dV0zCGrhy3vAbz4JFiaQgps8VDcjEu7S+bxHjhJDFDO8RWv+pNu
sdpM/UjGqOEM6q00LPzDrVoAuI6fXmFyxvliaK9hLOWmfiAjwWQVoaTj1pBrNysQCgFwVSe5u1gy
NY6+NpuQOjsf0hvtRos95m8qA0Zc03W3TDJL4CEknWzXTiwS8X5e0jWKyAuUWuGnu7geVzReAINs
XebRT0faj+0m7t4oIVLVQ4JtxherRMHK1dqFnQnyX8EmxFkvL0uHf24AAgEFEwB8XzHyJd0kmmts
4Xn2Sq0ZCJOD9uxbJJCZ2mtDA2+9gUEAED9CvWc/kRpQ2PAlwClRggHOHt9/KFio7n0aUgH37esn
MG0gRPJCqrtJ0PaF2LwmQ6uGLwdVdMgzjDISENOApN/iu4U6qPK5fPGYIElqDy3UEC3DgAuIhU6D
cp+mLts77to514lox6qig9HizG4dAXER/D/GCJM3KQA43kAtrIM4Ji/zzo1sf0JaTJKfVsVahPec
uSQV9wfx9GS/WJIX8MQuxce20XoTyMnBzyVDEr/VosRzuPuOtXrasMz0vCtC1Cnul8ciAYgim+y3
nq7EwpM5TlHJLtYyE8rA6Osro80gwhULlrx7fkjUdneqLpn0OReU+Wmij+6wftN45rQpl/e3Thl0
ggsXsw+dG/wwzIzjLsrzpAPZqdgHNWxD1MSdidri0ZopFM+YGBmLYPYY4AEH8MxpxmHm3kDzLy0r
bKfjSxDeBQNP3QL6l4khX72HDL12F1nE4dy2WVAeCfdo8tFxG7OEvQBjp6Y1acSk+KEgysq8XEtX
X2eKsQbdNfYXHLOcU1hQbKIsElBR0DoAC9rEowjee1yJQj4mZ2ycv9mI2M6VaDzVVfkxSCMgr77a
GGcdOJD5XihCgCDteWizryG5CJ/svjjg7XTdCCbCKWLUUt0omnuQTOnsWHvrZWr1m38aWxLNiir0
+msBZIf42jVeflJMh51QdjRtAOBlVwOHnWgABQoZhmKSDuTmfqg5jniJHaEp3pZ+sjHd9bSn4Wjz
vUj9MSDESNVEDhXbzxLVxDLes2pKGgYMt2SVzy1Z3R+ynm5cRTMtVDEGt64Xlw6JI1IAtNXpZlK8
1+RIX+uGJodLMw+Bu2subeJKZJ2aPff4VcWdmitXl+J6gMikUem6Hmp2g3czjp6EKdDdpw4UJakk
PZuX8J5rPCclk2dlbJHVeR53N7gMRqUL9rJKKYBP/lJ0DtW2/WQfs4UzLRCnzVBByHhiJY6nidRa
Ihatd1onmXHXfdSON+hg8ZozhhShCoCqMufzbp6qhiUWm4GXEre0vZMznbHp4ezit33z/askjTQU
VBVp+j6rYMcQq0mCkKTt/6f5lakMUspT2jsnG2eYw7XNvKOY3ePGXy5WAFLveG/nNu5g5+vYU5+y
5gc75vAndLO+Qe+JJit9NRCsJob27J+HuHtoE3m2rqnz+c/RNrh4P96Ab/3FRGeacKBTCU/7Eowa
1BvaJzVZ5t9ye6IszVXqoM7dIWybskLyTH2IXv4Ldh5FH8emWjiOCLq/DCj4Ym/LiwfporRSaW0S
b+hmjp2vq+CF6n4tazarTNYlpspQir8dzH5/+DhoPC2FJeOYWEtza5BUckvLVtvMk0gvhpA3qZEN
7krQ07KKrUQbLkUsX3CGMtfPQdSl6srjLrsk5sF4Mh6ZcLqEn40Xv9c7a78erl2AGtyyx6S62eok
uoN5xys0+WlYDarm0YoxXQmd5coBl7TiayU4+kGFX2A1fcK8rfzVywKVlKJeSLoCrAoLfCoYIwEe
3BLra82uj5GU2A+yHita7SC49/pF/2Q8m0rY5YKTeegu+bhUqqBBsuf/EHqQ95RvxhZbNVJ+nLZ5
SD0KzZ1llq7SQ2D8AC09kmDqYyq5t7GQP+3q+8z1qx1Jq74rHEdXJFvsTCGhAQABTmEVArEz9H+O
/PMsnZ0bfg3EjFa9BiCwO8MVOIx9boFkrj5p5OWaM0s1zolS44yG05+ud64eXVlE6XCgaXB1NuqE
0adlmkEXPZYlT3crtzYhNkAPIGDaVqyBKI/g9eEKnZIwssXaYgOvE9euWWBUC0UCioN1HTBJqGpI
D8dUVAW89AANU5NdxliIoMOMV3BSUPIVl9pL3bnY7Icxae8aG9mCwWFMfcQxrPJduMSD9nDtt7Q4
izsR3OW6EnmBAAb33Ph5b8xfC9rRsO7ImPcfR9OhKmAh2V9MQWIT1IfAc4JHJNSTPlocyYZ55l/s
LA0/gVl4WaeGPLx0i23Yca+kwjgD6ntTXV9EkJqHqrLveYoI9FAV8YrCCaKGv9I6IJcT14hUtc5I
gT3ozNMxXkcC4tTvJO9kbdDf+K4JkdP/TtWudIBhVOQLnsAHO4mJ/DHFagVdo/AYYXBhpGsy3yUk
AtJCfZUMWPTO4hwGCNNsv56RmelH5Hi8AqKtgXSLz0J8+OZg6H7XFNaOFrNnw0ANEpoL3hP9z2e0
bC1vWEHnI4asPyJeOZ0uOlOOUry83xAo0adz3+vKuKnKDBgzBAxV7RXJ2hZhdF6eJqeu6sjChyM7
dsE0UmI9Ee6JnwiCn6Tq54Swu3JQyPlb5gnbGqGUyjwmUwe3Hsjj7lB7cFv16MvuhrkZp+leaBQb
5EI9ZALEwsmAqm0LIaQvFDIYUNzkKIbdS62RE7GvBUaeBwFMmblANyg9PpCMk3gFtJAz1VAFlVZ7
VlX4RXCmiGw/tM6gQu7mCK7daayQvA13Q0Due9a5bxA2Bw1nGGkzkAew1cjtQLUPQiPB9JODv/Ow
xu/6ifTvEQ/t1g8F1wFBT542cJ4bdCABqp2rWxCp6JWup7Mmuo7fOSzGCB6wkG0Pms+K73ucJBZS
XE/bnGgrwIbTe8b2eN/gRRzaSu+zqB3stFp/UzOyVsu49b5LEp5/LWHRv9qnV62LxTI4k55Emoh4
rFIXAfZ2Vm8Z7lw6KpMPEL+dF/SdXrB7J54ddAp3tP6xxsLZN9iJThupRMdMmdIKoFR5yyxcqVeu
4yvOQYtR/jvrhrzb7J9dokEljMm6TyNUB7BJl77UMiKY9TnYgVqpzz66I8tROJSJbWZaEAKg4SE/
X+y8Dq1iOgq5D+cYvYkSNA3ZV1hUnpbZdWNs+SXpm2BykyekvZOnllSzglN3jVXyIBi1Lep7Biwc
6uOjqN8goD0yDShU5D5rtoFq/w4XYyHwjKMgBC0PfI4reh58MjcbsOmdf7kP0sNW/XkhFKpZNCia
2OFuDoz6dmW2ayCaalGDhqiapm1iGTX1QCSW3bbZ3FInDQ+mx14PdCdVtpIU7IBIWRfVdweDQtX/
GsiNpKdEX2656pmeQx4PcS/4ioK6b0zH0SnYNJpKbU5o7oyMtc0N9Y4JVzyp9wHzl91e8Vh74fKd
B1FkBeUjtF0jk6TZfI7/X5aOIBPQSCu+zEjBxkJHCxF7eQZ9CwaQ8OteK5nrkk496EgPCOrYRtlD
qbP9FC/GfYNvRGE2XH3uUGtR5HyUQI1fT/J2f+OZ+xKQRi4vrqny6gHP00Cp2fiWncz10FjUq8v5
W9JXRHplpug2tzqxhwU0HWF9H2+cQ7WTkH+Jom2ANwRnXk2n/nda1F2ZWi9Cs+4xrM+Pnj0AT2uX
iSxPxhkVEVwMfi4fhaBkMA7OzPcQL3qxswXV+K7q1mwoaorED7ceshAOhZidLg8kgOi1mykkP2QC
n+iOXPDCemgEi1lZiRx0TiuBVP9PIxUAEly2k/s1SEVBbQ2Q1Btz3VmgvJju8qBuqVuA69Kp41vb
pN4dZQpxs8DGbGafT4o5Yg9Gg7kQbNd8Q25zobDenL+7NmdTTUf7qwkhA0UqVQ2wAwlZT2Aw37jV
IBN0jzVEXu2FBhs7pZwGDO1eQbY/MSQuENQ4TBKHySefMAXRiEACgvahbAKZRoVaMAjSqKO+KJA4
TWqyU9ExhgYyGMAIQbE1NSkmdNEumHxoWWtlRUgwrGSQpN8K/yoc6Souan0DOAnU3WP94CC9+YaF
2Fypn932Sfy6+cbqFsSZLEo35vtJ2ia0qZAPB+SvMWfDJaXuVN6OKmEJ1ZJlXTGQLluYtA+P4FSm
H7PeqpPJLKYrI8Se7MJCSniYym8xpD5U+QjRrp/q6XJ+T39euRxracSWMDA0kUV42Sdvw4Krw2l6
V+9+kFkVa6OkCC/uSXes+i5IGFntGg8ORAoh+PJuT/4zbODFqjQHk7EMDmaHK7YIYoOU47U8/mOt
TcA8Y6EOgQcmylGNB08CYdcn4cFG1gcYoCPTuTypo2BBloupRq5OlBDtw7on61kKPSBeQMnMKG86
5nhIdbV235pv/33QOq96UPwZf2SSR3GHb7A+S8bPHMrVFImeBc/wtUgeKcYYhBloIrnstP24Fj8s
+094UwPHy2bvUsaKnZpmNc+CHliMMjI+roUTpLPHMDXOxaoXz4Z6uClh2UCHbjaUX/Dao76uSqqr
v/nk6rr4VbXHyc7y1VRCKVJhhr5VdqAUcjs2ZBw8tDEg255G4l+qAi9YL7K1S/+PIbLGdB38A0VW
7itDmPhjSFxmZkEE8OYHSlaSjjWadBhpjF3Pq51nwaG1/C6ODzdBEvis2FgCufKQoe3G4hGYJB+B
CxEEQYBkddZI+F3JoT+EC8+7z8ITFkBWCEbzn0oip4H/b4Q1sxia47ltt8Y5cJ4NqWsxeQpUmA3S
LhbzvTa5RUQ7mxAssL3v5/DFYFiSh5bPe/69Kgp59gdDXy1pYBGFycfAXN/cVkAbu+jmvUE/YrjL
oDB94JYgXINADJP7Ux8kTGVVaG+yYj+PmvAIcNDCRHiVkMpt9R4MvlmZ5yOLM5/r2rPtBvMB+k2l
x+MuBN3lyNej+6ZMeqHSfaBtWxw4QyDCGXDNABNPT9cAHYHuGoPGPuIuaJkITeLuN2WCWkF2SlNn
rIIGBsaKB5KZZuVaQ8aBQRqfZTrqn8g7Dk4CyvLgv26ig495mn9i/AG6a7+deSVBwnBSLh4h4WtZ
HpF1DfmDm9MtC42u4t/u3EhX4LUepY6w3PS9nvlv+0oXOhvdt/74BJORakTbIEsWuMYJqp6oXH1+
GL2xeV/WTs4DwSpSDt1iaC1IGxkvYwELQxtZ3G/sAEe/n05+rM8F1wmf59r12//t2UJmxLGGwu7Y
rh6Ur4o51BcsK1ME+DmxSd4/jXkX1qlqdbflX9OmLoHruSrZFaK5gc98OQq0XYjuuy7ze70QFJXN
T0gzavSgHtXuxSzYBKRY3FCnfoo1A7fMRMPQkOi4t4kH0/3287DPAqBhUX4Do6VJzSZApe7uI37y
St7toysIG/OJHJxYKKhutiA4dhEqUGbHCwirZhk7LJ+FPuik0b9ZW/NLlml/YwemSdl3a1Admq+P
hJRf32AtPsNr7/Zt02n/5WYjWPWJOqt/JZnkd4AUPdK1plrMWKU9rH6l8uXhUEtqamxR2c6cP7cm
86gaNZn8MRs0U5+Y+1HV1u7ophfSmB2JOtuMvTrYOh8mhqQZi5q6Gye1jn+5jnfpokMDBUaRNRSq
UUPxknVN2Oe2jTWSUXfwNfDqSB0lgVP3ensAUcIQiCr4G7J+CfAnPwlLa9YozHpUUPJPaETIm6UM
9xtMB1GYcpE7SICQALBzqFupAwacAc2WjaYcoANHRcJ5jldS0Y9p2wJPz2rAULcCHRPoZsL8QA5D
pAZnw3vTHXE1PsxHQk9007Uf5Pn5Efd0UToyWlXgINR1vSgKSNJB0BBU3PPfOuVz9NNtqG82EsaV
0oPTYomqi7NshYxxhQ9TXxShUhej79075t+ADhivp1HDsABkfO/088BGNRJkhcADzTY1lUjCbF4P
XZLlFarzS+sO2pMzHTdCByrdDogIUw5zMXP/ukgl1Ux8AzLCamfOguNe1lMtlLgI92j8rpGc8BvA
ycK4sAX09auKByNDUmaqo0COFqHW32b1k70cIqFF2YE46zrB55MuPBSq1yvjhY+QB0KFNIV3f/A0
aT6mS4pbEuvEcMjUqfCteR20hketwpT6OPL/nXdYpY+uZ1YjinDQZ35JkHOj9BFzM2XdbxOpPCjH
UCBEOZPdMjzS5wGvNV9bvxIoz6J19n5svNpdPQ6fxk5QeCHYw+aFIc8QoKuRrn6+f2w3kOmKch6+
KQHBlCmCP8z0zX8ZWYoTsbky4XfDXaHruHxrvG29tZRdM+Dl4xmgOHOzZjDEAxDgwvx3trBIljUZ
iuE0Sm/sLewQtX+mXtpERCcSMY2xVJYkHMq2nrVK/saUr2JfFzeo57M1E/TBVZh/K30Zw/45fAoB
Kjv5CifVki4X55X18LHcXkkrRaHDvbBiSJNRsCwSdaljCrwbv0Pw8R3nfknITm4giac0ii+8uEEi
9q9stSWWFgTmBCgOYaQcUPU4kRO7cY/QZ4cAYZAH8AYIFJE7lesY8AGRBhqsaCNHOu6tu5HZvRMB
mOmUjxMUWk9eeCYIU7qCd8eWDhbgkPQiEa/npIhX63Q3m+U7Aj6T+S5PPylAuxlGYkBOFkKfBPxr
mD9suBD+xGjgZrumXYQsETyFAb5Y7aVzsZaejbBp4XrzKifdC9b5cGEQtmLA5W8/3DIbUw8A7Pxf
xLx5wcuvXl6QfgxbqEK3TMaWKZ/exs96MOMvVUyTiioLmiJ+eMcD62aLdV1gEHFkYa5P5fnK4Dpa
/LJJV7w+G5M+AxVpNLNePcZTpWbFoYSVJDuB/Tx7dV/kxB8YMkt6HDl+HDiX4OLkRygrrG9t+eI+
ZRk4Fvo7DjPh2ZhaZpVaXTvzINBf2X1eobdcHRbFe0E7/eOnjgeTarsVcU931ROksTKB3+SO3NmQ
L8rDfp1N7OwqrhGxmdu76+593hVe56V6BhubX5qP/aYNY20BcOC/j9SLQbUCI6AYhUVg/U3eKdat
f5hsNEyWH1v+4iAKo/HhaBqN+tILcOLdhXMaMzv06C29JJkKorhRMesLPZ99qLcjH0VftvvO/yOj
M44k+dmHlqgvKSkcydTfv5rpgDCwppklkp7dyROUIrRSlM3BAwftUeV6Q6JJ4E+1PbowKOI664fl
Jdjk3CVnqkrNGxVnSVzJ9RiMgu9qEWAVE8qcTuiVWDiTP/jjn58JKywQMxsXQXBQ03blLrbeWMQf
2x4beMj85u2bZkp6OKcRMpUcXalqegJ5yMVbHQK5mLiFpVYjt9ufnSGSpx9Vp1BdPbRGXAOSj6AY
g3lQqm7b6lD3avXlnHPrFO8uyN3K3UmfXJwhVIfVKILRMRQgIVvJjbfNyTYq2Xj/rMVd3bWR/zks
lfxFKAsYt+xpj3JfhcO2GS4dKmlShRjSfhMmkVQaT5OH8DXy7hWzkJQlGp49DrmUf+i6tP4HYq9l
333nfGDnjNFltbwG4RdHzNC+QZwm5+U6tUC40Xt8Kp8mcSg1+W0yyIQjgpRMRmabF+npEUT15dNG
N41gTY2qugpt62qBeij7OWZhoY0e0WNjPnRkYeIN0QVormn3KSpk8RpxGUW5RE6m7tfj/uI+BdBO
Qte2dW+HXWFyi2ZXXXfdV0KuNIYsqJ6I+vr+21EfnCCEWLp0UMXthNM6LM8ojADALib9dprOoEgr
dmd2zU3Z223rpt8r0cmgHnEKvWKapjI+ncMtUYCCY6beCecZiTKjDN16mHsEO3ACgwEmYL4IkOg3
0b/zdfEpIXyORcHmpifUQvCY+bqFiyd/xv0U6OHyHhWdh1y1hDgj9cUgN6GpqsDxJe/BY7NrFpRc
VNouI4M1kFmParQJBaf9lrvfQPh6728nc91Bgh88/1V1qs1h3fUJ0nsgpEzm21Xg3Ia+5EhQc90u
L9O3NbeiuR461V0VnUPUX82iVzpWGPL2ftWaSpFKbTkXulxqr0B8i+TkZbtU4m+xNdfJZGFAvjWl
KJQEK5urgUpLwMsqlWF5RPC90NOiBs/zwU6g21VmjYKL9eFhTGFS8lNjGTEP8ILeBkbXDv6CarTw
o96BASXNiC+ki2Y7NkA9KD9KgqEMHYitdy/m639PtTL9F92DYhhB+QKzJl0oaWwhHQtn1sUE6zKE
3IdhHAz3sQVH+pFjHqVDydkkyv8wM8ALUqaxHua5ViNyod2Sp941jPOR3dxTtOovjPsu1o8UrGzV
MHKI1A42L0f7ywRz9xdVV9EXhesJvuuKO2We+0FOeHj4PbEZeJvASLpL6tuXS77AuzaUOrN0nLLN
ew+eur8owRLVMPYD7YA913LUJQ8Lu/gbqCeUtvs3Bf7BpcFGE8eVYMbKIOxOYvDWlh278C8Ny6mA
D7zLeHR6QfTYLyKH/X8LwjdUzxQLL/zLxLxnErCIhQ9aQFkNo/ByD2iaaQeKDygVZzDW+X/lFnUf
a614yncZVk7DkJGMoq8p97MNtm2qn+CA8W09eEjTFZEU6ujbkONBC6KdWxJoUVYPDip+a8qGnOeM
olOuXJ9YH8Uy+P27LMQ7E7fJXGnyFxJsnXPrkzIuyRSQQXQafUNiX+p3eA0uV1VSNtpoflu/FTiz
vL47/6qy1r1JFV3X4rhbhxaE+GKNi2+k8nT+JFUtCh2Ova2t5QEzhyMsZ4bef6e2zzmNNWpL5DX9
DZur34flc6zo3UbWChGxUqtPd/F3Gw6hnNvw2nh9s3ETpGYB3rLDopfI9sGes4T8/UJP6uc6P0Iy
ZdmKEOQzvuffvvL9AK0Pd9junrKPF0IZ8bDIsQykTNFLlH+mbgGdg+pnXQFF5YASPDVw5pD0z4H+
D0yp03QYvuaIneS+th0LS3UpSKN3nTxMXQ98xhupis63L5+aYuBjjZhqMv/jFiQMnKEs/gHubi+C
s7/ALF9qI4VY2xrxkNfoFtzvApLK2CoF9dYTK3vzmVH09a49uTmRwSjezPz6O5hLGjN1jEWsOF4T
q5RPVx8kVd3XQLEeEiGbSDsozWiDnjm6K592AIRCq+zmon3P/YH2V05Jp9hFWDjtb4WS7UNmo6t6
56OLzwe/8yQbKVkOQ8GurNl7nUK+oLU2bxx8SgU3EvCj/sMBMlNUd/6FyHLF6hp5Q0PR1F5qb5QM
ezQcyNFw6UM11MJCmreJDY1DId7Lg619ldXArTZYEH1VqlQZ3hHSSRR5xqgmggMs6af9mmLmZGWK
Yv91wCNBDU6Aa57mznz2q2IYCuL9eMGaIwFKlLLX9fjZAXqF1CZHNxGi41RvUhQv/UeOq4Ax4dDg
oCsVOLMUPWstt5ML9HXWJFuQm9BXJjV1tyBAcvxrdLo/PifRhqaoKWtkhE06y6f6Opkwt86zqQLG
UTYz9zZRsHFzEd3027d1xlAEZdjFfx+cr9gFguxJvisM8D5m0fJdt5Do4XWeJVcNLumZRtJbx3U0
na34TiZKjk6+3IKkdcAuYaByfAPoqV+cTppXTQNdrpduXc0emRZS9SCq9dIIHCua5o1k4YU8iZtn
f4vILHnpXrKzUIqSwa1QiCvbroBKH2pWr2PbU1QAz8HGNGg0vvK/x9dljfEXUsZRNxp3aeEOmpHN
nBImCOlKiz+BdLtQxElfghP0bQpp3jGxkkYAWEbavTHsfYk1zAKCBuCt/I0ZMDaNJIJvWlqEKRpc
nS37GlmZ/AIaP5mGrPzF3jsjYbODxxuMgG5Ck8SjdggetLSOo5AAd19/VngLUcsYELZu0hvau/U9
aUQVKiFX38iYPdkHwkuiClYNvbZR/vw1KkAtCKrqE5aRWiYbcboWSajgtRuXYJvwrfhiNBi19Tzh
OwGhYQ+sGRmg2IUFTBIvkVfkTtZB84xi8R+iF2i3+6y3hXJ/LT1BaE6uDqtpvWoK8JXn25wNZcSj
JSzBZcfSxBsykb2uHmO5+4F58R/p8Sk42yGR6OFrFhEsQ3gPJDu7tK5EDc5HnTP4eH836glQsDYW
Q11zSnvgoScLWG35HQacSy69aKuETGNILeUNPeii7vxlJVQEkhKP16sI1q3SHXyE7lkPxsBgvUAD
COoTXyIcTnF5WT9LJGyCO19JCfMJ3fgVklGUUhRJyk8oIi6jllETRLiz/zFniCkEmaQWor1Kf6G5
Naxg/7eLNNNQNlcYxqzt1XwD0fE8sbag6uj0x2npfQFTFBOhSl8coBZkMKRoblQ69zzC+oMZCHr5
pPR8M5AyK/Hn/ZqeOimafCkCFXUITV+y1C/WvnquOiuVcP5hJq8p1pKhehb3Hvnetufrt5NWYyzH
2Og7soNR+PBa4Re+TTefSfLrxTPKwHdizzoGRORiwsoiTg2YDfho2T5i1sI7wQJTDtXkynEJ/3IK
DOaQzBuFWOR+kDiYeGS7PQ/bQtDjp7rG8jYH1Vws666hnOseiB5Ii9OR1iJ6jxwx21OCZk2R4wO5
q8TOrp0ciH3zGLJbm8jpVKTwWkUEPVrIJmv9Rw2WZ8mmNR4b6te6lFHlHRD+8cdD4/ZnqfEKvokv
TmdeXYCsc2s2PI3zS+vA5U8PDl39Hj9GKh1mxoO31YW8r26S2NWkMkHlZsBrQnIj+ulnxNpbJzPq
9Svqb6nNF4IzrP07KSkSN9l1B8NZjvSI3GnKaXmT/e1sXyLr5kZJKCtjFAzOz30HmySRpngGXELr
OZy/ZGUvQvdrBHxcjz4FPvrtj+RByl2AYpJamL6vJJVb5xud7hO0rw14H7oZM7IbzoN9m4QFYNXC
B/knO8cxXtoY7nt95GTpUVQKHLrs7nLXVDOiLEkQp7H2agtkwK1mh1X3EAxbqc7bLTJ3+ytQHewJ
pAT9stT799IOaOW4ypiJQ1yFw2TPy3XcyR5GVRK64NwWZA6rRSkSazVfg8HvmlQHBz2AmzOvW12B
zm5Lz7B1tk81Kc98n6WsFf/Sc5AiOjRNJdpgsprUZvru2GUBmEcjiFsMb5QwRI8OaULYSE6kntgj
et8kJPAZ//U8IraM6FoEzaYvcTkMGUOqTBfniubeZ6VLY1YmgS0HJ3W5pqR3oneZv2Lj0zYmpert
nnUyyKZZMVSkbzwXQI+mBoPViw4cwbm2B3zOLfAxXOLbgmdR83HLrBnLOF5TnYTnzkb5WLsmK3cS
DCt7G4xhHshGnynRvqofeg9nrZ7cX0iTTvuKH5ZJHy1ju6G4eChenUrdGY2av4qKwWgfSo4/XK9a
9ZTxFQ1qgPXpKH41ZRtvP6FV2i20NjUHNJcRvf/LReegvjYqhLnulmpkxBquNgIs4uDGe3VLTo6R
TJ4tjyJZJKAJOE/i4vyHrwVx9Cw/asO3ySvfvb8/N+sHLwCblVUNxtUJBH5Y4HlCs1jdgqGlJKRR
sm3gsMtXZp9KbkgsDIr+Jy1e6fzF1kjJdX411SLyXbgAFlWUjAiFmbaToqt4/PpZcTamc87CDlAx
iCbFd198mU0C0L/fotgbNZXojnYnJOZz8mRSnZIarptmAYqE/XOzPk6efD3n9LTV+S0N1NiLPC6E
sjzSz0i5TwCdzvabeeuPMghoVZTk6EGhQ+/bFAHN262xYu0WkFMHy3lAaFEE0A258cJuoxmcZFKj
v+/ofbJmhAi/ow25D9MF8ugc8MlncCElXDIgCee5Gl0Fnrt7StjbDC/mG8D3aGK0U9QP1HytGG/X
nMUjRicC/fj8OACp4Uc74udWM8JEHMs8SewHW10dvbzRSa96bPdEa3zcGhWq5FXLtbtTHoL6xIn4
MHG2lcV1Gfm8zNekvtTbZk1gJdmF5XVdf9iWGKyhRHMXWBDKBP2BjHGWOqENR7BJg1S2A6D1nGFq
N/QXOBrGtbKxwt/tr+9jx1+iq+u0+fDe9YkzRHH6khRkznguSWNKMyzHWf0FxT65BELfZKt+qcjI
vQHUCLCFR+/mgIORErPmsw6waSyn7lQXUfI6yuq83KKxYL83eY5U8RVTWqGyD7y7UiAw2A4M4ID0
0MCJFW3B15/eBXQfXlL7wEy29gelScr7KNVbS/Wiag+XE/bUBJgPAcq/bCuthJaCs2TCFtUn8Syc
C8ECksSxzPjAGT15FurVDaN10PaPn4ye3NaLfZ1WYczvqs6qLgadMRCAmX3bLn//1wLtOlMhh2Nn
nnGWl6A/dZIVpXTQqHXx7yNqCoItXi9WSEbT2CnxL/uUjNFL6NJ4fDqIvSZeCtaiV96OSEsgzbJ6
HT/V+ssjQNXDE/Pc7MMP/zjtYosz6F3fHqGxwIku12eWrYvpmVCN1+0cqvmeDV+T+aZHxebZE+PV
TksBcLVS8aZlIsHnNFXuSXBM3d05RDRi8TLnqmPrF88j/PlrEIXRW5u9816GkIEXSAPWnOQkl/sd
1iH2MtQNroc45rS3QmlgZ6wYY1YkGPi7+83hR8XdKrezMh8ytqtZ0t+ta6k1gLc6eczXu1FHdT26
GnpGxjwjJlwACDwgO/Ect03qqBmbQTXYvC7uNqoNUc9WpAS7ke+d4LjEheTpbbweMJxK9166Otmb
ToCuUtG5qNnfPIb8Nd6urfWLGMFH7Q8BDIPJqGKU6epgVnIz9uHvRBNasNNttSfXWE6ZymPzAQDn
qKxSlqqvfY5/LF9ea33jDfoy8Iw33+9vspKHX6SNv+/hRutyEJ4cP3tN4CBfFZ7uGgIQjEP/KVx1
ooplVxjDScMd2mQXwYq2AYBfNWkKsT/o49+e5qioCoeGhQAwoq176x1bOIjgcdA/0t9AoahgVcPM
aFaCUKF4M3t7msL/q+k7p6xSQUhPzF9j+yQD9bjy8aev7Xum4XcGrPAN3LILBgyNEinJT7kC3vt+
X2BGoULty2vDVWBLJS+EJJnEptReDC8jd2TLpZY7Nb7V9ukaG4EHRGUPUgfNT8AWwX4wejj1S31H
xqgyI0flyk968ZTZ63xkvouwqymF5nalozCw+zwhEM20eLzuJi0jMpL7v9lLEgt0DsVq+NKViTUB
iXSlHLYZvcDWFP6jfzJOJe97+vXeJrIv78N/Vv2wdqDsaUtjeaQwt3A2u101RKA+SBm+xRW60vId
46/qF4JJ70f8cQsVXIDZ9XwIMqzrh5t3boF4/YponJmyVIvig1J+hRkC0Ff20Lc92egscfzRdmmm
D9uFzKk2ELcTJncdpX279XEO5nUrEl+DeG+xxsuaxdu8qAeGpOrxk8qumSa258w2uHZ32ZF1gtAE
TkztKmn1awi9F4QpwqCb7PDWQAqdQZePQenn/1Tiz6d3H+KM06dmjStF2ycQta6iRuD0faJ4kXH9
RJj5goG0VXdDEt2IZanvABAuZZba8urkkZkWQqRX7OPyardnrsK24kprgIGlLVJa8Pm3Nbldt0JV
x0I3KDZSr5E3L3Om2lpFsaUWM03JRy7Tl2vWukEEQPtUGN7OMbcvM82hrftdVyeg2t/UfAljekj6
qQdBpyrIk71a+RSnZr+bHKdj0aHHmatXkU3YV4q2fLU40C/8yD/zGF/3Gofu6h5R47DYlVNtrat7
z5SYaE0/c7/VZe2fWzdCUfRtntC6Qmw9G/iCw3CgyDruPbtXdVRRsvLmh7CHF40DaJcD5u80li3i
/TWs7olJXoyHxRcGWFr3VQkCsyZMzTBWOo7NSrbfibjegqC8IjBet/jjDHm09O39+u2A4ndw5zyB
m8kbVvXGgsvtDywcCM1Nl80jyKzaPIXx40MhCMdy1CgCPwP9vYgHn81QHojQRLQIU4AUvKpEwYsj
uz9A8On86REeDDr5CA2BE6w5tsTAr8a0jVQMqEOgERO5WO5XoCQrGRonkytsxpIGPgYMY6anQv53
tYJwlLwY6KVSpcXtJC4U5oDmpx3oEgCYg52aX3p97SGlL5nE4Jvnks8BTr2e0v5QaOwhE6C4R8IQ
cLkbLfQEwPf2463LsmNV7/gsoHgxFstOI8X/HzfJyanfMmuwRDLZYR1MWmytQJxvPDVnC3EyMliw
5DJFRvB0deW4fjJmTOgKx1vOfYBvdIJn49emjC9U3GyQ0GiiTdE+iNXgz3CC1Eoqq/CIA7uGiHwW
QKuX938hv1Q64eVNyfRq7Pv2bUhZ9/RFjgLCH/0XJu1W2IxLlQd66wWgV1Ei88fdreS1k/CqZthE
wuOECWbDC7iBr4zYjb8UWD9rwUHGnWYpJA/1sr5R/9s7bfdUpV9+zqB59/I5PQ3IPs9QZygM4t/J
j4q8dPvNNPXh9SiDRn7z7mP9a71T8Pt0ClbWDoT3yWymrdqPp0lEGyaMRN4aBGUovSmBuqFIyVzu
L4hTtaLpa/xyI/xZlmLX5lbJtz1N0evYoP4157Nn2JZ6fksIxl8IyF+rdID9IT5xESEejVUasbaH
yV0NzTQUB+ujHJoRE6u0ERMUR+cwXFs5QHbhZfTmQmH7UG+OZOdkYl2XCFOG0lwINNNbVNJ9EmaQ
haS9iSi/xAueX8r3JEA0XubRaH/m6BcCXFU9gekSyCx64ICp2KGcfzB2cdr4Qay0+/FHJv3Dt43M
yKlXWaKL8cUT+jCz7Xm92keFCiGgRv4JaSGdq7pLVBzuEJOmfZr5Xm338phuCvJs9kV5uu6ZYuT1
aNF36DeoGvAYNhDbdWIWExUqP2u1FrH6W1L7hws+P4gIoggF+IjUk//UxUPymvwiA2CYDBBAGHLS
XgukTh7vkfVa8fs+8rNEiUSVuXuXmqWZW0JEIrGzLt7W/g8MRpYvJID8S8Kh/S4NhXIkudTQLwCZ
QKbyNB1Gtn9B2wUC52FzXGxviQDMA9ut5QpeY/U0jT/SSxHLwOlG07XD1suWnquz3gAul1xCYnTf
i7ty8z6nPF6HYyMYu1sk6NSKXyOrK6BLjVuSAooJNcPAUa9DjUP1NDHArEx1Dz3oMhmp/w7UWS3l
9ar9TR7Sm07hCGmFWxYGTfPDanKWD2iya/zrAZx7HZnHvcZn8WHR2D+5Qe31HaQYk1Va0K6Fv5li
oibvuKwtLrrD3Y7gIsEAR0BCKfzCuPumNmrtd4huxGgpIabpqHZDYVA1lWjAIKJkOvxlSs1z1lTx
TOh81K1nbRm7VH7PuVfT500znQdWg5cCF4g83JB+OKd4CZ8k0dQaePZJ3DNP94AWzbVDpz+8B/0b
qq3Y9dvXDjDjpHrEp537AtWeQnS77HJsD5wspl/cbCcAZcpoku48l7fEiePD4fI+3CBmT5NeveRW
usFHjuxOghTl5KsrkNaMjZXiwa4gomZn3sQXQXBnsCJU+UfsBRdngaHKAiNDvNPai/wE7qNXcg6F
smOs0YrVLl0tHlk072uLDqvaiEyB3yd+PkOPrX7ubBDkc0hUIxxtMxFf6Um73VW/sCHuzrzWwKKx
hSgMbyLAMf8Fyp4ddj1xSeRhek6wxeianpcCjUsBoo/HN1c6+cShGKCImgqTR3sZm+kW9GLYplNR
q3x/otNkRTLc8Jtp0AgpEin//VmIaWHMwO2tdA+lCYPtjIeoGdgi+WDhaKVIBjJtGxevaV3uleXz
Czd8l+PEf/wAAii6+NuT7XDAOCsE1eiXtEgNrC39tKNpkJI+IWC2j6FT6pidwEWZ0oU5N8DRkGfX
ICQNge01HiRTExobvqYs0HYU6mBGmlZQ3mRIInNQ6JG7aqF+0eHioMQFYXt8PJ3aIcEN0RXsGsGw
MrJvQYxIAieyQ2ztnUAY8PmUCXtk2mVYK8kXKbg4TXrf26tb9hBBr1K0qOW28nlzoMwF61OmPCJd
nNAstxuJtLxfhsm4/xhxqc6KWG9aUr9UeOYqr0QHS+YL243U1I5LTw/x1hG8hmc3Kgo0KwFNZ1Hc
1QxaovBbEUTYqg7SgyyPlwEhY0QfVPvOuhNRwRoXUztDAV4MTn5EtdAgeUdtNLDxAPQ1o7u6AbGd
6UWVx9khdLtDmJYwf3lClBIzPAJhDN0iRX+LYcg+rN97LsZSl8Z613VwQ/B1ylGiJ1LI1DnMiMP7
tknePt62/NFedKgXI2FVSjxKth6uKKpRJhYobqGkw85MbN67QEmjgL88QQve9mB+GxB+wYPAYJiz
i9UsjDnO94hzdO5U2V9nZ4K+rzlvlkvIwlJs3o8cqTewJCRlKMXx30d7sfZIgf6mPZO8AJ+G0Wwz
Pg6nd7uNZKGFtQckNXEPlPdzttUFmUuPCU2MhiRpl0hoIXyfDmYqJ+zbVaFmXRbtFb9WPGuSQehH
blif782wTmN/C3FQa0+r676iD4BMmmkizGX1pVVU+pBvTJGo8exHaOA2PsBSbRZlk/TLvFdm12mS
H6MQWlkZpX1EfrYd+z3m2zjIT7iDCL+5MhyYw3QKF5now3osj3WNRw2yTmPJxWKMky75w8sQSA7h
uluzj+5gxRShSr+E35KoEU4keZ4UdD6y3QQ2uuazhaC1sUANIezRj4NDk8lQp3R1wZ1SAWM6kHRd
nFHIc5VBLiypF0UjG/Mpi97F0DCsgx74W7fEJp+27ozh5IFMUnIa8fRxkT55lbnecbqNeJr9YeX5
6ggM/wsW7Do7366ph3jSCXIYdDuJXhTAaSbpripYLnbnc6nTkcFFJp4E74VRntfqB304ENsGv3DG
Xhi9PhqWSc3HeH96rJ4Gx3yjl9rL9jvbAQLIs53hjuLCGs684csPpu0uyctvvmFT0TTXBLAhmTrJ
aFua5tTpnM9ZMfO+/bCsYIKqmmj2CvFWiiVlxdnMKe3RgTuZNWYZQTUyDH9djo370ZrsPDDQyUYm
/On3gQAPzHRG/4/5dCObJuZVMs5I+rBw98NgW+L0AvPfcTUuyq5CF2LMaK+YjJJZHE7xA3Hdm1i6
wC4ejR6DAJSvByD99LIfvKb1jJmVyNy2EtZ6KALOOuGsyWRXF+8yUh5Q+zZg/wKpQtl/hTVb03GI
VhU84beLpNUShDITCJFIJ19KfBiDEQk7bSkHrnjncgYYXb5afI6hqNLOJVhhK7Qhd3ro5m6ZnQ5Z
BELpvkgLR7cXAv+tdhpl8hazxc9vUzyT5auRZaw+0zZjWEOUZovEsuK+FwlHBT8VEYfbbvnz3tV4
R+m7Pj3dPLz5+EdeS+HvfrtWr3pxrvistRS5v+FrQibssEX01ZobLpvISSHNOjo2YjjERlhSkeZ+
BwdinQt19m5/i3UrBOAw5stDSwb4Rgakc6ohsOxJN0YTzEZgA8eYkvTTn5tw55Md5VpT38Kv8vEc
uCzXYjmRA7aMm6AQXvzAjlvtVj/cKx40ErTyi0+NUBOK+uzVGM1cvmLFOSSw5NoSeFH2G+txCiCO
d9FtwTs+kfzCYT9YdQfOBCD0ZjbWuk+76zCfC+mbu/aIOPFrirlhGJg9/pjdW0apqSPLu3HtI3BS
+Z7UKtR3TFk/Va4qWp+YyKz0m6YMCtIqeMo7lwd/TixyL1D5INQ7mtcwmyR3aREY6fumTs7Lgh4t
7QQolSj57D/tKf13QMmoVX9mnu8AhKQiB5lFmGsO83k3qHhRXHVI+whk+9hEW/UwtU3cm3MxI/gy
qN/JXHygjMZ62DV1ViIvrvb2xvzD5afWvUteKcWbjuiLE+HnP3b2zswvK61rJ4ehskJJufz6zVUI
bDUmMtk9q5J71bx3JholD8HeQR5mLaKfpzHSyxDtkV5+qdT2J4SnuRAR3NXvDWg9flhtrowhduld
M2oVUezdnADRsx45HCg+XhDJ9YTyBU22VHDfqGi32cALQs9lR7X7vd6qKtBzDj+temgRqYQeTW/B
o0gVcI1IGVFGg7tdXSxW86MEZMsH9nz1FXw8ftIMKiasLW1MfXR9rPjMmgfRLJJh7tXTET3pq6ZT
IWYn32JFiV6NNTpx9GpRr0x1aPDCfNeMflOkFJtO8nrviejSyMg+k+uLcOJPcJCC3XXPBvobf4V/
Au82IlRVQGp3Zq4vW1/o3HhfiY1tKrt7F8MTostINSSyEMPmYFxoooCwJBGsV98UyAHyEvwWcMS2
c1mea7pGoMKUdBcFHgIEFW+QGxjSCEmy2JKh7NBRBdF6Q9RA4vhAGiURKwa0FnjrNNu+n/ZA6CFD
D+huf8r2oeWvn3R+Jy+EPEKMm+bgqnV4ESFcCdJ5Vt/zt9nmyfgsaKBVzpja8FmwUtyR67FnOVo2
680yMnEgaXIPPh4Jh7gX2xYq8Hhxdx/oU5RR8FOGADR3t8fLgQncsnN3j0QQ67y7L5NA08PYQzV8
vH0rq5sfdgtW/3q+bEy1rr8MO8qxbvMQ/A0lYHcsHBY9RM1Cgof7ysRrrlBk+GDkiTe2Zslpq2L0
JcSjIUgWoy7gQNor9jtrABR5LQggGeJYWEbDOZN002G/ZThxmRM3bsyUn7wylFDTToc8Ii7H6vwi
ukf84eRYgea3AdVCunQXyP92k8UT/BZFZ/FubVdKKEBCUn0F6NxM0dB1l66Sjk9GlT3sQsC5gUa1
UIJ1qBh3tnpi3dNLyJJ16Gu5Rt9ugLcVAP2N14+O6knJYJ5OMvkZgOWsilSwgxdxBmNkHRUgiTBg
a0gyPDXp0DbziehFul6r0FyID6wfgV/XkQ7AapgAV5yx+Lu7EVGkC2sY8R3yekvGIw6rk9hC2FNS
/RvZPgDzOn8VZ9h3kYkuk+03U+nAghbpyCelL8DCvPuAlyxnBZDheQ2In0b6G5nbVjRarSydcTYp
dcLmBkRJGqPxz81sCeh37PHKw5jpci5+SQCUHME2d7eElMG1EQTL4sUyRr4GDQdlGbtHSWExU+4g
rg7KDJ1ktR4ur3oC3uQcmyLTxZrDabXMpBAcDuW+N+QDL+n/1aRPQOzF1zOerYpPF4yeBNq6OGxq
zY7wRYdHUpK0jvnD6p6OwHpK0o5SlyEpeI/szCTD+lntLLmId/pGJ5wijMnGl//TxuK2Hcru0Nus
JRUktB/bLHm3jO+xJMIMP3/Lh3VIMaa9jXwO3dgdWht4rItL0TzBCyvVh5HLRZJK9Pu9kJE/nK0j
l2V4dgTwXl0NYTjMzDsqbDe58s5HQSQwV7P7P1p1sjnwImVHtwr+smzJnqnE55LKZnyhyxmgHAJM
Fi/Lc2jkxvZAS3Zj54/S9yvwgKruFDRwyso/lpTiVjv67Gtk91Ts7iKUDaa7saTWR5lhvsHxlk+Q
vRD5B0AC7y2dGjWtBLl7cViu+/m/5+8fY9rUKgT62+4+HtARhHY9NyqTkY54+o/NABgsbqFMhYcK
Nl2TVSG3LjOqOtPmYDq8tNfaToCf0yzPUeoYHxfsoBnjz+NYu5Zu5Z/jyneB/2V81URnEn4kudJb
f21G2mkE2fc5WRW09/W7pKw79aj8GF1NiHlERjp/M5NJkN3rO7l038/wkMzEpu0ZtooWl5CSMdNh
qzLNUA+SkmovQ7B/t3jx3/Ov2XT7u+olC1KxFoSGCl2UQ3aTdZL+aKsaZU9KzJVZ+2CzF+wTuIQU
wSwU1eyPy75SKsy7rOduG/ebZPd1bEbOrF7h4JCUVoseeVOHfSlTa6oB7jEnYAREeOZDRKFoaQjm
U85L+8KDd9CwLZQtFW+G1PQL+6+Hoo78eOBkgfW2zeSy1zwLyudVDrMHUWJPYKMacV5wFK7+cV5L
n1TRy3wFy7b+FLwDXx3K9VuHn1VdMimpuWOB+GctEdbPDnX9uTP0Sw2f+E6b8wlvL8gDryytPIRI
IxErKzJkEWXVrd9nnAJiGprCD1euydnHD4Nd8jkGDBd0B74DCQEMJ0SbDubNdcvfBpBWHNFuzgRW
bTyzBUpwrWOLeXw7l+Jj0ntGXmTKxilhlIzwCrhDqnwtm7o3BQlMITQ0p83jMp1fdhnrXFUS2fr9
sGVpSCrcfjCrh7brV0mVqdV7ni5cfzAxBzLNO2QTOHQtRwX4mUvLcRB5Za89LWqQ0BWaUV9r0Ykm
IO6AZte1Zsm5QMxNOwKw5CcPSbs5SZWterUWiV4JgYMPo930e17D10z8ieTjL5LckE2ugcKwdSZ6
z4/qFpiatf9YUBOqbl3in6eQ62ddzmbXQPb3ZcwsHy0hYerfHjEV8Q0qIRMPFqU8S7LlIAXKjemY
2iYH2z+fHzjEahOeTGsu44fMTYtCvFJcvd3bnw0uZ5th5U0duf0P5QMN+COryiXnYCPNm8Plpp1m
GA7d1FnqWshqV0Y7yHa72XQqcY/JfKwqsiyoQT/qerzI0X6Ong+H6WVACCGexs8V/DVWVkv/L/BU
mDC0a9fGpGmYgLWlmT3Nr3Ari1Lb52BtrR4ec4ntYvs3eVl54u8BS0682u1mKhXzY0ng/XxABA61
Wp7uumIjW2g2bVw+db0txz6zVf0mzOAHpDZvI9tPN0GWwLeJf1SiZJLlXg5fac0gew9e6q5U4Rhk
9pelTDaijvAxuw3+6T3HZeDooo97igQV76UvpJBfZjqzx+uxZn+nyDWLmPOy8/4QWRAfOhc7XsDZ
rE8mYOr/Kt/rUyfwaFXucxFRBXI7K6AU8b8Vwn1GyZ2OIwZXn87+LWR5cNEB8N/dU7Lh6eqWPqy3
fOlypdU0AZyuPFVdsn8YWWpuhiXSup5aeA6nm5Q9orxzRR8zjMcpRkap4aSTD6NcoYt7aHW6Ia8D
r0Iled0jELLE+j+ia+ResTv+k4rPVBStAQqm6SMEAf9Xh9+aGGbdX5y2t53Rqy51fJJ2mtteWGOc
ZY+NI6pf9/jcxeyvvFWX/j+S/O6dzFJzxhEDdBuMmxwr0P9G62U0naqS+U5OcJ8SiCZ1vNhP4UNl
543fwHDWEBjueRXxAjKNaBvyyAPxfCoin90rLJHCmgMwV24UJpikmZykqngAZ6cHvwSpOYrBAlGz
7xoMixAHGMaEANqrWvS2U2dJH09F617TdgAe3TMtiwBQALL535TvaEqWVVwqVQRMUtMF7mx7YrZd
lh4kN3RRFiZDCeuL6uaclBdcql0cq3oFNjbykaOE0Sie3WLs9YdeOBz+XhUQmBHHVjnENBQAo24+
MjvkyfubyRsnS3L7xB7BYThLfrPBVrv5/RbSuKEyRsR2XJ6YdJvQxVG9hv9H5OSiad1Jx22NacR8
J+GwSnlFWt3I+ocXR6q4XVdQM4qwt+XG+hVGKWhNlQHimwDQ0AftlPnUM3dBNDSnMtMf1GDViHHw
ki0PW58w0MIcpcLd3T2LYV98diWlFEQcqrAJg1vAVc0QxXmtvqTmRo4Dm+AShCns91weTNnZQyxz
ztUCwZrzhtm/djbnxDD9cpCA/DImWHzDWQ21O1vI9pVkTIQej7HwBZq+CaqWdZRkv39NZxwUUHKJ
mkxnIUzGYVhfui22gW0LP9HBdiUJzedb67ZiwsRgIFWYAq9np7JcDPuld211EjVjgtV9kj7q9epb
SpcYGQoFmCCSMf9rT0ebfNI3gHZTb2+JM45YAzu4QdDftSlizuloeLmnxRDq/8wYrztkJu7e8yD0
lYhWBDKv0PHkWG3OVGq2P9eZFNqumow3Idj3azwDj0ExoqlXNjHug8CvmpPQZkONmTCLgIYxV7Mu
0O6+nAX8TFqRu4LkVtGo3HJF6dPNvH9qK+s1+IX/jJzBAUr+dkXVwJBZqLPhP7yrYiITSA5mdKbI
m/QFAgemYU1I2Rk6k/8T6n2iVPdnTYSyVlSXkaxsup71YBh+ftzSlz4EiVl3H5bMCR9ujct94822
WTIb56Pc+vn9M9Yy7pqKhhHnyChvoyXHD146/CEa1sbN3WGxJQC6NmlK17LjgCfG+hYvM7nVrWTd
m87faqehkWjTPheoFEM7bvb+MXnKsVPwRaLZTLSeL3/dD0tKXt9N52Zx5Oe+SkkFsQBzsEFadLLV
4UgHum/WWTeQlSn16DXAbBEFPlJ5CLZYlX3i7LLyp/BRdq4zzGoygo3JAJdgBXSDnFz6gCJ91yGR
mtfMMx+HGpTCxElnLdHjsnLxjRxw5huIFriXbFCz9Azu8g38hVU5prhoMr13eVQHv/IQzB09T6VH
StREZcrMI24Od9AsYUpD6pLEYU8IZ+ll8KnA5uerH9QBc6vGVu0kqnsDh/wvuKWQUVslwPNh/C/X
8aCHN8JlOWVhfX86Zx8Gig7mfA1+w8lsEwhen6Hz1ZkXWA6nxXGbGK9OKuV1XsviMKBkR4BgBcSk
6OoQMPbaIyh8IN+a1bkBcul4KD44Ru78G/8piPMduEkzKPOWvePRZYqytfkCmjp6vNdbOHt/ImdX
DZmELcQQclmAqrAdPyMyIL+Oq+skVCZIG+0yRBuIxOMmIAdJ3tDeJHpspqlfEDuhIZQsTv9OhjID
0UGgEyTyIcow5BSAR1YTZCvorxwoguyXEl1llwcjgsJOKgI8nnHVEzY0hvpqPKwXQRe/MiV3dqZp
grq8TJ5USiHJoAdGICMV2plDYKnv5/liJHbrz06sOr4J4Y7ANWcrcaP8u6LK+QWVpBzZ2r5jx9wc
yn7WrsCG2UvTXknnwJPv7wXHZhXS3kuCSxEWAjp3QxA2JJyeQDwzxBPAUb049nDBRSIP40ptT9mU
OVQueAIbFPj+uWnfvBi9eh0RaEAKoCltxFEEalQSZmsxH0XDQyfMkHKG/rPZhwTAcBLLYEG+mOiQ
1mqPxeGp1uwEKRUisST/VxSgvMGOUqDTZiarZWpKI36LdxIEdP2444uJZfKMIu9WDwLELc3Vd0h7
WS5H8v4emB27MYCrpCG+Hjtjhj3QNs7/kafFe8qcIBN/e3EpT7CYzRhb7sywaOiNS7781WhtKsyV
rJdoKMXVbztb/4bbGAIToU+IOxhwvTvUqxegy1K80vio4rz1szYqLkipLOwhGSKQIuE4JeZOE29C
pXCi5xcXlh51cwehUVIbXvljTWgumDH/BWPPJNF39G83cejy1eB715zuVKbEr1tWLG3P23BUPUOQ
Zl8UURQqbiHi3hqeAy25zEDSeHVANSY5u+gIXlnmD0LwlR3k4zY6ECqwi7p7JSnjHrmdXteqdzfw
dk7pDbHdyc+HM2/CMA4BBmNcTX82IQlmrgaYecJbtFUXw4j+uPZonEtFSEYhbZ9KmxrWdKW1oIxN
cirCsqO04WRpmusM+BT6eiQFm31EgXUcc9tPJ4OnJteT2jXyloKRp5zE2t35OEEIuCjHibP1li1p
WaU5Td8Sqs9rCQH8mu/zkpdgY3ZVrfqOS3oWM2Cwec+jV8KiK2FTUhGhAS3Xl0W3jbznpiFHPTz4
zONoMoLHVnYX7K15C6T8x402FEIbUVRUxKH1tnZnQXWvdZ/OZGp5vbuAWteATjmNWY4UciOEI1Ny
9pee0VlHZ0F2GPnqgAe4l46gwpIvepafDGzcoylHxD50ZvXF1YOQF6jgtaj7D+JX9iOf7GXdp/OZ
m725NspaFofKmwP/0cVjKhEBO65LgAYqWOzLyqg0eK7iE/azT79YXhAyVfI8xg2QeqJIOlS7umld
7fVCpJvCkmJwm0ELO4GCX9dYF31MobGWdaMpmejEtRrZWdI0YRT+JI+xBcpcLJnVDrzMFnWhjiA4
zN4lvkJDxJ8iV/Qxltt0xBflLPSv1yAsz/mVpCaVxQ4tBWd0XeaUROHvri+GIZWYJxua9eJKFjRy
0j6bOisAxr+ubgwBnYvVB3mNHCjayfNFcQSXldlDAGmeAf02ulRA4qlFKWmSCxGuLd3u8R/VaPRE
dkS/FgvxnpZgPftmS07RRm4yE0lZCPNXAQjkmaL2kpUrAxjiePeQUXXxuNpxq5IDTThagjkMujTQ
nObCjHG5drbdPU2Hzgm7FaZK8KS2ol/9EZE51Rayr6qr3ufzjvqcwtgNqRADAT5Jw8/ttiO5l0kv
yEabPTWvDDo2N3jZh9z5AO8H6AZzuSCyCIvZgg2HMcGsFf+DIw99I1Oy6DvyJutQLreUpiqbfRQ6
VMEiRn/w4Y7rDU7zi8QrE+SX5t+F06b/zeYXoSEspNj6ManmQHL7zBs85mP9uW8CEEBfdnqin0Fq
m+9tdUDiWZ1cEPxfmZnM+QQDmCiUjanFxj6sttT3B+1moh2TsII55Ft/6+DzoVtzHgxRGfdTabPR
Sk5PDJSrpXb8KiLqXMtqEdbtnHcAPTNweSeSVo145cRZFmJsQ2U7Uzf/PynD2cQEeRfPmghAnQ+d
I30vpNq0Hp4oIpEwqiMD71TDg1ZbF7IUtd6JLpa1haVtLNj+IoB1h8fa76bla8f2ClSRoyQRXgLa
z9YRgKHME+czHAGmQJ1EBktFR78ZBWo7ErkLaiolf68YQbuVi9RTxoN/wkjJUk+D9K3gkm+OX8et
M8lyRgSNp+Wj4JUTwgCX0OH27xucHXnlta2V8PNdZSGSAKS7HqC1e1N2TGiapO6B6ln0wMDWxyjR
52DOMDOny35FFtNs4S7J2xJTIXjvQNKzXFFPzgJDEz57Bxg/1hnT3F2laqYZ875/+a7obG2bfdMH
SlPEPuL64WxE9GRCWFWeYZt5t45Q47RgNJyOHotyujRm1yoeXVhlfqry8Vv6LWPnFD2SW/qAkjmt
qg4rvynDrBWKJRSUj8c6LTf/ZFCupTbC8m87kTndtCMKWu9YvqED+l5sd1/eWu4/sF8mzrRN6QEa
DWB1g9ZbuV3N7AT21TJpQz+qmRh46T1uU/mCUSkAPPBxDgTaaiROyiXhZVDhHCw2nY0+DvJOB6tc
iOr0bCV+vucccKjgrNYFhbrEg/bOjBOTLKfLcH3VOmxT9LovPpjmvjifJHcgCFdbn3vI+wcfBLGk
OlK397UDUuvYDewgHcOwYHVRADVDEF5ALWK5AtBVYGgwhsUpcvvW/sfeZsqJlUtdLclII1Qf7N3U
1Qa81B9f7yuSyXjPKFPtK8Mzieh7Xn8TXsgVkRiRPfydFXcjVhN6TLSF34rNRlhveug6dVcEo0qm
6rA4TRET4nUr4zDIQHJvsgk3NLO1rN0o64M2QJ1pUsUkmAd3qBmxnQFHPVYMLX8mossRcaf5Ff0U
rsZNa4YoXJBKXG4iXjHBQOX9n8knvCt3lln5BfuzDdSq/S3A7iGu64AcTNQaJ1zEcYa5OIROFbCs
oEVMq7tf4u60LWj1uFl6xpJnWyQvHqeuR8o/tLNNaXQJB+tibrxD+q/+Bde7ruId7NPd2a6Qzpl6
nUQ4i+dslU+g4NAyYlMVssEo9IIFXpHD1jx0Y/N2wVHWSHxJfJvEQ//QgQsg8UYvFUGM6WrY175x
VO4XGupr5yDYIeyfvkqRLqM+UqxwbXH+UJrEhARX5QXPYATGSD4UYnK3z3gsApajchn8L4+4nfgV
erY0Kntw8Ot7Ru26MaaETeU6VxO9f3IFiG8iY9CUDXWIUCDg9poas5pR2JoNfkyq1GALVz8IlmP2
qCK/nJdpK2gtjFa+hDmDYtRGzXPCqFbTQ8rpN0jE0pwGiWtjdhkNGoQZ/by/oJuqQ86WiKy6s3rb
9vtmwkuF1FPu69zsqt+Odw4Tfkdk+aqp8a71teTxIUInR8ixH3U7z4TzbMI2+PDrBzT/yGWraD3G
RpLyFCDGWTOxkMfUvprXj1uAdrEa6GRmnuXaZyB2H7x3vMpXHHSENrRJeE7+nCxZ5Bil/ieQoGBu
cb4dhKdLllDfvs6zkFXpNdKKOcpKk4dMy7OGL+Z8L0QW/sSgroyZ4AUSr/WEqYXjDE7jgoYzxrRo
kwjp8FtqDKBQ8wvbZ2RG+Kk0T9EjsejyDOi0cI5z/b55xj4S+rXk43yxjEg86SIqPPdAJf+4sEEd
Erz30FqYodIbgolkdW+um9rjYZ4w4+QBJ5JULQSn9tnZ0W5SnV0Px/YQZtoA8f25oO5gabL8DOT1
yB+szBKY23mb2q+N7FyPgbpqRHdooDeY25qjuvuD4PQb3oavIKQNWG8ITyCrMUecR7r0xYHvfsJS
Wa0NmvdfDmlGfC0c2QKnKFyAASUyXe5he922nPCeebqL6cNTCwWZofJyt3WpLNZvT3L7aLaX536E
KnQfQByM536D/OGclVOgG1FiZNRwjUk2BFeLoMWZedIS8eEmHlqpsVwszbMS6JryrGAeM0Oiww9G
kOPPfFy+Sysgll9CvzGDKDNQBzv7BoF4wfTt8dJdT/WYnsYc7mRk/0MX+wjjLQ/vw9NjBDn1PgNp
hQtUQKSepkUh6sTZ5/O1eBQ78r7oI2n4hgHTbeGxBOGF8c9QaeejKRqwKfzcgUY1rgffKin0799X
JEmpBF9lsqMDJAZIh9YuRfKCmSBCENiaNrMJqx1mDDNslY1h+cliqxOlGmmJ+eoMhUGjJMc0s+AH
pNZNr5U9MbdK+FLcmYiR2VHh7z42ljzVn6U+dBjl1zpwXvRLtKGAl2temdW6Zm09vuayv6ePV9PO
aI/ge26xgTo13cERHZWiYJOtknPyKD3Z1lV/cWFgg6umEzX4Wl6Eciw1vBgMBbU1Te7NRZDrFR+Y
ikmLaf7LenlPlfl9eO2OtBCC75hf0szqUtbhSqI+VI/rq+O4Ij3Sy/P1F7itDEM8/LnpRfH2vG96
5Lq2vPLUdjlwiZQ5teD/gAudmEIJF0l76J75VSgS9sBtor03AkPt4RoZl1XWZvnIoloLgNShhK7F
k63hHWKXr6OmIjBEwthnWEnpDAg10ryHqtG7fAWQQid+8rcdVEGidKOwfaipUj/9tpPVaVfRF6bQ
CGd5Sam3mw5ojzOFfAypWEg6vdnjsW204mZMgCVTR1wiinCzBXkXs7XTDiOfShtYqtTRxBYEzXTp
IjqdUrdiSAWaBECvKJlRmMeVM247YNb5mdMG8Cd0+ATKnyWVujx2ZKpQhE+5x6KV0TDOcnG6jDeo
SmTEwc7kmDG4hEJIRphioRlV+/THQTEDr1IMd0Rvye/X1f3FHTqHZWn4kYUf7hMIfZ3WoL5k79T0
l7ax0zyAO/93+R4RrrMRjipLKCvyjxoKcCWXjEHJLhcrcsHko+V2ohk66tHs9KGdS3wIJUAiHkqb
tRyGxCcyBJdN2uxJ0o0tMWZ6Sm8+gkHQ39iLyGmrxA5HbgzxJJujfJQh3lkrhGrembLDlcvs9add
qZemnwX5npPgRm0KBg2ck5DDrBOtI5pLLeAXfr2dDn9xy+Y3n7d+sSQtBeDC+8R3+NC4/m0IfTVX
jhyOOTpuN95bAoHz8byscAVEzgIpY3NZrb/o+tPLMSN9OrhYUIMjdhoKxVj+4Mc0ASBTIFGdkDWf
mQQ99rJv/j+IgzwF8dGJQXzGj0otZ9lJUTWgsYobWJn6avi23AxPrnI7aeXkH7BJHjJyhnurrX1x
oIYOpfCzP+yBeYMF/6OFtxRZ9yrA/37uVofzrEkbnx4eesESbOtjQ+EVlsv6Kppx3EJWIauy9GQE
x+N1xAlfn+AEnCOEKH6XksZ2A5W/xaCAv51vyEpf1PEeZIWyfnMK/b3FL0T4MnGtLlqZ0o2O/tR/
oSWP0ToJxQeFX6rcQCcq3+/KOuty/+0BKo+2EhP1B6teOcz5Xo6HPRwBJy16ToU0xu9pttwpv/n0
Q7kQ332yZLoKSNgk3konZsxky4nXGVyO1rvv3Gu/2W26PCTp63tmz+yA427Z3bzHRhP+0PYk8/Lu
9KTRf1e4Ot3z2lo/iRYlC//o/zHw1qw6RJofnn1pJIO2MkjtubTfM3+PTh/tGZ7I7sEeHVS6044Z
mg4Eed/FYhgRl1/lr4yoXIQOINdeVHm/Uq4YGyqGtpxCmOgjc66u0Bf4i+tCi2jGg5gnZh27BbCp
h9p3Rb4hBxmOjgxbogsl3WMD2n0B/jTJeye89C3XUcV8/j00g7I4p/Zn8VP3LbaNn/aVGAqbpjda
lxj55LSaHUf56P/LiDM4z8iQ3T8TKLhvzZOIR+fuHiIx77FJzCcrfPu9v8oErwAUzb4FIaUmmr8B
Zi25sOoEb8lQ9eXKzEgdJVK59gEQL9ue4JWGZed4FyiVa5g/TJZNoO+mBBjvPJJc4BCLytb6Z5Mf
T4GP6C1Tf1k3MIpwIVq15CCtVxg9vFcvAB680FBM13oSgWMhRARCupNNxKMHe1/rIUvmJHSINbhx
n7XxAZ5W/hpdFn4aB/AtYJSJfXzvUEzhXm1XjVEpf6JLeHjhpJa8EqSwmfxsZtF0/nlIN8Jh/eZz
Sc4rNHtyACK55RVcll/UoWwERrCxfAVEAEOSXQhO+7EbSA3zoYB3KvCo9RIAns1l0XVxcip0tvfv
nK+ja5MZrfiGn0UCpDrTkFMEECkd8H3hQpwvC84myGUObPf7Ukd4SVVBW2+oJ+UaBdhb0WjpIWfI
e6MUhVJ8tD2L5Htkt+RiXrzJY8RvBefG5FKt2Z//f+g67b+RR4ygN/l3p8faFtpxuR5779OsQ7Uf
dMnCrkZCEefVwox6+vvpgC5OEYBD3rFDDE51Q6C+Wgn+1gyTrD5hJShzMkKmcwZSTbAEGy5O6eDP
v0+BeNswJxxSYnXdzck448EjpgNt2S0wL6JafpVYZCF1QYB6qnitCXrrMuRbREa3U8Ymqs+ICQaL
qwatKYJlVWjDP67UTA3sSmTwksnUDZ4KdnInp4ui0NcCx6zwRYYmleugmQdjgT1neCslSuqAtVqy
1Cs9J/BJ1rRy3xNUbuN4OgWnRFf5wQF01smBOsYwQ6e1ALWgQ4I3lOHtRDE/OPaDi1pvFWGezKzv
JFYPX2prLUUUPLZ0aB2Rb9voEuKXFHanjTajqMSEUHBrCaXlaMwYEIHR4uFIjSuMoZ0I4DgMKNzx
em0DPUAQR3RoAj7MPBERRMnUhDL94hTzNty4QoA9/IjFHV6V8skVA0keSx4KzX5SgNlYngMDRG89
UsJyfTwHjy/kxC0CriQTrNZgx1IIuoW7arPogwnp1kBkoKrT6vuuJMdbIPHJi5NExawMhyJx0pC2
GktqRle+KNuzw4Iq6YcFlUni28G5FRJgtnrrV6fKQVbHnePoFd4ioT6lYst8SJFYzOf3AY0SyPR0
LVq9fHdz96gYtHViSk3CYJoGd9lTZsC+zNKA9p47HNzJ68bYv5dV+fSnQ8MqxYGszhtRkZMhWwVn
iI/S6SV9pf+0w8tubCuDZ/SC092jcQaEaqGwaDPnv8z8SpySG8Hk25FqLHnOKzTRaKsIDb1yppH2
6OxXHMQ2sPm8JSK4k3GL8KFN+kdpapGv+/HQ+OdpW7Z7ofaMuSTFkHCUGWw6NoPhyiICpbbxKICZ
N7D6d8Eopu0kY62yaIqpPWD5BvlSiQxK7hZgAMKpbwELeRCD3MR5HL1ny2hFajbcGfQu7gQpDpKQ
RMouiDoliTqlbHIqMhD0I64C0ZdkjnFsi41/HKgfQtwrgB8Eyscjsi6Sy0lBlRJksrwq9worEYAn
T9diDVOkeeHXQMuj4m9sqVk+DMWwonVJ5MjJ68UlofUS8ZuBURWxlQJ53zmvQagTpCyox5sOrhl3
TivPoGFSJzIKb5rnaZSepcMo+EFiU10CPGaYOY/wf+y0jLjeP7itgu9e7yRnBAAXAOeivng68M2v
ISZuCo5xPlOcpagtKrUbDkFzzFci2hUfuzVh9p/cZXglTRFZ2Ei3uivG3vXzA1M9kCLbymHerdhR
rP4i+E0uDnmmj/GioKIhwmiKwHkzp4NI1Z1X4qMt+7YfbmG5bPdsQG/1MZg9bhTWKhNtMIg0R6+M
NwTEaw7xUTzbGD2TWZed+K9YLwd5L2jNFrUQfqxT1Xu7AlfnAwwsBpsb1zJsr62nCJYgrn7dYUSK
5Fkt6bbJ+H8vl1MwfwzRPdfNhVkIfD1/5H1dPOfLQ5k5aYBIMYQRa6ezFoxbhRyTYxGOFLeym1tY
LevlDeE+r4Gr84texECC/Jm/h4IPIDj/MCPJ9SCSkEmraZNmE/eK1Uq2f/BYjnphZP0f4PaL4hMv
uVg/nI42d2ot/FJ+88by3tqh6rKaOtaC8CdtrUDnDaCkAo8Cb0rjD4ZxQxUfq/CZPcex6TIZtmQQ
hd9D2kHOIO5L8dypnhUZ4W1NWJzqg4wutMoF6nFnjUfLXdN3p7bDl/9ajMwmmiQ5fMYEoXUt5EiE
SAc/+3O4pGkdvzdKJJjSdCcS9bRL+kR7MaO97pKh4j7v2JBjGfkL0EGqBfIpdSnVRjMN5WyAVCZh
vmvdotYUn2U2NCb9JPKng2nfPJUA4jfHHjbvgZsS11+wUgjnvNFUD+HKHYLJwKEt0U4HLm1S3K83
dF+rm14Hd80AkCM+0F9+lRjDvdtft5/MCRqKiLFjLq2X+55DWju9xPK+2diaHvttpdM9NyYocdTr
nFJoYwkr5hdtxtImu3KZ6iAmUoPWcHO8Vjg6s17MTuYraw7dwFbyvltcB6kG1CEooBVIT7s4d8BH
PrP2zzkO6Rcalle83Y4P9iwRDNmSN4PPiO5zFS86+9BJjW6bDApbdLm0TJt3mSno576LvPXjuDVY
uUd67VcUHxeGRmA617uOJfJ+am7M6geTdElFCbB7lz9u8YRF7xZ1yN+8nKdzAwNsstihCCiy2tF6
gqBZEbqMxzTpbD/6nr989VqQsfD8TtzQe0ndxs+8NH7qhumJDBhkbJi6FlgLh8oLUZ8/Scj19oUY
dWfHntLXtJ/YBIanfXcjWQZRNKzveiILbpYFyXiXm0NP+X689IZTzoXsjo6qqTV0FgzEikHm2wf4
fECW63FKpGDGG9T7+7shPt5+jVcKT54WmCfVesOyJ+2yhEiFnQofqCepccS6Z5f3jS10VH18Hb08
2g0Zfdn6hdNpVXEL0CqJcPmpbku1SNQxmWNeVsURgMLXVeChFkS3JjXTUwEtFuIXNWbSg+tUrm/Q
Bz6MTbby49VZbkEvMdjHLsTgIBick+j9Sh80iOXGC26BY1NHEMeGMD5ujT+u5Kgqj4TSh8TCrV27
42C0HQueLtkBaEtdvQhIJI/aBFYww+bKMYW2M/5PxHRuMxuflwEfNcszuqXtFa2TVg6/tQdMtNrt
+WkZn+jkKqWJBcSEtWPYUFg5FcjwzYnlpGjWg2tWQfogbwTcXoiIQcBfW5/UZqXx/ifQByMiTT/w
V9gJz2wB36qtfME81upKC3rabNf7fhhuVvESYMyCNYcABxt/7D17pcGX7jnS2bzL/HdU2/++Y4Qf
+rK3qMtjMnjPwynzMGhTrpJmhKNK6n9SRfQoOPRLXcYTpK6Z9i+WxyEFlukPpvjjsWNYAeQyiL2x
tzelhEpaBX0Obfzb0PWJQ1fKqlGx6l69qBiFJ901NylPeKjgdiCtoZbXPrbxcy+CtWSdRdMhjyig
aXr9JMye79dAdAIJg2o03lqIbfXt6PKcPl10EGeJ47p7xWCuoW4/dVs7kQ208yHjFwy17dxbJD1S
y/8fCq/gdrymP/foVujFz9qc56xcMS3gTNAwg4Z6Q/Ize+74bwRDoVzv7Lz4kTeNBJfvqYDOedEV
vjI6TeL76E8LBY1ZQiGWoCfHEDwDmbaRZlwNW67hBumiDAi+WiIsHE1nisz4BOWNOBPuouCGDaNy
A89/9Dlywj5hdSJSOBOiB8+f/W5kQQNo7iUog6YznVpqra7drqLscPs96nttzRONXcPW8YQ/Y+BA
Fi3QnUM4YRw/AzyiKlkEC+pG1Y+pXAuFVnVa/1m8BQnqHx0p1cFllGcECrfo3afmMp43QpcJ395T
ftRcSbRXBg6SGuJ3+dwe3psKl38/sfPi2fv9Z8Ft7Pe3X9zjbOEoW3tHjyrwf9GqEd4i0Mt0XQ9W
r0y7OuyhbntJslI17hVOAyPqjDgvcH9FbRDvbN0/7xjZ5DxXJ82FSQJe7UR+gKxcyLgrEjwQrR9q
2ty7f01kSyYUKtIO+LSpQVnWhFzg/GoJSoArKXl38xuZLde0ifYYteKu1xDx89GM9k9FW7KFplcz
/5ARxxhz419KaHOTtJ5W+8Zp6c4PzxbWCtcjyC3wJks+fCzG7T7LAyZh+dJDUgSqRMZoqyZgfAmL
mDtwq1LhwWsuuB2BG5WIPCAp0A8/kqqQBz0RunpE0ad5roqUvsW6ba7YDqKzskF2RkH1XFHPqOV0
a304KVhZAQ1wiRDLKxIj5AolqasXjjloOEvXFAhfjV10C+bnsjG8e51i8isoxJgmc6kyD0jczLoK
yLJoUAE5qqz4JLIaerzRb0BfudaP30nROeu7vZM+oZYVTQkO3ixpx8zSjd8etNurJ7TBQIK5BP2h
/4ZWVPx4EQ961pK5RDPWNatdMVEbxOcg3x6szc5iURLtw/g3NwTzwJcbAJ3t2n3E0sWxEhZfvqAe
1jc/geCu3EUoHzn4AF2LcQ9XuY9Fdbu4p3TEPY/oQmZYQzLAJsfSuWvLRkUk2FJ35+Na5GTSAwHl
Zjmg/G/f/Yf9MhIq1M/8EYHgCg0Fn7PAEXz2/0sZvuQb7cXjOPBna6UBinjsoqnFURYYVU+miRNz
Fjb0gjbeT853277Egnf/I7TYoY+zQosvSNkuf7//DPwxOSTIeoHpZp+9iD16AGjpsAXWuRI/CKsL
rabVzaDAOsEbc1hf7y6SDhAaEk9CcpKrJVudhKwUu3cPGBJ6FGKbVK2Om/1wTFLJwQeoWC007ZSB
QIpwMEII0JltrPX5MCOAo7CHlI6383KXhpsZofRoN2pVHP9qoW4oxnW7Qv8duQIBaYMyesVKK/Aq
8sxs+l5Df41W7uK9LMDDBXWcH7ldxzxnzZljjbd+/oIwXFWD5qvE//sIHpKNX1IWtLsDJXjw5ttp
czCTObhhFoJMSZTnOUr8MwiO7N7fJ1BfUqagjpqS6My8nc+/i73xiEAM8NuLQ/mCn6X7WhMeYzcB
jhqMr5J2Fl2OcTON5drim4BYkbBZG0gDIETK0fdfREsHZGhw2+tmeFA4okV1+vnCdaY9GFdxcuIl
/eI3AXlEox+cc2oDndQzljHJdxFRtZcY1D1QahfoUvu6gnKFPlDKL1B+H9hUcP5ulTzpAZ0I6Ax6
Af3tDyPG9vAWk4jIzU420FWtciT/Kqz1weouN7gsTZPU95h8evZdHRH0R8+U/hqkTXa5x+GiLmGA
9QuLvjwWkZ3MjkDtv+LzgMJYxgu8NG/5Kvordwt2caiBeTzpjyeefxT8iSsUOBhMMQuGQlI9hPYr
RiNjEq2wam1Q1FQuVxRgcDeAegLMOuUQCKKN8bNbgCKY/XvKJrh1lvpajlFPmDBhVfjXYFWroJG/
3OQbrAL5hzaI2manZhF+eqrrPE2stn5NnPD9o/hpER6QzrhL1rXrfOIkVekSmwALx6dvMT/VpK6O
hovNtzHH6sXaE+kjYM56ActjZ9rQT+afZezy8tsZ9BcL679hwqIfZ2qLF1a9xJlRLEl7XzpIcZa4
wEUxsigxxXoh0rSxe8RL/g8jGol/UVPrJ4ckU9trZJ4umFdR7imJB+RAUSooC/9CLAj0m6RyZgOM
B0LZgj/nV0B8SF2q0GgBZ8Eep6yxxcvgpTPr+6IzSHFIzWmsitCAttpjy2DInPI0UApNa2NNGFP9
HaC/+VcJood5JFilvGlU68v7yJXAyP0FjDnG3qiZDjTAcwiDsa9/ewFbXXxokecR9D9LBa551x8t
Gw4ShVMWwZe2BQuoXFSkDh9cQ1tKpWeXBkqp3wI/6YWFdhxUiafWk1CZDyes4Vze5QEFDlsdE3oe
ASczu9MiijGpsZUEMLIavsRyJdXb5194wOWN5sS3uRIV76WR/QoDqS75GZByBJ3nvG+BeYrMiNto
Bn/dfMZ8OEedDmi4mw2zDN444LmHL7GLCSs4hkLOhB0pAqVQpDwvYUzgpxP4Za0h8OmFjGvuW1VS
7+de5FmYFY310eQwUXqOS5nze47CeZpSWygYjokRak6OnSwGEH8A/sXvU3LmaroKXZb4J7DlCnKR
vREiQ2OgoxsZeMbUqhF4X65LPdj4bYpY8L477w9CZku6AvJ+Qv5mvdlAueAYuqsDBGIKT9VGtYbj
2rPwqeTn6fR0siQUdrRcX+JNrtAEvM3ZALC3UcqtmOe14fT4S4sGQAl+QHcxhkGKssd0+/JF8FJw
yg1ron7ckabbySl7NzRmYMhgQ+P3FiXLz9WpbOif5N20VWtwhJh33ksMty24QbGT0cKb6d7mTjrH
1BE1yHjth8yi4msCBX0FxZtxibbctsz5htaaaxzen7/6nvb7njo/4WmS3F++/LB2y9D//Q4joRpH
B7r69PfSzAG1gBS1/m7Uctkfiodhoz4tlEwZ/D8+PYDRrtoLb9Cgi182Ql1h6d/S9LVRzpApjG40
KWHlQdAzumpRvpIz//iRjOTBDMf8SRSoP3XKK94pxyZvrjetEgbfjca7bi8+5I/fBeYDCRn1uWT8
MMw+Uk00WfYc8fMjwW6p76lGbodoPEgYAgfrKXVqpldL28FvDtum4zD4DHJHOBjYk2i+Cr7ZImwq
B3khfCVs/D5YM4HX8+388HKTDHHIAOSCDr+PSvnAEgDS5OZ63G2DkUqIm08xqG+9ubLB8Ofd+Ts8
3zZUsSd4oKr4B+SvJaVdsdLuF29I/kjOLmDk1IQd/h/2eg43i3uyfS9kFiiWwVL3PWI2Oz9jDQfG
DeBPQ3dS7vu58vI5Y7m0O6+oWQLaQ95wwMCKvz0xl3onstQ2lNneZmQqOdyNFNbOH37hWkZaaucr
NfN/3e1AxPoD+b5SuWDExxQfZsfKcFLgA82LIKegZTjy1JCNQsvgjEPCdw2zDCWve+51yyaP4Ppq
T1dkGNudcLvK0INLvi3qNgRTfl6Hvfi+KvbgvRoPLFVF1m9rlw9D0DNKgkUMZO7bjYpbgukvu1mi
OUJmgqxlCFYK6tipmI7Db34Ojx/E4vd5XhrHTwKmrXJDf0G1lRyXSx2CDhQqm9r9Fr8C2ibKxArX
15/VulToof8sXI136jbY8v5OEiMHZ70rp62OcN5O+Dr6WqUfOvFqWpEJsIOGCs43VwJzkhNYNbjg
Vmp5Nbl91TN136UbLofXgUNafIMsF7fGU7HBgNSKYTPkmpdB2ILo6wCDHPkRWGWPybvG2ZlOMHHE
jbH/9rmnwo10HEBmhJmYt5/NaYKvtqGFtP20EUgr/NufWrGQijpbPyDZwVLuOkue905eA5C3/Irb
gy0UDZkjyB44U3P0LZ1yZex2n5n4g9DAq3FGaDlgUri0U6MNp/YX5ZxBIhG0FjQ82ItgbCseyLHf
Or3SlAKaKhFfpO8ikJr5MqvNJFsTl97VGu1oWSaXPlB2VmXHgmvSciufnvcrDfmy5xKAfoN34bpf
r9eQPwEACJKiqjyEHvqTbZnuyDEfoLmavHaNFhjGoQEcsycgyGrGPgc31O338MNTSa9vqDTlNLNq
eB1VmKtUpAl6dE80OcJCNA2J+kRGbap9t+3w6Ao37NoysuEI4dqWHbOYVAi2Ta83Z8khLmD+YQxP
TEqsvgd2+VbW0noHAHuhDmwFILFUMF/oXiXyUli1hEwF9gz/E2oJZM6i3c2CtWuceIrZbN9TfivO
CRbnY0HX6u5Q+HXu7ver7NIXW4PYKP/x4MU0HFXaopzdeXyEq3mwLoAd3rjI9bQPUe7EXycMH5/a
OtGMJLqcZNgyUog/uatkar6aHImA7jMiB3DN9ShAYIrY2culBc9RHuPN5MKaaFNKcVK8pmFmeNok
sawNlQbmNkUiAKnNmvQ8267r2bAZyy+pXUPgCTT0xesmJeEJBySiWOMj7ePMSLJFaJmHFC2u6dy4
WF6ahJCYYUPWNZEs4yBgKn7a9roIop7sK/GHN5uMjFKE4SBR4j+4rQDg6zoQe6SkYS4HEstUaA9j
D7/cest6eCzsEUwsKW2m6JiQ3wv2EOxFY//Vhaju3zWjA7ZGOttMu6LVGwoubcE7EuDYl0ZHq7zz
7xfOYLi+RczgUdzBvy4l9i1XUzRR7Ii0PLrF9nKlvYODgkAV8z4v0TvcP0JaVAsf+gK5ZusEmLRa
ulxUj0qiQxmxnLxWXbJaGiyLyupimK3dokkNqDJjrNdCIDhqoT6JzvliFnFj0Hrziu1cNHH8JGbK
k+zJh8dvIjtbSKkx4WJ+cVGDkWl9MsYCHGXszBCycPuMg2iOwVZkk6KT0+9LFkaUExd51mByHsDv
Hao3KncvESucdZ+gRRJl0l5r3NrMRJWFlini/HHGITATtbYnxFIt//t8bqU5M8MuibI03m/VXOAi
TiHk6Sfn+jRKFp5AIz091Mw6A8+3T4vw3MtZdRZ1R/pBl5xMDUtEqGgC8897dtKGKXZ+cRfl3R3G
kJuZAjlZPzk1IITiqyrXnTRZh1qybU6bae6j5zncdCM2WtlJbhlpFCNOPIIMspH8pFvyiD57/Fx3
dNcIvlYBY3twLSBSQLxd7DMu5/jFmisIzoe/bKd4B+hj/QKlrziW49yuFHPLwSYP/iCpjLVi+UQi
Gp8D60A21SEPLBR6RapNF0zSVHQWRvyW+2+6iNhNJD6A2wPe1lnE8k+8ak/kYHWKoOjYCUuqokzD
2j0huO/kd44ORq62VxhsSC0LILk64LYINNmngerB0utpLo0t6xQWZmsEwK+Kz7Kz69wwHPg6vnrf
Mq5q1VY+2GgocsXORi2n5HNME3tcFuH8CxrIOgLRcvS/cd52IcKe6qevFJ2SymMfMrE+V1LXvkLx
WSiB/YqCeKPt9DbtWcQ1F3MbnVLaoroGOw6+NKad8EKM5jmqpDe3whgH6Xc13aBfFRpCL3IntXZ6
Yd64h7ZspG95IixJc2fzWY/7mRt6Nm8FEt6rkUOEN4HxQ0pjndXX5Ef/HWV31RVtivpeYpbhWxjE
kJwscksCqRnngrzZai4SPcN0BJ2WOWy3I5vhFDZyWGMVoFYnh9Fe2SlNUwU6Y1zfJMN38yk9Ngen
OGlbRF5HmR8Q95BoXyp91peZOkIcvMcfCzXZFF50HX9Qf9Dhrk3e01Jg6AtYN9Y2TOGRb3WVYQe0
OYcAaeslX7mgR2nvXI9ljQwi/W/2GCYdlw+NXek5nWR8rkeBEcWn1/77oA6Rri1qQlp+GsW6FCDS
hE81D5LAGuQjZxfu74wyyv/iKyOjqGlIrLxL8LImp/pokuc06SNi5k6C+JfIFBI2p301pyZ8t/i4
a5pTJF/e0JDQ5Ps9BTiZqtothnMLcvWlvEYewLmkx2P57KjhmOw+Dn4YLaMyyIMkt5FUwMmxmLoi
+ifDZtq6C3nvSGMdTl9j7tBUhcX0Mdl8lPDzCXk8phz41VWiczVNvstz1n5x9MpwfTQsxpveESDX
5Xittxj1pGbs7u8BxxXc4WYoIGHOrkOZbcmjU7cC+/htX7TRf8H6ObqgopTCvgCEmLhcowFFAY+6
bLJwwAe+qRHmPwGXKqsBfUrokSV42NQoOyOxdsaYXwkipLga6CfWI0/3r0TSNGcvmO3YGiI2p6vg
C+TvgkMQbYFYUBNG/OaVtkRRJdcaTeLxTmZkWG7EouAjJ76pyUN27m7NH6nsQgXgyArddExzCasT
burUH8rNS7mrMIUuGLlYD0LwsLim4KwCcC0gcUWwo+8U8u0fN70mUIgvOOLZFB+9kM1AgvA3nHsx
65LUwfqPeN6ZfkCVTvDPNYTVlH6Dx5bMvogGjiyX1BS6iBxpK6rWGZlkpk6I//ZQN/SFiBkG2X/n
7KJtrLeeHUZTjpXVn1yIrmgI/yZrFQGpPfKx7PBkSXTir6oIaytnlxbb3qwiLwmPgr1cYVP2x2xv
oHZjo74lNks0tItUSl0kf4o9T6MNV70e14uBk5r2Dty1WlWiL+oPrp05W+1lUimLtrYSG2GSFvIg
gZn1lT7ehctgsAT7BdZJpUEyG4l+qQZpAF3Mg3ez6QyAzzDi4YSLoEYsx9dRnVpAJ0KNlP0ITpWF
PlkRamWd3CxgU3flAfPMNMrapI+2KIwUDfZP7jseFfmGXjhN0gN5fUEYFW1xZPiI4+JTr76F8n/k
9zmOhRst/yGxZec/13nKm2brsEBoVHKYEBPobgJcKjU6OBG+36SUmiVqVAwOcQ1QaUn2m+8GFiyn
5WwP9U+28YrkvUFgwYVBiiAxiuaIrojdgVF0qVxnJZselV775S8U7T82juMHk/j25bhwbp5IhOCR
FSjoSSEXYtowSW5ZJQVB98caLLGgov/txmPRIWCdV++v0A+pnd2BmBITTLlQRHzIskudrv7zy69j
e/vVUxmfL/l5H/zwT29mxNHcZhJhdGkys5vfiLShS0/R8d7Dscy1BCkSIK3Szz05q8Fh29BbAXIh
MOHqBr5aYi6CQdZlfxRgFRdsoBfHzJ6decfnFOcRF6EVAyEQKm9ttxbv6brs6R8aslQfLtThFQ26
RGzmXdJJOaGyRPx6CNL2WKkODBYvtLuG9FrwqeEZw9hhOWFnY8bNKq9xtKjLOEMQZv9d9d/ojerk
JF21KiD247x/rhl2nwLS6R9vfvqd1SeBI7FxVNeDWVHbeLYFvO860AG8P1NIrN9pseNHVHTj5alN
/g8jzQtMG8fjOmzvpR/8UXf9B/RxYZrcgz0YNKqOG5mf19NBPHR+E36V+V0UxmAj6t9G+xV7gsKF
+Xr4S0PY6wbtZEqx8emGniqNowvveYv7ET5GzAERaNT1muepdHowqGGmDWlEhn4Un5A6ddfgEGHx
ItjAH8WuNuuYZkF6nMo46W5LJSq5fIxfD4CIwM0rgsKjnsjgL3GCMUQLZwxxilJ06Ny1ZJaKTcde
2yze5SV1wn0CX7fomauHqX9za1i2mVY6ktQSCt5YHhPZ4mMFK+V8ECkBkBnwj+f6tFr3Nf98At6/
wzIGnXj5CGINN3IxMwvh3HxQIuSDKLsjEMLQTmhWMIKTWYzIvdCblUS8E5z4ylLsWnGGEoGK9Qr8
DcUnMT+GJCZzrqVwchwH0NsSdM0newaqjIM/rxVU5tR/czRKcXW6ZCcJf2tqwXhTyWwAK/rsEy4e
b/VlMIvzapfRLFq5IdAhdVwhRcVUJ7ZeCcgkSc2+9MbgN9NRSwOOhvj44nHNudFJzq/NQA4HIWXP
BDdgbfSjqb1DyRPuaNw1AIS12gBHMM3vZEDtMa+53T447J+VB3ZSbNOXvxYZvDs4z0OUJO0Iw+hZ
SjLYfBxXpTg2x+33DamTGfcGcx308LQ1dMre2Uf7XxhiqOJIQP9cxCR1PKxtMp7zsTB4XMiw3nFL
IuJUNhsVeZHz2pgdshBo24dtk01nM2rJ/5+usSl7Cv2Z+t5IPoyHTWWhBCzi+Pa2a9DCM1bK3Gtj
eaodDvBgYfsykxQnw+++xzEBO0wFJkZ5N2/fR8uYUJy/Ow56A774q0m7o8INjgJ5l7Za5+Tt/p6y
BnHjJ/1CqSwj7D/S2i1BEi8ITsUaZXUo6WSDxHabKf7o0/w7/m7xNPM3VwBhqyZpuiMneyrFaFHj
90snI5QyaCxMEyqAXiV8ayLruxM76OmfaDszX10VfKNZ4uAT0s9iw/5U/5kgybsKNdV6I408e5Y7
OAII/HsdBERm+90SSyQs183MzaJgl1/2JXCrA5o9jcfmL/sAwkFZZyflVZDQ7/oCwB0mpQIEfpnd
QEWQi3eIUzN0Dt/FvFhN58zYEqq3+ESX/Y+4bfl8Kjx3N+vkx3g17uFeFRHDL1/OMYkolQs8BgD0
ukvntK+xYKCIY4cpokE51XtYw1Be0kSpzYvFpcj+B1a6csx8hqcWiQyAh0btrMpZGBU/LWLcD0se
hejjUh8O+SGzyyxL0qytdeOOhv37tZKYNONzG6AcUkAJitQIlf7IAuu6fXDRpZWZ2HKo6giz9STn
sRzLKVyDUs/2mU6/L/nQnSAMloBTLYZ6hYWutBeYpHYv5FyrqGOINH8JTDP3zzK0krwlrfzILVAp
5S8OkERit4DKqZ6DeOv+/IotaNoFYfo2aY8ASShFOZUpXS+6OIzkD5hjxK50ys0iJW0Kp5zr+xV6
Wr0KSgzSK9aRUnRGep1Rj+3WwvgwT3EH1xXU/PoN4lTdQU5Z6ZODuWZ71s903lWoM6qyNUsY1nKj
g6a4D9PkJgXYegZdE1qPEW+vwWaAZduDiZ1v8dPCSqHbBXjHabDZG3tfXzzgEPizSgtvVRKbPCjk
WK64DlMewa4Z9BpZyUFTh3FGArkfu7nwYFmKx6EKLX/Ahr+MWxMQMfVv5jPpWpRdar1FAVVLhNmU
tF7O6zUX02WKN3V0BBA2Bw3Y/mMPPoaL0bajMZQBxF8u07RdH9Fj7RiPzGpeE1EGWa4oTtHtJH+N
PAOAMXWrOiYL+g7JP1ce6kz6uGI4SGSBPIO4emb1oIHk0TwymNQrOtQF1QtPBIDlucDeM5v0IBG8
ErlsJfISEfzT7YoS2Pp+6dLgkOCu2uBk1UtYTU3SwgAV2E5ALS48hLF4RTahCDu1LlKk+TkfPNNH
5J953ObwYpLvQMjrIHTs4vLN4yTTXel5yZp/wHCQ1wfaGOeJY7zkB1caHa5fbFBqRXTdJ+cfNUB+
TJ7NbL+T5FjBu/m3a+l+FUU8iTYuTBMI4NHIkTVmyi+DF/6+GVMJe3X2LNEt/wOWOYRJmzgBdrk6
dkr2xksBpbg39vz9ro9WYScHwNOoxltWkm2SYkbH/jTXs167M1BNdFzm7rDL7OmJNHkxs6VM9nTr
7mykm57FN3RIbK7kY8WoOIy3HxwwuEhFMHAqq6nD9M6EQZO4gPSi4zyZzn2VW+hqk93qWoi5Q+RZ
GeVh830kBC1oOkV2ADlcFkmq1LlVAERKT0bKwcGCuYE4o3Z1euQMq5o0pGxuHOsyEaEiLBiZ3xi8
xLIjKkVZikJn2tfSna0WGculOXdtdAJxb1YOq6yFcBBagCNvsH+L3zV/sU8kfNbmKuup4/TCasgA
CrYrADM+OolCP9slg2zBNp5V9+y6+1v6WX8w0RXerNVtM+Y8L9NQ6oNY+LJDAZc1CgChkrt6F6sA
pEQrqv9LQIufz/GCnXf34eaj/TJxQESY0s5vCgNV1cYfUUeTT90CkiCCxNoOrq+4d+kzsGkSjVWi
vVeePDas5Yb5GpU9pyYMwxXjnKnb2d2Zx5ICPSmz0cak2YCM/U+UnNL8jkcASldIP8NfOaNNcZx0
9vxD879WefQSlgopDTQf+XxpSnmJyHpIscJ9VGSLhq5hX1d3Wo1AqPZTkbDNBHqOMU9JbtEyXSI9
8y6duv2Zv/i/xPXH1t1q3+8QveXrdOKf9jU4ScZKn/aYR6CPUNjj4gkGF+awk4PrBBXdwOe3zEsX
U34uuZUKZ0vQYHmjLmyO5up/BtAP8Pw6NfNukdPHHY6I37BFbXZ371wsxkARPIMeASmxYWcDWOH0
ZotSsQsztgP0c7U7tSoXO3YX6fuWGm/34l1zUmNK2zuycG4/NHhiWjvT7e9eLtxtJzAfukfTSOd6
4nOtV6DguEX4lJBh0hrZiQfjL4luoKLc/dhwAmlht8ZNqv58kR5Zv5GwPmnf3+Vco8qtGkFHA9Na
u1JH32H44n1lF9k+jm3NTi4+gSIFFwr6y744iTNbLgEK2s9qwBOl3zhSBmjIQ1wSL3A2qF/KYJ3p
eMS5b+T1Ni63Wv5X+lECaNe2hGcCnMhFS/eHCncNhpUZ/b78+PHNndnbSYB2zzg0dHtlvQZKy29D
deuI059cgDRpu75YoeENHU89/Q4/InMGrVwHFqGgq/Cup/ePKguAOq/65v5N3pq3SqeQEi+KJcVz
jL6u4Qqk6bUe6F0fBrPAvGcWOkbmVwt9u04RUzpoFXC4OTne5CkLmuyqdA2tik6ywROjZfM8xWbi
UK3csKr/+w6DGhZU2tsWW73F42SkPHFvu8ny2Yqlq8M9TWQRKFqm6Gltbwp04vS8Uim/9kaONOF3
M2DNX+TonqKMGfU6GZTBWgwW8XFFzZUXLdAVmvnPNRvizmlNUaZcXbXdmMd0QLf/AblkCNXMbLCL
EPXlcD0vtK/hHMhkyiYQBUqn+weOQjESyupFvlbRBzF6Xlmnx9PuIV8iytM8obGY5pGbQFPlEW1Z
p5UXOpbuoTsINBN4ONLAopx2TGynHOaF7I/krvqkZD7YL7ji9qSTT9HsUD0lg0/Vcj4+INLKdpq8
vky1sHlmVjAeGhALyQnLPvLV8eiIT/tTsdO0hjatJfNiVS9zkMhjiCZ9RD/l6tWguhSaSp3IetwL
ja+GKcfbIHelsqMcyQzN9j4iMAVc+SQVsSiPlcn37VBoUNH9HQBj6WrEwv/V7hR18FB4dR11ykS1
YtPq+A10TB7KFiBUCYnvfuLn0E69eGK3tcyo/fIy6vJVgrpCb6T48I3p11QOJZRZ+2qw+DWmgwxG
ggx5DRdUCiz7IXLXlAHdeMInb0iIRyUWJCS2Y6uM2ANs4MBN3a5vYxHiMvFlwsLVTjoqhwXRn+4U
Ix+CxCXHnYT0BGD77s2XVj+PG2HBOUQk32Q+VM/TbQZuM7ihBoKsE8jX7BN4KwohJI2GkPPTBpl+
X9F+Y/zWaSq1s5yhN4VUnx3sWn4Aa2lHplMqWhgWeNO2jmKzV86LkPATIEsAw7D7GFqrjVgHStTv
fjMM5XxQ5k/FxHk+65UlSkPVIRz2uIRRYFO6kOcLG1noAR4pKx1aiGKTzyFUA0AdAd64+chNPzqH
v6aQ4DiWIVv0q3JxgI8oPN+XqP0Et20PH75OKuybwetQwVoUvtocd0c6q8IMitP6BxfWVuwyK+R1
JW6iDOWHxlIPmhT1Gf/J+hNDB6jxrqryb51PkegdwUQseAeDAQ1FNqTr77UkH+vj3dRxrmzzyxPP
vWCs/zqJjeiR8yJRmZWzjcsMZW/n2C+ULs7Ur4kdgc9LX9OTlqwJdl7ZgDf5RMSlGfrAU0HM+STh
EOWEARGYvkRMrx5a70f8L1IKJpp9sjCiUs2fEGrmSNmyZSPHh3JpiS+NKrvj7AcTHvGgQb6sF4WU
ni2ndGPDcHFPl/KxQ9EkNHxJ6uq/c4RLXL/xZheSGE3loZk4RVlE70ohwpke/4puJjy5PoGMSXka
ksDBdz5Xc7tLl1QKgo+EsO1OQqs/fxm/DtCU75YHT08K+39q5Z/SojNDcJ3dd2D8hasDmANvOI1A
oC/TO2ZAsXKSREg3Wl+iENgVhIgGSSeuhsCbsygCOpk7enZUos6AyD57JxQuYUrBLy/jLsB7SYGK
CbgsUDGaGPiI8qxeD7WWY46JYHEsfWFU79Agy+cx87sEj3//Lp9HU4CVXDrofgJXkjNUJFObMS/5
45eCft6V6v6d4wa7b0EvQTPwfsryfQS5wpXC8cP7sXiAhcsEo0rAJBSmRdMRQZ/joCZWIeRuv8nP
9pDh9+7fj4Xsb7iLwdFT4gxZovvluBoc7G0QT5l+u54CTZc7HOpX9QbT+YkJDAzHegqQuYhdV/DW
iGwbtiiSl6t2dopWncsjHCltXqc7aYRjo2qu1bIKdJsJdupcRdXcGb7Ofv6WEI8bHLaa3ge8EtyK
4S+9gM6h2LGckjKTsSkO3RfkjUMSKWTQk8clQSsLWrvQuSPXdRlsY4uMapolkNUgR0DamXJAyP0Z
rcUKLHG7ZOKTrtE+kbyc8a8v711JZjog6wiI/6JbMktgnD8pI1mHrSXBIdBkXKrYNONb/Waaizvr
EL+rfuKtJYeDzLUQL8AyFyI19WoBWqf9nsctR6PL3TbjTYjNphSt58fNVsrLHiWg+hVjmo9dSM2z
aCa8SDGQkM51rvGuEUEOwbieouK/VUoMhQiwP3p9L3ccJNp0mOzwY9XB3BsvVZNiWVPnnTYpg3OT
SuVVRST/r6gDdiT/xDbYrcg0fLPO/+7ca7LG6tzdEnjGSPgnjDRAWx8G75ifeIlhGmjrZeQwq5Wl
Y3rFxOmI1xF9RlitglP0obuCXMWr2qWY+42XAxyr2RnP0wCfuH3r8qDoBHMPmfzvZ4ki13OjbQAN
h0P9AyvZQhhbOxMuI89S6ZBUkI5eeuc5Twpo9UscWC9Dd1Xy9ujhPKY3cQPHaQ+y+p3613YvKB5h
/Kpex7k61vyCZMCYBbrP1QQgh2uBXK4P6yPrHUTnxQlQLYvdx/1o3/SU4Nda2/ykwzJmSrq9UQ+i
t7ZSlcNqVuUvxbErNe9oYbR6xnLt7U5iKMyHlHCXixGKVx0D6Vep/nRzcfAfkepR69O3LpVM5LrA
rTObIDxHkOJYmS0KVvb0GSCfIYmB0vVnbZLYl54Jbj6C73Ktf5/0zDvcDTfXsSxN+HBEtaf211HY
tSr+aJIMjL9yydH+urQXM5ZAZyiKAA3GKgeWa7o2+GkhFqnp68L4d0F6LgjFKf71zenynfsL7Edq
EBFR8cPXpyEx6qAEaRaAPzxeoltsQFQlv6PmH0shY1i6DTmXJOyTLHHF2XfOFTlgChrHkw6UXB2S
5m7kTgcHyrnfRPZi9vkbC9MpU5oaBcIPd+bUqZ2a0xectrd8xmfXHt+ZDnw0EXvMGNZQxWDsdxMs
EjY+axMyYMl+dfL7XGgyyMLN9x9Nt+GY9EP8lL4Bw06vmppexGy+hpXCp0IZmb5rHDUEE3xPy85D
d+F+l3Y3Uf3MLi4SJkcBKfhmAAwoyxj1ahXTqIsdok5ahQb2dI/X4R3Gdubybp6MRFiHzIdnCJse
4FvuvfuFGo0MsqroBj5O4KpWtK2emyeUSWPMWyiD/6/lMIGozzPFzJXS9MOwdNlVx/+uTnrRPwwm
GwcWNvJGJw4Ao3yYXeVtfsGGvShz9wZLStw8TSQIrke2N24DSygrXDN3OMs8JeaiUKUtkXNRyyyK
n/WlCuDsqFpA/EJFAuWg0CECA0HZYKtdPwa81J47zWnDfF9wEiT+1/NrnwN2aR8RDpwsn+/4q8Qh
WXLnsReCKTXgCfcfbMrEEmilssbTmCx0+iV+yDlz+3oAuwxLKAWaVIlG5H5KWkALJfyb2MceQ+FS
W95T2YGDXFuxFABvSLYSb5/KPlzCeZ1YYq3N3MJBmt51zRbz//3JotUuSo0QnayVct22g3i8lyeW
BGhT+du/SwcDlgx2yEL7rrFmapwS4TNJdMRCKXVvQ3IWv9wlix/n60LoBAe4zE8O2dcltrl9glFW
DvpryQXtgH4X/SVwylZ5Muonvi+OuemZMZK9drgXrrzX+qvNxmPrnUdoTswQ2uH6RdydaNBnEjXH
wQk0x+5/aJ99fkcM/VlGTj196TfL0ggvrh3Phz+YPEFaIHSx+eX8bz2kcLhIiU0c7Cmpr3ajOJ5s
dEktj+FIDnRzOamEcLuFI/ks7ahkS1vIQbugow+ZJABzS8Yjtph4pwqAhMMnXgd/IfDL9BoBHwTp
+ql2/PWS+x86Dh76oIgiIdUn992Zsylr/B2KX17Bt23tLskGnGf6TTrztjNzQMNORU8CsMOOxx+3
JVwWNnixz87pMwy6A/woniF5GxHD6yL5QVpnfWLDoLiisE+to1/DuoNJCzaXRpUlsBX6WTsRh8DO
X9/04el5xNIVCv3V0S/646n/6sXhuaenYZzVYI2hFPWflb3f1NadNNfthtmYr8byHmbl6p5idEfu
M1KZuKTHnjOgxHFnauEcCfAkggAvvDovjAkUMkG74BGCXHcOsFk2K7H1HZpdLiI5jJ7LOvq+tnX5
eJVGm6bufKZDAEozrbWNf7luU9jC1ML0lbt3RlHF9GXLJNb3uAgvI9nuSdhEjLrL5rZN7QvIp+ze
fk6yTh9yWA8hFNgIckGZg0auGd/6ZoQXzXs1qATbaCEsaPJTBnxHqJfsqdqnE76N9QZpcL6p0xmB
u5k9FpkEsVjIfOH9mpC7ISzIu7Ujp//1oBPrPQM7xmecJ1JRr8bhvOSpFW/2vKye7zuCL5sjcRxY
P5Y7v7O+dGB6P8QzTz/dfxMBiGxtFvR33avM8LZrPb0RMv+rP5XcDF2V5KSv5I+drQmp9KeskyK6
TRMzeuNKStsK9TX4pP0evuY97R3oiub7Dr6zLthzoEsaaYooYLGWT9+ezWG+2ywCwG+FepyHUmpQ
sq4A2Bri4l2HMqLWZ8XohD9HGNqph+pSn0Kql3+QyoSNt8P8nLU73hvVHS+heEHMVBilI3EC062P
avKFyCPZZTeHmSr2HnRTdVFKpddjpQyFGSVNjkhHMNNLb3FdGnKhEKUbZ2WwCe6NIBSaNMxD0smx
pbpA4gS7tf1ByWZ4VbJZAL93X6rLT50wSNJ3a/ow7YlUkswbq/w0rIaPixTmATn907ydWDkWu2NW
uam3VdNSLEkk2xQUkNTuWn25e8J47DYLUz50Y/rlZBBXDiQk9ZUE78J8vw1vKPvVjyc01//0MrFi
K4YrBwcSI6MuQdKsaxRlDFbQnXSLOFCQRJAD+2hz2YGRKgT9hK6CAoF9bA+oT2RQcS7XmRM3wS/6
oMbZlNC2+1khBiHYVzOuZy9XwKGCEj15C1dFv8LlE8GVbNiWBL0R+IR0TGUEGIBZq3txw2/atw33
CLU+0FQ69C7+IgI4qb6CwoMYuk9yc26HR08V/gLNf+dRxMQqLl2U/5wwo9GRikvDYTFz6oATmH7y
lP3VmoTSTE2PRr+iN/OuK/ub8W4xjMAHU4H4g5hQNWARJ7C7rgI3vEYNtam0FhYgfhB65UFFbKbo
EnwMvznWXebypQf44GsjTmyTkonrmmyYhtPiVbcCvlu15Tbl5VJEiZWzBhZfURg6UBMdXw+09RoE
pGz15P2QigsO2Wcw2A4D9H1i0YdFZ+lFq3oAabBgvbkHSJ9xplm++SLQPYxmsrPZDOn3sUByOpH/
2xIGR2gVbv++L6ooxd3IlIAqBMR9DYZ177oD+v5NiQjxz2BmJSGlN83/o2dmN5U/4o7F3djJnVzw
wrxud8iTgadSLpv9aJJsQIfuo0+y1XPIqmwJolOZRJMcdlqVVGLaA2Wo98Wq2jUZ2A/iFebLQda8
YFRiUPQMEHBvv9yuIaqQBOOcuk70SFW5AL/a7BxF7eoPSS2+FkpO6LlvWJFsxslyZGGtHdNk6VWC
8qiFDRLeK50Z8DVFRn8WcGZ46Xcwo//o38omjNMVwSZUOo0ZSEsDQHEb3u6myVLZMoVrAwoP5eD5
fwCWqqfe0d8iIsEPu3VhgKPfrpnDstJrqLRE5cqDIwYQBIJylJNNJvwOLrZXbqQrii27mFvHUp7m
UVWuyoTaEoy2Um5/38AXwR5Nmf2mGSRKehbb0hBYnppXhraeDUs0HelhGncWhfii6mJlevK9LnCu
q8xu8aWvcRZXtBDTdFXBDiUKbeLnzR64F8zkj8sHWiyPs+H4D/LT1R6tmBYZQBcsXcxdzPGF8UBR
9RaP3NMmFgJm6X2LkIAQV/v/Xo7nWuo5x6WN21kplgn4xOUOHpGPQMd70tl+EocrC16GfFsymgPM
1JsBZdxvAEM6ZVW3CMn3j9N4NeGZaqGDkHKMGD4X0ldd/GygkarfZRTZ061F0z2mRC4ifbWo/cNC
si54dyzMIjM6zAqhSDctR7Mrpqc5kgnKHbvHLZtFDfKrHegMVroYYXOedhNR4WlV07GR3Lrfc1o1
KyXiLOzw3vkn25XqM17n+w3d491ahokk7+x47S4FVLRzF67SB+NHmJSNeT2b7GB1iv+iRpy1CEhB
h3r3IueSc2vVVDGbpKGVkbXi4j3Ox2zeATj/FefkrK1D7RsQqKXV9gNBkBXJ+GrrfDoJS/7D+iTs
Rnf8IHg/C860OftAvkbnnPWEPL2P+jD4l2dwtwj02689rFCh1qO2npU9QnbjKVVHiLbzTorVbM2a
HoUL/6W+yfc8M9Y0tHE2gm9QXb3t2Wnav9VlrdmTEyX6UtnQ3hzhjm4mTjVR12KmuVfD2iy+BIJh
K5/PStSzzVIAUjvP3GbbN6zdHC5+JmH3pNldZCy671VkiO0M1nSyD9QXuHqDGDyDkmH/6+LDNrAU
1oLm/6fwVNxoE1VQ5kdjzp4xRrj87QHr1e1vZJxU7R2H9Q77wxFlHCoJQK7BbEEpFhKwRrOZ4Xu1
ZzYFQLStL6xQ0jHpnPaoH8ypbehOP6T2TlbelC9FGmV3G+o3T0Jg6gJCQcEV2PRF/BqdKIE7FGBb
q9wswUJDFjOsUYnORiBu+yefuCcwTCFKTEnUXZPpqdhSHuoDMKAMwBZIYmFn4GQvLEa6QstKiWmk
h/dKsxGgkeBq8Myb0wdRtEoF4hzq+SyB/xJC9+5cZHs0ZgkrVqsMvuRd7p/xL44i1Q1capFtJDik
9+u1oUsgqAZ2ZZZRtxRFWGIBTpAG8iGXL1eNg8LNng2c3rZmmZVLp5K1f5kI8dsd0F/xAxoKd4rH
oPFw84xvDK7ugObv882XK/SMz2ziK137ZTKiYrfW2A+ymlEdGTBzeLAXSJBgvq3+rdQG68j1Gwln
6pmsrAiakJ8/VHENkXUmYOXMcbqAWGeyHT/I3ddjOx9Gg44FgCTT0vXsD2In2boMkOMBsRPVacTL
1KFslCx9Upp/Yo7UX0E0Ah55JIWPQ3fAYA3WlOlcVwUHa6gUp83TH1eo6FQHXALcxMKSBqKam4Ij
io7T7pSzEyRz7Qpk06DeHqVG4iBRzqr94KG4D1xympyIawTIuv8QmH2EBtVQhqjRHavk7b2wq/hf
Ed3zMdCFmg4SQWmpERxU8qPUXTt8Tir77Cy6yRb9GA5RcwmfnJeUKU3vA59ea++uCx+V5hmx/gra
gxCn44VVC4QAD89n3Yohlq0r/w+FnIh8mK6MujsZpTTjttBI0YGCZpszujdZ1d6Mux3JpHLwimMT
QwhpAbFmjtb0UXPSwHI6ZvYVjegvCEowES2Pra9l0tBckyVyjg8gv/tqfJG5Qb/Sq1xks1SG3hh7
9404vaTzz0D2gI/hzLI5Mn7bTErWLDqnAWGqx3LL0uMKOcnw7YNvddxVvqegGKzOOgC5EjTAExsm
k0lgyTOzK+2vSae6S0vVvIsh0Wiv4U2+bmqmNY+o9O6CgFygvbcMGx/IXg1qLVXKOoSi9NILaESG
jxusA2Ap6YNi6DAPoKqZmN+WLIP/6NnGVrlWJZGb5BldDEtb6X/FAOukuhHo0F29MdHK4/86vmJ8
Z6II/MDFlE5FpzyoSE3hyJ83cMMt5826S+ZqhpYtJuevN0vTXA1Gq97aUKH0+qH9skf0VGUuJG+x
3YeHNaqbfiHRYRM7DQP74FrzTNqRIft9jy1iKpADX0TQ33nwCt99+0zgvBdH56NIdpCQPHfWcM5z
2MSXR02akCzO3VScXQrgg+6jNaC1+8AFB4je6Dx7udHdDFYrTZ0SVbAa6Hw9CGywFE3kphRxIZKs
qRUfFzTdVrxeQAqtCoMcVyODbgfUjB+V2CJ4g7EGqfDpS5engbeoZKOjsCtC0EyN0jciAPiXo03M
rHplK5gPAs/6QoWK3Ibn/FWwFL2GWlpYbUWI37rQ7cCklgxn7Pd2BYzsa8LratfpoGJUFQuFLV93
1QUoaInMeeP/ozOgAexQSqW0oG0LNVXNi8XE09zdStCRgr4tXuiXi5Ir3CSFZ8VK2lanuG+O820s
ShaMmitriaXaaZLuYHhv4dpV+8KXmR7mvX0A/rcWa7dRW2fONjrsmahqkySQeVBwrlEVX2ebOLyK
gilHkhv5RHtjzwQWTCZCG6qL6wTfLjT9YV4TLfLqSvy8XNAgO5GmMeG1eBd3Ub/AsEHCwe1xwjUq
vpdrxcsBVgo/HtrtB+z9mEpTy6mkAFv98Sbr+J+JrQFHIlBjXunFKcQees/D4GH0lzX5Qlmvjb83
ruMoY6hpV8xxCBTapoSkekbCsWIarcxef9AtZFc1je8UXfG+beQ8Ek9eAdL5UPveGhxYqrJxrgq1
R+BSzjofZFcBv6w8UZ9JiymImPBmuBWnl7xaf1ExVelwXR01PH52MD0tbREaK3P62QFYzvIGhLff
WCcKu5qx97Px/mKhEJnBUK9j2g7zNsYPbfxY2FLNBTtobS2ZMcbfK146OENHTJ/QKlvTDEXBTBRq
NcV1M6ZE/T15IY0wozQXL1SgcREVEwPW8n44TOIDt9bREGhYfpL2NoHpCPrOLwf9e/TURFmBP9uJ
A3s7kzcdKF6gZB7HS86OyY7/5L5CpDs3V9ECPfX0Fg6v0TWBUTMwK3851UbbUzmI1Y2jUgry0ckM
CaVSWw1fH0uu1Njlya3BF2Ww3FJfz3FVGonrrhOuVpi9EMtT6QBrabIHUYobjvqNbyko60V4sScW
s+gez7v2RJLdFj3HAsCpV5Nz/zwgOgtdx3/gAPeJGqutmMR/yOwFysRhD0xAMWr1ISVy8XlaSrys
kpk06vEBV8+qDZSki9q8FVxh9dUmb9gxq44QHGn1HimLrRH+lI+lBWhe427buJx7Q7ihP80kgp+y
ft2ohBgAKFvPHhw9s1+LL/LJm3ZRoU5JnyUiLHXYd2MjbtcU8iSpj0ORTteQcNTYg1XQTNBmMyPG
ho/0KX5/4d4aRbK6mYkZrVboA139QMGLsZDLFDDXc84U3h/MvbGxe5HhKznuCgj0w22obnzEPxot
RxzEbtWjhdIxvmPcBqrB+i3Ab7s0rwubBO7ITUonlL/S6xo0tfhX0ZlrpItKePLTF92nLnfB1jyr
fKB6fWMdk4YUEHtSR4ptMIIoeZ9OlGwUonTpQ+7z1AOpz+cyJu3GO7S4j6L85QiGsX8TUBe9KRXB
c1BsmIlg/bEHnW0+ZLJ1XVcSq/cBf3Pw+qrdMOhRV2fCiBnT65iYlOvehPGXRkqagPUisZLj1GdY
AIimVjK8UqjohamObt9v8za4TYPRzSRFvw9DjFiWX581y9F9ew8btdshUiamRytNXXmw6Vc6FkqD
i1495RvtoeeweA3cxCinb8gLVI4aVd9HEbNF/doUdU/hFfdLVpUxwMX5YWBmMDIghcCIq1nbNOFQ
oP/MzWXi5IUFwMZrMQk9C8qIwrSqMapR2lucwKPatwSl7gmuqLY0qorwuyhIy7CtiSYmv1nHhONI
qcdDBAjPzFlknMN3tuVMQOlwO3ZRUfJgbNmxTpevEWcw+JSs2HTwlG1GV0/m+lgq8/HKj4QnPpxS
uVkoX0n70yr4msX6qKP9dbNRA3qigpTf3/QPAcCaaOEWNFVMlmXoyfuixv3tV+frlLHcQ4yD7/JY
YY9rwAh/GLLzkk1RzAM3bFwz6/L7iwf7kUFnfzyrVVIMBNhz67kKO/0pyU8UqgVIKY2sS8iRybpg
cWY1EOl5+2P969vr/GsWxyy8U1J6QFmtJvzPHUZPbGJ9Ntrc3BsH0jNfQS4bZ8qWJC2KIUdCJ6yj
8OBofs0g6PNDNlMUiJwXCNhqW7EG4m5pOm/zU5GTnLCOYK+UNshjhzbsAbxH6mgpz+DHYw+ijtr3
wPt/WFAEHifIqsc2VS+/aorRNgPQuV1HrLsDPwmsgg/vUzGqQpA2xCD+zZmeyrsQ8gsl2wX3mA2e
Rm3KzECKHZ44BQvMu3KQk04gz+Vt47h4z1fUOL2iiosnIE6YWs6rrstm96mDqKP63hDp9gzuni4b
HvxEytaeuaz8PtY19UR6LLatkVGPzG8r13ATPdzjeMVdmqdrJiENI36AaCprDYDtyO8D+kvGio1M
/nWHvTyt4s7E+CISjsfhLFPuaxt2QIroVLZVsFxjK5pQEnZrLQpoK4OSvdvi3A+xNrX3RNovSKnA
e5zpZDi8UEkbbvxxdVitQ08AzitfmKVT2LKmyf5x0YKVY9f/riMbqdst6IWQVvmXZYIilsOfK2rI
NCBp7UtY92wDobmn71l/YWjW8lq+Fi8ijyZ5Bcqf7T4BRA7OvpIu2TqLa1lZiMKKoU9DwBax0FMz
Qf9risViA0U+VI0z5R9ie54VSW7nb9LFXfTKH22QA5xfIU0Q+PZrBr49c7eG7JnShl7dmLUtfnBy
rieZc3wQFYirkjp2Buu03ZuQUziYJN9JpIPJaRHgDOV+MrZX1aZjBjlXdpiTD1Vt9XuJIr4Q/1jl
l0j2wKKXbOXfFVGaYireG2e3B6bRjMbP3ExC+7+TWO10LeYv7kMOvzQlW8BBqUC3wXgaGDBGxrCP
NqhCiIeIik3lsFIdnLTCoW/daLz1oq/NNNUH7gfpxNuVXaEvAJfx2RQImz7hOBy87xScpMZvSXyz
6t9vyPejUj5qf7orIpytavAtIImjXt4POci9fHzAB0UogjZccDuNR7wwovEn2tSiCHX7T/FsKdlo
LF5GpuzETn04kD58cmzQrrvzktdN0/xgGHd+oA8qsJjj9wOZg0GOl4xfwmLRstiFMZkBTZednGbh
+fevTJZT9mlJnhsUkOZJC+F67QGXKL6bNBo9vU7LQ/vZ3SXB3+Q6F7J4qGrhsnL+UzeyIOUsZ2mK
Qi8WRUEdlwngWZEmJlpybBPOHiYhVZ2RR/dj7HS0lEPRpa60ZjGVulo6HMQa699XGRv/S9t3DHtJ
jvELlXMqyxwdtkRFXFOoP3sVuShGQ8E/rDQ21DLxFWauc5xHh2VCAMceHyHKsDs8T2qck+o+suWj
ouobZGrF3xLPnxjrlnhBClmGHSvGKSSHbUjsehGnt6N7NqDLrepy2nK09XhlA1jXQSJeWIwQarOB
YON9RszvuBBQW05NGDUfdYY2LIGkjYgyyb+cYxj6CYOIcT6ehbJEvQXZhUP1ly3CLgDLQeCUMWrT
7Q295gfLzpdRE756U51zXY0NHyvZ+QV+OVwJoMlUzvbuGY7WVe4ki5ZjG0H9rpN3XPCCVL5FJysE
GwZ81xb7650kRTjlA0KlbCMNOlUNVrn49f5U9kJseZ+3kZbIYh9cX4uAYKGQFWKnw7c5nUiRe+A8
5z15J+lcxuMjJOhShnW/xbcoNWxQ9vU8d4ss713+iI2xe5YeFYr595VD5RXAI/PZVti2lZzzxz+j
JSQhVac/YbRaR87Ol+RJDVqxBKzada1m/5C9s0XRAWZz0KvoPQOkpk1Ot+OAQT6boc0CPEqdVHfN
LrPqmI7qInOxvsbbERAa9+tduROf+ETzbhZCbN3lcCSfJS1Lqdb6poV8kLvTu1xB1+92N6kwkC+4
ZSM51mTB5jM6tLyby3FPBXzSLLXHCgRFZMjevB8JrC6KzpkWCm30cokfJOEIYNw12sqObCDwEakB
Do/leaj1sL4RbiwLXHj6s7qO2Xra0Eg01PUaFIbpqOpNyN1vMOL8lTpAd0DnyttNtG8ewV4lh0Re
vtVAR2mIL2dkyOZjNaRSNqHKOEVnOM882W//P58EzrHTHRfKDIyuLTqYU2LUWJcPN2DVzRYFQ7mY
7J8vv1i08+lMjQKQR1MhR4h2KqUxrU7O5eQiSpvZriwe1WIHVb+29Zyh60TDRUTRKRjioD7+vj+t
oSmJryiHVw+4/WzOzX7OcWU8nqIjXvi01Hcs677o7TOigNqeZrX/KdVgUIaxX+rvjvn5ei+cuZYU
gvTZHBDpPSG4T5/ZmejjKs/2fblQ5Yoxo0BsmFxkZLHvZH5NTChBQX/e+HsvP00s4SMfryxKXr5H
bKxn3VVVh2DB08glr7LY5f6OG7WIGoWc0ehggnETAzkuqdOuxXZAEXyMC1BbHtj4KU5K2Wnkjq9T
hfabR1VhoUcqngunWZN4zbbtVOLnNixkg8l0tk83hOyDdS0U/DyNgsdZkLFUOeRKQ8LW9y9KCM6W
koowz8bX9cJ97SCO81U8wXsMo/yj6UaU5diFC3odsh7NhJ2znlxfzOSh0drDdKwhK6OHbR7ix6IP
PgHDWyjZdk8++NMgEqvfzBs7e2RDcRD+CNriTtAtqv4oSW8Dw2QiRtjA5HmlE95nivi8OgXze9B3
QZNapxjlOpxkEPoh/xEw52Eyx7oEaPpqjIC55C7YkH0yN2sq0Ls7SBvVs2AlCcxfKe/DOqemZcTb
QrqrGuwdn/IZc1zRy1BNTM8Nfa90k6UagYMKVrkrob74m+X+9ZOiEEQopYKQMBeTd6kHxn4Z9f1H
vQpWaqLBGF3rP3dQX2MOkoyR442jaH5cOa/ciVJmV3LoyHhS+tpYbu1elUyzI3YAV/l9cMpgz5xo
vJnuKrq3EIYu1E9surNCStkSWYhE43xJbnIIQAhUObGKEFjb/9tkXFm+GY1IsMsPLmhPzfAZ8II0
x1+jUDtjJfUPx7uzLD/GyJ5NGZpI5qwKzC5o1jxZR063ukGNt+62lqdN2CmlWr40papnFnAXWo8V
LnGf9nY6sZEigMbF7OtWCiU2nEj0zp+x3USG+ZE+8/R6ibxV/J0O6iLvFDwaW6FILH87fTO6Aekm
QM1m6Nu8PFBwlzKXqExw2uPfL+Se6F4VPq9UnsbAE2XE+oNM42rwts/xdILwkrL2Rh1aVR5mIZxe
B9RJe2IgD1d4ebmrfS2kdbdbwBys0mwkw6NZMG+eXU5iQKEsQmjIXcAj5/lI6JwInnEPJUPMl6Ls
2Sbz+9/SrZPsQmWipe+MNNdOaOrZxul9Ddhb7zkm+Bf+ASTd1C3KC/kFFzrunzw040Rato95lAu0
p87Dy0PPu3+h2AJpsfwRzIwuIPgPQhla1T8cHec9r4Yldm3UcsRqFo2NieHoEsU9L0xbD7fmzATe
VASBrWzp1T03Gpu+EFAuooj2LV84VuvgYumPPcZnctCi9vDbm0ePh8pvfeDvOmAk3/Exv7CYkIsf
g/myDYiupmFVFMzME/aSTkONU9fgmJtgLnI/juPQ8M0yKoNmwm/nfyDw22mXDpG6KINVhSWuBwoU
BWLPdzYJFZdg+Y6o3+hIHZkuLIIDsoYPxGAK4TSbO3JdEKQoFDFB/9BNlW9mDDPExwpOYb7N14ug
36KEUqKbwHxjgowqYWDSQvNXtxd9N29d2Vg4G7sSwY9AFmOXgNwzWWzKQlFXsL2t64NX22lUG2cF
NfuR5mtWn92vFLeERN19fZjxrv6Gmv0EgH1eTA/ERDJUF29rnGIAICZyjppPWABywBH1oKQN+0mJ
bOCMoAvnDmL/Bwmrs6mdF9dfU+mvNN0LUYxlwSzo1bZhHLM0AIAJUOfTdn4UHCh00wVTEuflWjRB
7dPBG1FazDmoNLm2uFsttrkI13ZRXN/UDsfCWAitGrUppTwvOIeAR5dzdh5xv6YB+6ov8N1kHDy1
eRPf44R0cpFL5ARa5mzHhxTdti9dvTUR4LiE0DyCD5nK4r8xymajKq2+hTje69tFHWSqhvPh8Ha1
IsYA40GRipR+hwoDHlhAgdWSTdVBJJBc/XTI01VMbBlarxuD53jkvGBqK3J91rR/Ga+dF3x2J0DG
t0L4z0wQrE0lX/MOu+QYRY7B/PB9n853MXxnpe0C/pP1Z9FPYZnK+ZYd6payEfJay1mWuklJLZMn
9k6ARJj9zPQe5P6xSMTd2eP4S8agVawxVm2CiEwXnkpGQE7X5Z4aqiKHVzwLpq68PULQnYDoSXMW
+2l0RZ+qlHIGr7App4YFvL14725OGwjWOViB0Xh7xJBl+DV10XzfHb8jXoHER61W5C7aCx2vz21d
Ha0/N1uSUQmrVVNATp5LWBm+q4T/ABCc/+2uvMlcIzF1xv1i9lOvSpkDp6uTvZQWY4Ey1Ts+/Uvt
z7BC5IBljXK3Fgytj4K+7p+srfZ75YJpQN/UV0Td1+nc6Tn5ueQ7QfNoHZ2h9S4xOTFC7FaUfmju
QT+ZV59hUFBuquNAQ+OrOPJ1iw3eg5TzeUpCarIGzxj8Eo3a8+PuW8uVDtGCqEjDlVXdBF6xjeEn
UFSWmhDu+CIwuaac34CTo6qCBdbmbOoUAcNDlJEw+Ppe33iCsFXRwdXAJwebdBEbvdxFeqLZVfsQ
76cw2VWzVKiRnI0udgcGcUuw6IxHsfp0k14QAyF3SZzqqBKr5ze89QsOfGS59n4+7Z2so7szprjs
Q5EfSXNkgci4Y1XBbQwoW5EwxMNB9El7+k/x7h7Vn5rlmRtW46oNmCAUleW/l3rQOBehW8SQhu5D
wlc19z/SM6oecHnxSeRSOtaxIn7lfdHRwNz09qdRL1gJD0ZGbYw/THH6Hf4x4758ppV7AK6ZQHoK
vF6jhZKZw6O3DC5JvP4adNxiDO0hfKrasgbO7pRvMcD07w6CM6smqD88pXF5dC7VWuq08SZSqErL
05g8JeV/dgmEK3Jx8wU0VOe4TNmkFkGqD4tBtXFEMtTW+xG74WhTyPnruyc9HIXndIXsS+TBp7hD
iCZdgh7f56mHSZgxipgtQ+98+vPJNRQduRm18cdGHZs/iMLaMj55qP+ZLeeMDh4RVQ0iqRXSjFYS
PH8k/rD1EZcWO4bMuLXmdTVKd6hA3Jm0PZ4eT36gG50vyX5W8KMmd11JS0kAavw6XJqj4s3D/nAR
e6q7M72EmB1M8S3quLnDMPfOXTu9BNAUa+wjKwhH3+ix/rZU8glFvPx0FjVS30g6IaUC4r9+GAgY
RQsS+Etd2hDXgdyebqSjdtapvws5ve14qiYlBD57h3JOFXN7PIk7bsWaqh+3OZmPHGd2e5YaaiCx
06IlL1gNW75DNJczOYz+nFp/voOCfrYtQ0uIOk/WBdqnMrSmjgF024fy5C+o/Tqy6FbWLPtGrP3B
vfIL7hjO1Rk7N/BaNIYIAeB+o2msTCyanbtbcoVXdn9+z2fWLnXCvOxIcauWQfdYs7dk2IV2SkTJ
iLBFytezvwkMNMFDkM/3MnIxKAzvwUxSe9z7q5gWP7VHcbg1wwtwAyo184T+Ild9JnODWcFm6w1o
bxE04SwtDCS1b8WAUQ26cUcCVkKJngt30+jfPS/jubm21268DT8RYn+I7iuACp1gQPS5/RWGVvwi
Ql7V+cleerDKozyZ5vp/dZXNbXIN5as3OHqBGUKwrl0njoojmMwNBqzJ9hOb8C379juT7tvl9/M/
au3MMff4nUPWhnIyt9Db8aa3R4RkOykdmD5pKiBotDR1D+53gFbmSgs+39vE7C3uHGIYTsGSJvP0
qxWG+SQ4PrqjEug8ano0R0ImbXnLqUG4GiaZHWCgZmkAT30s2HKZVKCR7f9NLBi4SZIg8g7m4oUv
9xGasFXYt2EQIDn4WTBSEZc6xvbufCJW3T2pTY7xz5hgDgq2CwhVzWVueyRDktSfPh+QNO06158D
HGFQjBbE10AgxDVWYPp+IDDGHuV4aUMlRNQy31Y7qK9REjFR1/Pigqao+t4X8FKmRPNMlxtI7zSI
TebMTKOsGkcBUAujYVSJAaLVJKXPf+zVUfidXr8FmZyFBU5r4AmnOa4OnLcOWagH2hxXr9gShpGP
v1vkTJqj1o9vUJl3AXgKDoZDPaAcbvVAABL6XyVCOJmQVlF7bt3nklIQIpEiPqJg9nRMowMdZJeA
GToNgfNI+XBhfXAEeIRzn1H+l+zZXkR4f/fOuqyRmZi+acJAFe+8ScLEqlgp3qd0+ckSS6SVbA4H
MD1Yc7c/O3LbuRm8JzJIyPm8fqLJNC2C3DXoLgJKUkkY7uZAjBBq/e0kheYeLj5lx9dEtmCxo5ml
BIAYrQxhQCuWn+tfGSKQIINQYrtQWP14/8xQHUKNzLjTE93/LahtUeKS/U9/ni3Q83GZeWMSFZoR
akIwi9oeyKvBC6019siSCCm4e4aRITZjvBeQ2jOiStFq3K+4gmUPbQoxGjTLtwibBTBaSsskgG/U
p71r7ABJe+bIMIkMqP4JI2Zl2KyQ7kVtd4FDB8DeEi9V0QtGgoJJkHHfi1nA3juheApvwtbEgwjF
oGTdtInBQgfvZ9oxGL6+GxvXQx0gso3WIgeT4qxrfCEsaLqEml9kY7ZoCa/TbwFOM4KKb80O4EQx
z/MeXVOn/Wev/FojXmXYkQoLdoLQJyLRMZqsDcYq1e8aYye0O77zHbG8VQ+iBM8Lz7Ct5FPd4Kzg
j3ylIxdKY6jA1+HDLE+JLyj05FCSNOVwQXUKJiKqMNvFDLU6F04oqUotGOBdToj+Ct77mPNB1ZFV
PxmX9/rMCgxHYJA2tpzXsVetGASuCo6o59cN0TBRo1fcYhA3ubWMpx/VbB6ISzBW10q8YjAdnA+I
qRNT3Z0XHQKZvLFoz11CBpC69bYTd4ykJhBj8ios2Wk7nrBgFjSFhKbtrjCUBtima0mn+6nM5mDu
I3b625QID0Y581UMrpCs8PxEuCRsEE3y4kKFY7LFXId3x1ABMjcKl0g5MgTST3Lef3XELCFVMgRv
xdpUTMO+TGbHMmA0EznmZcZW0FOIZIC+FZn37H+ypOzMbN0sLYuAEyU2MeYaACMV2qXq8nQWLazG
i+fntpzV6JheOebgT+buCAebZvv80bn7c0LDqRbWcucEwIWG/Afscc85JvkK5JPXw5PKUpSnEpRm
MLxan2oEsXzvpMAD22//RPk0bwUpbNFjonM8UgckKhHfSLNAvbh847hjDnbN7Tj6uU1IElMyEa+i
Do7TcptMoU46ihbVOzreJd+VhxtHCQDIkOgSRM+dDHtxs2IHH7SvpxZJMZu4lBaNyYD7bezkDnZo
Y0e/cQdCrSQtXrPAVXZFPlG0ftLs8HOOi/tlNC0/2KFYInAk3pFt2uUl+NB+tF3QoedKV35AtE9a
CgOz5j1cLQr1byT03fLWv1ucz4E6UE40EqRQe2LgEQKzAHPvENH9t0btchVLjo2BiObRr4iGzsD1
PE0zwok0wdTiCHEns8yZU0B7uipBrSO5vNeW9+fdbtM6um/uYOrvRzT62nGNy909v+V9n6hYGc/e
JdomgJ8+DdmBygZJJib0UtM/VU5cs+GQtRc31eBOYiOS8g7A8jULpfKdlyAUmNOPXn7+zI0l2bQ0
sxVBBWtXQnGYb2DhjGXOC4enD8BdaNo7LkheShXvYmCxHvojIAPDLkou4SEESAKhXiwsbU3XSUUk
JlNOyaVwhv32S/qchxMMxexqgg9qf9tmtOl1UQWVHGEyA7qCAVb1MLoDyyY1d+Q+kdndcLDD5ZL4
td7W2UBxumx8Hy/yNnodLug21/LHBGlg0uFzwLmuOO95ghUqij3MqwfvkSeRb4ws39114+UixRt4
JyFd77KaY/TfN/h6iyaxlpNrbnbEI6YcdTeArHHETL1UThDpDSvtL13kjaMCzta+XC32VVXLCep1
MC1Fsjuym6uTw077xP03JQS/1Py4Kgn5PVx1AeT9j1o6rAZPTkklO2gBJLBBaTTFkCiWXZW7qGJY
Ex/gatIvZMOkt4ItgHkaBBm5RKgrf5j52OKDDfnNHabcjY/i0qGi3JUmJu1AfkcFdK/zvEBCVZDL
IMe58k6otAHLFfh93G7Yt/E6oPERtPkhKqVLS152rjDFSVpydUso2VD79o73j/CkJjFwlBBGQDZM
xLxkpUWGwCF13NE77VzxdjYkEdbE9MqRWSCLR9d3rh77r5FlSidO9kU856jLaEDHKd/FYK0q1Urv
SPRyReI60SzYFPctJOmtyj0WK9KNjhPqnwcJ84pWYYwWP9oo5xOd6+8PqLaRDN4sSC/pQLOMAl4r
q2uqHWMruYeQdY5dW/1VYo+Du6guQnU/4Xp6TX8ECHG4LB+BuRF+uTnLqMyq5qqQthbGxyOsN6f7
TPEzxqmVg+pk8jezOwtgy/ZkHr6Bw6Zdjbqj3xZaTT8zMMlRaz8lBfdtYGw/0nWXYC8NLlLj/iXI
xI/gDAZRtMTeWFCpzaQ7Pj8XGJifnjhNb8BXB9/zV96/P2XTeJTbNe+obEbFyfvjj75pbPPpu8xp
MmmfbJ4y4XG9Zc4DCuYX4kWCE1xo7XqkA85B9nz9jau1PKBKbN0j9+KPCLCxvBgHsfOom8vpQ0UY
Vm0WuIYTdXxJq+dqjGLq2G6qslgS+myividJtPQzUIc2o6iinlApCNQuHrEHIJiyD4fz+3vYjVqx
EPuODGR10oByvisEKxQzLXnXf8fyxqba4Za8Ng9m45f/qdJuyaTr97/obJ8HRTmEyqXzP62mpbWu
m04CtB3yZJazXA4ZkvTZUaL9cQIBhrdCesQdgSvXxlnlJrV5+aM2TipJbzyOPwC5MOFUxWCSKdID
/N8f7qC1uNvfsLgT9rEQ13DqdyQq+ACe34TpFR9UeyAME5OFvs1L0TzO8AxS8AakgYhuW2DCInkD
ZVfHy2kdUybULEMJXRt+LadFc3C/Sjp4u50d++TAq3YZ5qCMkefOXxdtIojyiOclMoMm1AMvDGC1
MFcCDWBPYm+SsS6XufArA3vYbFFKwlCUIkC+5zy8YpjvJzf5sdoyaDm1JCHyxaIW64gMTnl9hvny
QWMt9UfaYUmuhl90WeyWBVA2q06J0l/DlRozqaL3gRCUsHsYbccngKxO3cwQB5zSUNvakYl/82MG
+P4xZLqWpKmllvfdDtSYpQ2s60dVXr6rF1RAFS+NHM7mWKkbRpQRtLRKBZGjBey17vKfxWrcoyhe
kDTBuBI1Vw1JU2xQZ+UzVm7fcICXi8B7qE85Xgaq5kv71AcBkoVOJ8za2eKaba+T7PqCHaQL6s7G
pJ1g2ajNB1PFe5z56obksqUPOvN7H0+QLJ1fVLEl8HpiqcK8w2pxjstfJMAPA/8nS2Yd9ILFIi1G
xCTYnqTLpbj/O+9PcUH4qM4kq3xJRdCxBqL9cWaiX0+zP9jkPQQTnYQ3SNxKgwJHfFo27JbCzDsR
hyIl3rPrGrLtCIsk1gyCnImrVTdEXjHbhj7TggbwxvZ3YHbZ2q0D+n9vVqeTgcuf2KAYJPgDy6Gm
9qc4GkIov75Vk7KJLcqo9zBfsY2Wuhdwh5t7s2UhtsBPotLZG0hmeH+eeYKoPR5x8Ljjem8r46jL
Z4WUsyn51Tk7+6JYrLtal4Nx/9NBaozY3FjXjTRGNYxgBCT8TIRYdWFKA8/mpi8abiiIrn8XI+tB
xknpnmO6rplYhvPvDTpU3bZo2aMCG5JpR37DFCwys07pE5MUoZtVbwVSt87S1uXNjBcocKfgvIIl
GKvKdMG9iG/MaFDM2ssSavvxV+hPvZt6Ve4nyCfzxhGFlPBWMJUlwlBSrR8REEo5nF/fD8ynEou6
GpKGBoV2y1KyyM+tPfO7yY8ff5iKkt7yIedsFKTcVfr16uC+2Pm1LYY8H224BEr8oEovLf5w79zo
gi31xktPJLqF0JpXFGB7qYI6vGmyes1fy5BL2c25uBqUCeak8WonNHXqDrxWYlBaBRJQzMtRiztI
/kV+GN4ktjSYhS/IMUWsQFBByLOaBSHM5WJhtrxEw43u+RiQEtNxeBBPhOzdFLGdWz6xeb1U7GVD
6NKJKAp5+NoR3cOhgF00Fa8LwTs5Irsbk1nWb1BAcBDs452N2gnWG+zw3rrMoi7s0+NwDKdbpUIH
NlkWYQHRUZbuWkuRhR8nI3nFdfech8/KyBnVJW6hWW9wmbTVU6WenrQZCURsEIg44LjPwNuFX+ac
UkhHfga9n8U9r7x8DSQVNyf6Bfxkkc8f3djyZYZ07M6Ys7HE9Kbdq1FI1qF8dH3y3w8J6t1/zEh2
8wIAsx+G28d9fF50U7c5zDXJWoQy9QMYLQPYFX7BOZj/TA4MqVTrsBmrbbaKW2RK8b04IJSDc/wP
3/0Wm7ggO55cfM6pfMbBkD3sRwtMbiYT8gayjramUE249mnz4zRNw+OkUsm5SIyGe/6JAdkBOTkG
Y7tqNbmG+q/j6qOykVvr6a+qT/hirdxFIcge4BAf8UQRZkhbIdtztmzN9tAchvWo/Kyw2v9SzB+I
oXLQabkHUs0JKZ5nB/4oSMF2hhkabFNP1aNnjY7gzdKp2rja76ZFBib7PrixNFxBdV/dnwYyA5u1
BMnarh4TaZ9VUkRw3LAmNkyeOHiSnVVxFecp7GOxXCe02vD5QAXHQXyCGwXYXCuX2pxJN4HRD65u
ZQcCw+hleirj5z6VK8IttxdJRbidkJFK4whQ+r9ZyFj58mGEbxNrKbNbeyKzCOuoumYBE+VtzYVu
JlcELchRQthwNGsOTZC3k3IXAAGBqWucIb5Nkb3ikQA7uedAysdXOMxqzwrnEFIM22mvZ/IlTpjm
Xjx6BBAE9fyvhYZbPycu+TmsSfAEgu4zYHX7nRI8pjxQ67fiIJcPA/7uVp5ejm780fF/sD68KuVa
yhc5HIuLjp/eNI2Bi4X/kK/ReOUrIbf22OLcobWZdFCL70g3QYtPOzim18udPxXxsjdirPtTaPA9
9lVfF5Jo4N0N2VVY3ocHHNQNBeMzGEa12Cq6ipsOzBk4l9yRtH71f3lzqu3RgrhCO5mkzDYEa8gQ
c/q2hGjaiB72PXb4kDm422OeTYxjXu0q9QhQ4NzslS5sOvUb2ZRfnVHnTyJcrIdA5j8bXX9y3z9J
ehCgb3vLxUBMfoCkJEW57EHdvbk5HveQ6xuL8c2g9E2ZV3Kw2/TJWE1xg98xn6l3BaZ/Iel5E/52
wCvQWC9FZTB/IBqSFmIamUJalLriAvdDTnoz95C2sVQfKRASAXqUuB/d5S2tW5RAuBBvWtcJ1XNl
el1pcWm0cscBfSBTUwQSo4i7XvMI6T+F7JRfm9ZOoIgnxnJkmenm3osZMtjFltpyCMWAX3rmNmOC
oEcikhy0M4sIL6wrzWK8UhKLgJNDRuyCmXA+lOtvUw51r9PrC3rhc5gj6wF4A6X94+utXeVIlFhw
vAwKopW/1H5CFLQEyt/q37ElIvP8q5+MqKPL9K9VOTRt5aItYBXOHCfdnKw+K0CZEFSvXkPCmlDc
6mAnZBMSow2tFOvaqKbh5oY6aVQkO49GkjDwvu1a+msJSn+gcZFkyctrs/RJse1KQcWFSg9hySSR
rFoHXBKlnqOm9BY11rDRnmWn0frrH9qRy1PCTQ3DhZ48D9XHuHAARU/lvTvnazY90fqk/R4fOGrt
o0i4HQlzaQtw2f4Q7YKm0YPLaOI0JPfI4kadF3PXhl8bk/Cl0kybwUrpK/54wvqioX2SYP7jR+IK
j1VfQDsc1R8Enc0MCq7ATjtJsC9w0PExMg9ZPPgVy+X69iKYGUOfe68CQ4hbBUAkz3tSR7DMFdMS
8EdWqLg8ssvrET+LGP/foMsTA+jAKimzM63JSZcyDQhDh8DhCPYUn/YPeqVzJUa9Qo8Qrasp1Vsh
OpI44CbAnbhVz9QRYAzGRUYveBb+rpWF8iY3m7syuAHkKMgSwNsEXlf9+iqrkQv7XZ/+CGoflswy
JMo7KvbciG+xU7c5BH9bhbJXQfrgWxZHInX7uBPkFVxCf//35VmR/5KKfzPY6nuhAztTgbW2B2g1
W9OjfhNxEKvPzspozy9IfYl0iv48cI8DLut3v/4dbN0nVsU7Pim01CogEyB3ErX7JvDZG3gqyLaH
6h0yBQ9Mlf1uFOKxR2OW0ZSz+pgEsCY/nQcS2wnCHjsMp8bM2Kb9mY81nZnA8LrviNVvF/80eVct
Tngm7PIqoY3e3z3kOaEnr8ExHPNiJyFv46BCp0pIDJUUfFssPIgtBMmSKFJRw89xFr2CRrgew/EL
ix6bUwDL8KQMYT3aBWxw+ygLL313dRB4wXN1JlFVIegeFJg4t47Q82JqEoEdr7h0v8NAJ9hJykbT
uFdJwK+zTfeHJf8stLvHmCyWVhxrqEaqCXc9DWxy+RUqOQMXpzpckK+s5GeBkagBF3xIV4w6vhr9
fZ15UThfQdu0jlGVIoFclr13PJ7IESpGsJs9UnT6uqCrWtfI0Omv7y641T5BPM4qCNkTItzUeULH
sALKdnRGhbSmYMBUU8Ii1qeV9h7q4tPo2xLBZPnnL79XTTuRotjMXFj2r7U8wHfrB0+EJ6DS99Pb
sMXvI47xb5dLNXeznQanGn0sWQblQQ32v/qCzoyJBTR6R6sSDNUPQf5L5BuTb/KSQjqtPB+vx93y
RrfRj1yYCKB7ZOHnaeIWvFurPNmJoY9f3cWc8DwCWIe/zlitVEgsVDVmv3035FDa4WxRsf3fHynO
nWZceNg8zKiiGBu3s0C48+0UJrPtRwGFkacv2V0Q7UIpwgZuPTbnr15n3UUCmsYRNvLTUUfJuCRQ
W/ZUUs+jtgpf1m7G/ZMBjwGvl48Yu1NvWz0OagcXhBnIQ33+Jcc+kGUACUMp2H8kYb++UPXtnjcK
2ei+XJoyCrb19Ew0bRQQBpW/gF0gbTkwVzNpyazCxFZi4K9iwyHmsjRgSLSc1V1vlv48EHb28IB0
DxVjZbj9xKh6eSXHI4NR9D5P3arCwgCMizuj7qKIcmLSo9FCl1P4GeipR1UiZjq+8hY4m3r4JJxE
IGq4RhUkTbbs5ClkhF9NTJLTT9YCOABmghuKeEvbi09x7gxQ8/YJB83PpjlEGQYo2sWYg2U0q0oS
pmv1caxGjenlYkgpLCFlxBQA861Rmu09O7SyzSObOBymaX6cYsxL+nuZcJbZvjg+RSuFMrIXWAtp
X1jOn0GeRLr+/1vb8yRZbnw8MLU0jO0YnUwjU1rs29OBvo7ih7ggdxp2/b8paL1x9nRAo48eHI4v
FwDxeM9gDhHFkM3Uw1BKLT3fmPXfp7m2N3crHFEuaVZ2g7mGm0MAicQ8PDevyiBXHZsC4IuHc1Uy
ZklyTVEW0UdoYjaNjnzmVRpcORQXD/4ofETifAL+LIuzmVDj3+pp3LcZ2Xqb1ZFcXhtSBx3xtk5K
JcWEPpH1AlaTBxVIzzkS+T7w1ZxFrAtUyAr06AAqSeaOPjebJYvZaHF9eDsZOhOdAiUkMLybGMOt
6K7NwFRi4j4g8i2il6NF+SfmF7k+uic6loIi5NNlNR0oEc3dmPstw78NysIhbafa+B65c8cyAjSK
AQv3FuHQq24yQ7KBYWSJgMdPHII7WTWDgQcvs6VBBLqjM5oJ3PjE4N74Y06s+QoNOTy4KSpcCrIM
5LtP3wSmMngNt8VaU1U/iPkAkL4gBWaqv/cqD5o+SEBXVQOvlne3rzLhQJImSI5xhH7jEVlGZ33v
5uicnRStjDSEKRIGcLDp39/fuOvj+aRBrGfuK+MbmnptnNeyre+xtTB1CmSXYeX1kr9zTuMAxBzb
AFMtF7Zj+0+EEgfLGAi7NiU9oWtRc39nlc0DvjdgltNhrPIIOCAehFjW7ylekq3vnC7gqBu4HhsC
+QtmdkHfRukwJeHX55NBXb7UN+R/xTkv0C2DiUUnI+200pwO31+QDplNtvbQ/7HJ7Fxv5CVkos0I
8ipBrUY+hV+q8qPwYF3tdp/78v2LV4z6SK05Uah4JEIWy73X6MRlq4KMhqAu7dLd6BilvaPE0sdI
HYlB612jeiULRfOUHCtdIl6mcNiRxHvPHnnM3F4EpwZEf4y91JdSTR7eNBPftl7Y32Ei/VuEjw/h
zv5e76+YSoJDvinfzuVSZkv/iwuTSmYHv3tpWmQURmxJh+Ok2L2joUrKTHp204HIdDWQiWwmTfJ9
7hcxzHVgFkdqtp5KUbORbQh8Ya75AvGcXE5cXnPcOnlIud5iDzTcmXya9VcUZyH9sY+9ScN7IEmH
Trt9TZg4J22D4KcKoLzGdeZs+1lkAjfDmiLts6pQIsWgaxqUClwVQ/ZVThpSODRHyqBRCAChYHDz
mqck+IOh5cM6h4gxUugTZmUR0MxUaXN/pdCSoRsndSojhmDkHn7AF61km2XKnlRmgUZne1iDjWcL
DdADDoYraiHHoDooRxbssnyA8aQKH1cbGK270hdGN79CbXjFW3himSci8EF+0YF1b7OHMTpVmenF
99mKUiQ/33lz7XWEkYshXzo/W3JZdi7hNMpyaZFTpafcbk6kpyUfj5sItL60TMyqGh9Ht0A8bTdM
xW7DlOxz1S3BoJxgOOOCd7ohGZmUXntXP595mvVg1vkMIdQZ9skbI5aB2o96wpfatDD+Vr8TG9fZ
S2fIFVDZbB9RSIloXdV3fGuASPQE/8uUIFw1QDlFyOKnH4sUwtX3wzAsL6I4q2+xv6IK/+C1cUDg
8JFtkXrO4+1sRR2O2cRed/fv6bkCRSVapeqweRaV5csJ7cd4/4f8Oggn+hDPwCzDQop6UbEjYnI9
gB2YDe2PCLRAvr6WL+S7bwmu8rRr5c1+8jidf5IjxtIESs/FjyErj9BLW+hlc2k6q+s1tnzmZ3re
xhrEFu7i9JII2zy17vH/Ad+CGkD971BiXcqE5ieMarYgW7cSv8YMjnYm0jD+ryuT33aXuNT5/0c3
3blhoxn1BL1lVtRsZSZOVTYC+EwwdiV7eyLzL2qRKFdyqYH/ZWeiCVAnxpFRRKuEzToEXGAtjcP7
tzeGloDWW+GZky8j12UL/B5aNBvWWUEo296eHB0zhXjo3644f4+Jy6+9iDi1/H4jMiUsW74ZXdrn
ceYMYDxg4DJNUjwnQhpUak2f+SKEwyFFlFbq4p5knIr0JG51tsI8mtjV8hYLToWaqvEiL700/Y0U
j/jAQF6oRfoFtw5QMkzI5Jh/bUssRaLSeo/th5UJhLSHbZrKIff0M5YK9EVQKH2RJ9Nva9zvDXa0
HVxyIDLToulx97izaUQGUZEOZKO8LWvvpY2j5DEDJ/YJ2E/zQ/2ZGZ8nDIJnfsPgpq+QsyW0T/kU
5LMr5UPQGXIfLfB+7R8kmXDm9RKluNhXJNngvLDC50c3havP3aeltjTWPTjra4AOrDGEVKzrqnxA
nIbbaRxRfvhztC5Xp3kcfAOiFMMzZhOiynqYivnoJr+PPwpJ8Cc4yaI1n8tpr+Mhl46/aEyeDDgD
zRzKKZTwywt9jyFzCdwsEtB+zKoxAADNJBmjM7Z3XVYo9OlJS8JGdWxEVkrcHKw47RDjbfnPbBUr
1SZXo+oc/yju2ELkY+RSnz0V8FKNRNFSxXLore+kDanNmBUenfNR8eMsRuorSQLcNdWMszx92NeU
moi6lPbc8XG6pnUzsE4bQdpRX5dkeSl/FnxOi9R6Y7uvLCWYigjcVZzByqlnkAwl7s+1AYqjn3Zp
6nI5TpU76TxSRCFIseTzARoJfiMO7h7wd7vCpEYYxNsFj/t3OHXJ6TveGrvruw6Gyizi7OPfEqSV
+tA2WMUzojS4HDzzJNT/nAbpEUDxcWOHADT+bKnYVE1HPs266Uhhwx9Bt5CiiEiZE4ICtV3H4AXu
0vemwJty+VCdM8vOLuYQxGreyC4+f8djTSYl93+p0jZmHLRL3aVCGF5tZ+x9W7ofwGYU5YrI+z0U
1ncxxw2I7hPs9mxLE1aQh7akFjA20QjhpXSCIWBuLPBTbk0K5fYLRIkm6SSwVtW2Z9dHJvv4n5uf
jTtncmV7cNMYOFzPkd1d/z+9FvriOa/qNHn6tOPyJyRy5973MCUFYMrPxSjdqh4WPw8C3eor8PMI
YsnBUiW4UTy+qdK+DC21AB6IKP6VWGscFP8nCFn5aP1bz9fFJH3RBmX3dPLWlR4IJKqOl9myh+dT
CPEvxuYywQ3sNgu4Eysmc2wwyUEQW5e8csii7s0ntcnMA/GG0vRO4jcn9fdlg7n0kjYfO72AVWWV
GEY92NjZn1A5wc7zTsfMBIGQqci2osnxNs4jycVxQ4VnZQm/Y+4roXl+hz9gkBCx+o5fqa+FZB0+
kyAezNaqXfeuZ2N+97X+1WNeELVA0Npfxd4EufNgE6gciTnj3wpxaDlJvgpjf8FmqPuZZPJG9xO4
/UC5P8yHxfwEamOGVgqI4GRyuU/q7JzOV0uEjz8wW1nBeIC08JLmLCm1zW5IngmpNRGZUDRCPe3G
0nCALJnh0fx52fBZAOOKtbXxU/sK8NUrnB5Ooc+xiNVkkeqrmobfEtzF2nS0rZV5CBtfPDmzCH2a
YmQJmp4wK09N0xM4upR2c2OOe0VY/cEAPdlUhUcjAEWn0WNa0aE3crxl/BGgkQonZ1FtZDGVe46L
qISBfohDF2vPNO1QHMdil28jbI1l2chCl1QdTz4xgVLTSnvKChZoFICK2bk/njA/WIX/3PzX7nUe
XHzWQtUD8GBhiXHp19duEz6akXhCrxbjsuEdGj6eVoHnRW7ccOTTToVESo1zX6Qj/eTeovvJwQbw
ZqWAgMIru+Ab3TKxuPMKmY/hFAqeo2ZqSHu/ewByfzwtyUm32eJwW5TUFRJt20vroByb8ItL6ze+
BToVSgH67TgY9Cun9gAHal+qAKV5Cq/oDDbnEh1Pyjpxhk9xsUzwR1S2LVSlfJVK8Xxh1IiKmqKR
32uCrg1I/uEwRM1ovBYFE56o0G36rlsSebFn/yCi+H9JI2Ifs/4NXMtJtihn03UWylsPfuqX4DxC
WJzEaUaWxkEuKYureHQl9Q5v8v9neT81lJnUN164UqjnU67yz3aByyBiUTgWooFaoxjWkWI/n6D3
zfTf5gZnLLTtFJ7mlpkma2w0rRbqyITZRGHF/1f15BE1FiIvin1XWZaCT+4EN+Nwf1+PKtPlM/tt
wDTE8DkQYxH77DgzG2XATGR34/ior2im6UfSMO/o/rZDnX2mJ2sCeaOmBFIcmPXcU8H92mbjN8ym
dW61fWpnTrCN3piu633QQ6pHkfJqplor27G/wGfArcFVkM4TE+WgrZD5EIIBkq5PJG77iEokAFQf
JOxaHMu/mnGFSOzM12W2HkZI8KPivE49CkiwlnJTh0/yjO6m/jvLdGT2xaAYBNoTQxxWBdKvVVci
WTptLffkCniA0EMxOgniwcxJfUb7mRhvLPalfsBVhV027KuqBKbtatozfvahdeKFdtDfGgiX9O2+
GceS4Mo84zVPIZnm/g0WRnA6/px352mJuIUP+6Cucd5wCSeqXd+gR8llMkFaHs436G7LZANuutdt
D0NHc/erz7Vwdvumk7Kb7WndcxDbsNf69fTuvWTrrtGGAZT04yMYJpAt4bONuS3bPjZlw2EidW1O
rJGwXU2CU7h3vkU9OybZhBUx8BswrFqUrspdXEjGVfiZxMSI8ipJzDpxAER2NWBNkme3eYxS/y6o
OEoYp3qQb56Wak1ME9zKTSAL+GZMPVijAYj5G0lPZMvZt1n7Y5MVmejIzf8Cjw/h9AMdoPFD307z
+9hdBK63DRkzGRCak4CcGSqMvj66s2sdosnqYDUAjU+kRbcSTtkTD7V0pUbJskahLhEMou076VQQ
4ulDQ5UyuIsF61ltZj9WU7D6FszEvhCFrScp3Wo557n0S+fOcVQtSUXjlu/WGgwdQLDgsdmGW0HS
JN9MRsUBN0uZevhv78Rij9GrtpoZ8nEUyFhXftbOtg4q5dOjHHb9iKcW8GskCgkL7JIziYxtdnif
3W19o3uSbSQ9dze8E1PwZD545Gu137GwJwTR5OAmbOfw8j41gOSaAoa28m0Qe4WX2TNe3waxP0HX
aCy2jRhCpyf88osOwrHdMdusG86URXvTI5IGLERTfyuas278n52N2IO+IxCbS7drwk7h98n05LGx
qTxRP+8Ymk4ZCB/60zKpI7iE3/5P/n96B09kM/tD0ULYY/qbYLhNdBfyjvcsRXYN/gqmLVdRhbrZ
0HiHuuJLAZ1wAFCTAuKHa9j2Zn1ZykGYU7eCACHzorhrTSjO0hWhImrvUo8Q445mvpD+ixprcuvy
4Q2fxKZH6YCG/LenKQO16AhIt+1Fmgs6pSxcxmCWsaXaE+V2m3YZXN2A+RjegEKC+TDDaSnfb6sx
llINwk2Nxr/7MsW/tG3t8BBC9urtzzlJHczAe+JgE23eh4GLCQ26YbiZ/AFxOBJN1zXmlTr70Yhd
f10ZBTBIpN6T5m1BFI44D8tIbLHOqhdp6FebMzE5jJOqk0/0SWz0ugxveNknozglk0z2RJVp2tws
PSoacYcLZN3b2ptU9BE7WWV38LmpqtuIn82gdAlXIul1w3EUj3QbuZ3SfOFcKFjv6rjdzWbVxZyJ
sdIT9jhdpIgYRoQQOBrSUWubAeul7lzgdDzeYPeEp07+ZrQ1EMydInio5jRPF1uP2uIDJbaXy8DK
h6QRJrkyzA+KQZT17RrN8hhhOKNeuu/AnhLxTKLXcn15aUnsIYh7hd3sfU1rGqU+BFmF/cK9RyqU
Slzn+B9dj6qwEKTVGP10Q/rqrR2nydvbKYpv2UoW7MKrdYOhOfN3vJDvI2ifmatkTt3bIRCSX6Ga
EKeWqwK6tEKBmSVeoDhxSM8hnAmjSoTYAYGpcvV9pxnahl0OpLOjMaj0Pef7AxLzAk7ZVHJBnwvh
zKHiRLgZzxjtetb3Rk1aR5f8zh8pJgdxXFE53tTFAadB8bQ0yIiMilxNho71MZJdwfvDRTSKQB+H
PcjywfOZfs8BWnoqnwV/yhiRQXw1a7Ggg+e4Cukb47+nyjv6mRpz5KStQRQA7YtCR5BuWVuO0p2d
cH8JymJT/IybS38tS6sP0mKXRh201KxiLYsFVR8BpJ/KDL+nnORrO2HZoGL94fm/6c3O9MalNoVN
cGVoDX/Ggy74PkmAOV7evoJq4Z87x2J+93sLvPdPmzrqYnmWc5WvM8i//0tJ0EvYwVNHx4D4X9Qr
D8ByWnGca/T5UE9SX2SZVbxos9gZFRmM+gvQxZVhIZLG6E79hp3fgrQM2TkwcaT4JB2qu4H5RNUn
6o1PEw47wR4zDXAHhPKcEnY8+HPh8HDdQRnUQID0ayz8spaAMxXK/uNKNZUFNtqgvUjQi8+tetuh
Zw25/yCGuoPmdHmU5GQjEXTT9AlezVq+6/TG70NACV5riQMTaHDJubW2SAY54GQPN0FEV0nI2K9m
dG2UWlaz2ZHc5ajaKPyRpieQfVWqRnzFoHjLuk7a1ze9M344S7cJ4I4JiNPY50tFAT8dctKB0/zs
ttV/WlYhk7UNKE+ccSl/WxOhJCWmVGf+zLnApoIHsTVGjCZlPpZinoAdhmia1qkl97AYVcLFiZfF
tA1XQ7b40z4ZSYjkN0nrBKdtCR7OShhQmrYtzTRniBu4aKoVRaAyJUrOWAgk6t1OzM+BgLwTXkQI
G++x/Zo4Vn4IEQ8zBft4QyofO/xHOgU1B0i21g0SWn0kLkIMC9J/+ra5xwvdVWt3gnFhGNdK1sER
O+ujzdwo3OnXCHi+HNn20w3FGsYrC0zqVLHzC/0IRNsZnXSeRsMFzkQquYij8b8F18Wk6hVYQ7Ee
C3sYFjWXllZbiYAQyQn+u/Ms5OPT6FGurF2CVUFu7ChBEClZyEYxAZMkVn+mO8dDuwfRFdJ+fvlB
wx3nc/8aZgVoUwkWOJCx/QL7HyqjpaiXO8pB0O4WzJcAAIvlTocq/wiBategfxIdtoEd1i/4Wozc
lwmYujOZHIi++8qO7E0nlpFghJimhP02NOJYTRabDuFqb1AEojUWeZeTXFujvwBVYWCplIclPFhC
sUjFa4H6Y6pqOT714ASxu6YXCIkgohEPCgTCWVDrcQcDvLZ3j9NM9uh4FAfYNwNqH5s8Dq1KTTtn
BaUnoAyIL/QQlmqKJO/9hyKZ23+qZ5H9G5831ENelG9GMAkTtLK6ImjzSwZBV8+L80dK/2bQY/+g
bw1yc87FUO9da0YRy83D8ljAWzyN+dYnJtYiYTFwEqlyLWBikNTB5HoX3N/D8eEX++Gcatj//FEt
Gdb13/eBcVxCuMggzLU58nfpZxVWi4ZIYl75X37N4yXsC1gnAs5bNRtckOvgSOpczFWMsYaHc+eU
58qTDwHNZrkx4lNBYpDmc/fZ/eqr4J4SQr/c/8pvJv/k/2IWheE9Cg9XLZN2uPiwUG1MpZxCh/gp
9Ju7dr3grn0dDx9d/+0j7g5Gn6getjOcjkX4+CCNvdci3e/VjB26PG9V07kzdGIwWH8Cd+yUl5LZ
kFHKz1twFfVjPWncCosCYbMGTQO/ZGxfWDGDssErKY/uSepryJxOdA/Dz/VmfpuAR20GXDIGuhku
/1FPbMUvzwFXm77dMajb6TCUOGyANa+i0efZZ7ErZDPIC5WVxoOfntdXrFOh8h5z6d1KvMsBQR/o
g5kDA/c4zZKLpyN0MFmuBFDQEn78TnnwwH3y5NkMMuFQ1PUMxhvUJ73nLT0zJWpykeI1EDwA0oFB
7CDysBUjoeG79ue72SWFgptG4wh4lP4Sxg1GrmsRIWvM2Va0YsdkYQlwC2APcn1Y9+NIZMWcXU/B
5Ygwduudjz6neUiuKL7RciR5jlrWuCAkNVHlK7uDC5IbRh1dAbx7Cb57M13KLgaFVEuCmSBcqART
JofFRXpMCx0Y/CCZUYoxLW7fc97m6dfhs2PVKx6Qc+WJwNi0QyC7Z+0h/qXVwtEzSYqvaXK3ptXJ
onHeG6OTEo16MEe/WuE0P/EHsGj5vMCufuDNR9/h6t0+qjuNqMzuz78t5uaGuhD6j8ZN7IhxzZRW
8pgqEI7ljJTDbjQOYnKZAbysRZy4+clAeVH15QmwTOi4iWP61/NtIOK5n1zudXNYDPkPkECLL6vl
iuQMa8j66JPdrAdHvtn945G++QqwuMZOCcnzzBh8cvU7OyQ212SYE9fwIF3/RbQMvc1uvJDkT55A
ruJ4yNkux/DjsdkrAiWWwOcY7VclC4Yb+YNEXxCJzhP+EDQvIU8hT1CL2G3ydxOO2IEcvWR53bU8
Z8ro08/Qq7nXjR2nsrzX7DBaq2m6hf9VpW+M+LRAknWuMGH8AVxT339MHnwbDa+W/JOyLIG8+6uD
JB23kPzrj0fgQBilpXsenJIAmFcHwlToaqntCYKSsgFRxIFOJ47ZnLzhmWu+Gr3nB2LBF546TW21
BuZeAYa2EB45E01IenexYR4d6j0VO6L31/yTTz9mEZgjAEEAcl/lBbCldHThYp4w6p1eWqhaXl+G
PksayFNeCUKysz6QpRRfOCZCOhNdUt1gjscoLHsCTx5oEgzskyg4HiUELmhoEXJcYFLobBRAt1cQ
Gfg+LlDpFKtL5BedF+gAyDUOExHrl59CogRg3bvD0LmOL+HulAeN0tYaQOSaWY7vGpNuVOA7+SMA
SE3W5mXZm7+22PDcXXFtJ9JXJs9JqmhwfeM3wawUHVGooRTGSLGv+GClSTVYw0bJwdKyBA2l0Et7
H8n0IvFa4AUm5c+C4Q8n4vfUnxCLTF4m8Gas9zGUVYWzuiNFhoAuknxFrPXQxOq1b8u08VYJFRso
5slSa6jTnS/bNg9VvSBtU/d7ISFDs47VWpLYD+4lBCf8ypb3fGO2jdSI/YJyaUYnUFZ+afrgO3Ox
E5Gt15ob+pOoJu1wXDCVToWem3/lYxt7Gg/z5KsYAPl8O/o7poMZLOSjeA3I7Bj1FP817AeFrM1c
pPIt6OVE36LqSI1nN6a0yFVSq1DFkDs23HcxayvPHGlXlHMS+PKCDDiplCfHeHDJjexUE4hXKUna
Fag8TIpd+GB+gfR/iwo212+DtTiTIyQA6doBYDco73NfchbnlfgBmBzG+LHfTxpn+gVsMIrT/RCS
Mt1TivMVRKSIBYkD2LYy6tgDxE7ktM2IZFLw3VG3HLT3Q8kCYXRDOpB5mx86J2745TZER9YYxcrx
jNYcLc/oUMFOWvaK0zscoNrVV9xwSBksfIdmq3woEllNxEsmA7sdizQEOYSSjOZvq2yHLts/RMui
84aJSMn2QI4YwqWZ+oglB7HXcmxYbbRffHKkSD1I0YkvLoED4J36FOq4DeQGy65Ff3I0gJ1vzngx
kNsKvElNldkiMuBUFWdH9Wt7VtXSgohaF/hO7CKtDNdVW+fitCCegfeyX350AWMd2cL/zl/+7G4Z
4vtQ/iG56vTJIyLw/EgYsMgdi4HcvUL2GbW0b1eHFyYaJESmw58KYJz3MDH+m9UMG47R/A//bQnR
FEnL1IcHwdyQAAez6k8iZGYkTAN3xkzx6Nj3PCRd6hpW6mLQc4KnFMWdXvsg4AhZDJSAmFkmPptQ
oahxwvKYNvORmt3zFp7SzerKfFtClwjPGS4HNzNGe69mTdcmEbcd22z8aKWLaHoMS11QkyAVbPX3
CmuKM5QrBF9ljruaUy/DfktTGPhikGFSQU5LPUhY7RNBaENXuozib7v6CP2HE/Gl7b14SZrO6jc6
Nu0eTt4FA0PorwrMsZL0oQ/QC3Fx2w6sorf2OZ3rGkyObJTQsXrjxv2/vi0QF1HVMbjwaMHLNQDT
agP3bJRo/2F0jh+szKf8ZhYJ2WJIHKC7ftwfD73NjjRQX28T1nnmE9RA1qp1fxG2zfSne46Yca4W
9v0Ju9CQhEeg3DCxZj9GULOsafUd5cdK7cnzytRZKbCWCLbo1ygZRENiBdZ24VhGU+br1yLWzp13
GF2WPgPYarCgJh6wFOqlrlaghB8UyzD59R32IW+M2iRPk03j0XGlLIB7BiM84MDzpOopLrH8TeEP
ZKyeNsl6GdFYkbUsH5HN4E5dJquNG1MJg/XjKAAtMBcunQiBx8/uDF4gT1SLAKhtB2bzjqhdps7O
vIDL1DWA2qosxg19opatlOMNHVIxvBlou9WdZnpw8j9GzXgkKEWPE/9vwBbWmbIMBLTZGk1Hnk5I
mA39xPoFQpLXhwCci962kRwl2r6axO23UyvOeMpttXdNCBjnQrjC9l/Ea6ptXGMERPIVbHZxnpul
sw5gpupj/fnyaDGAU8tKqORF0Zw9na52Lwe3FwY9p9/IMv2VYbL/r+bwtDxYLgDDw5TLHI83Wjsj
GPqi4BaDl5C3GhA7uHuBnogBiWaXHZcQvJ8ch1r0Y7Uk4SkG5Q+N2/hydt2CTS7y4UNt6OTt+ALH
0BzGMOjrhfHLxQkcw35OlL7B1JEuq6FF7HHCb9qciAG2eM1GggIGgbn8aiRAz40rz9dWOIn5YG9t
f1GnzAt/2LWJdsMlZtnwNZCnxkOToGnp8kgKCyES72adVHpauQ7xx8VOKcbcPRyBAdI3d45rrsrN
swNdE6uTca3d87TE0wyUpuNq0xzPDrIemrqgxR3lzsAWzvJyrtKUbpp6+SbteZBVv5Z6ttIKePNo
lOBJ7JjrTX/6lAQY+A+k+yxu75ZMGnFZ+rNlNGGPkRFfm7aEWrOhuZmMCXvSRVXs+8N+GEggaH4A
5dyjJJ57udZ+cyjNA3dmkZcajo3XiBKBnFrUEKmliGSWGEK294WPiHFd37gZL7VHccIFsx5WY3oR
s/HlzBIUAHju28PRhzHSLa8tVpHcCSc5SDXETl6a0uja0PKLU5UrP9Dal7XpTWJRI1wWY5AIUDXv
C2GD1KsyB+DX/GtXOv/GGYS4oyjCnZI5KDHihyV2eTM537UymCOARK3s1fGnscYrN9JNiWFt3GH9
Qw3eihpe+JYVW/qz6e1J4zlnDYDAQIl7l20KOR9c0okHkyY8DjEniHVlj0SxvBGPnNwX/Nt6ob1v
H9/3dX04v6PUwVzOu+Hva9E6rDK0si95qNRzssWTrLM8t90GRETLofv1/99FXb54++VnTQt+ErZe
SfWI8N1EZhyWt68qfZS9+v65yIQLHUTsfk8MLbxDkDGk2YlbpvHTKl1/WoQJ6hhUnmJ3azQOshr4
vEI0bmPvTOLgnA2RT8auj2/KbnJUNmsMARMw7HwkLM3vmzxc0zmXQtm1AQ/PkdFeo0hymrMLLun7
x3+SCMlP0LguueypAwCfOuPLzbe4I+SN4Ge/yNXVlxifoEzcRlI30bdkzuLuGDeAuNe1rTye9OQP
5Vo/GnMO3znIdiAs9IwyB3YqNtff8ysyTpqFy2WgZw2prQdDd0TK7yFAKwruzKvjuRsgi9jlEtLQ
X2YUDoccUg28Tca9m7NVe2BkJ+07rbd+yz/eNFsVwVUktadyVWItOucL/SXkAEoOdZeLzijpWS0n
95v3xzIw0BKsSBwiKYP1/PRlne9wx8VMUkcLqpMHeyyH9sBMXLUMYStemzTbwl54sjIM0mtrJXrp
IQUogBht1ViEiFatZX0TTvpVM7f1eT0kSEjO3+mF5VARC2VQnNOffzotdRVP5gTX484RoN27Te/y
I7COjWBWWAUYGwyyynUcwJWh1BH1/272dMJWjRM3ZTzS7Z4Gol4awqhe2A3U14+3ZYrfiES+N7rH
ivJWrF2vMljSybkTYIzMPh30MFk5f6iZsN8ydmA1JBTDPepa0luU0eFyREiGH4vO58U9vqc0VPpC
W/8IyNlSux6Wx79MN9K7TVkyElFKfQKrAEibNp0yEO2gIC1L+slEqRWFCMm4uyCcJvsnNxXfnOj3
PmN2Hw/7fwrNhRuyKNcNTHLtCDfo8c4aX0RvasH01Gjv3KB+Pr8v7zXflDHm4gpBye1a63ZidXOK
cTc4mq0bFFFo7pMjio3CQZ/nNDjotR7t2qTaoX1z4/02MDm/R4yH7EuUejRX6xbnIGgL//5tCfwe
FelRYqL+vOwvuTOtxRTAltwB7xrfud/iXtJH/uqikGcVK7wWrFoVIK04juPGvJc4V6wwmUjtBklm
b4lfAbxILL+FL3C80S+O3XJR5J78mFzpkUt2t9ByZ/V9WCxZfI4u18aHJXqmZjV+C1BCh8be9dOZ
DcJ9Hk3tu17UfvxOSa+ga6l90eWoHSMLiuFQC/8A6Z5y1DYyh6SayuA8Qq59HwuCuO9pB5fexkFA
E6B3SHhTa7DYsffq/JeAFxplQXgZpcWBk8dOWS69B5Mgj705aAHFibVra5t9mrnMuTiFghQv7cdc
6NXM4OCwdjqB4vZR06QLj9FCp4eVgX9/24vTnrz38BAypqdgxVHYa7JDeG28BvkomVhlnrlMr/ta
kDg8IZE3mE5sW3P3h8pUf64PZTfNBhMfb/5NEDFHsMY3VzplA9sB+h6t2bChl+FazvjNq0dAP7JX
n+6Sa6dAYECvi6NeOhhlGFMeK1Degpx5gCMVOW4VNy/A6VgkcGxe4Sjo/92E1rXlRBwTeIQ3nudO
ylMatdQD5vG6tF9jduB3JxM7shWhFiiPSR+DVmn5MKwRX4pKLPmWd+C9nP9rh0MpSUzYcOGFIyxk
Dg8hJlkR7xET9dKBtY0Nc4HXE7ZxJI/espEhmdMZYJnURT2EhDYfeIf4y9OSgQXGePtKsJew0QTG
5u3RdwrMTUpY6WlDEnrO/kn6ntF06kD85lCQ2+A5z/KaLsP6v3W+0rayc0SA9pOaRx9/hbibnFht
Ef+RGGdXJ1hhu67q9S0XEpguuknTqEBoRuvG/w0uGdPsBViy6kQDzsO76d3y4VtRErS5d8iwlyHg
8n7D7ZqcSYvmG6K7PvI5fNUcPbnej/HiUY7pb6okOM//VXvPe7Ux8jOgHoNc1MQecKTk33HjIpQ3
lF0j73uCySHBYaoELTBCsl0JePbDRa9y1tJiHP1Wvp20cNc2IYAsdQIkzwWSXgEvF83x4YZbGDIO
6nzfkKH9KZctWIM2Vht/rAB0i0uvZK8pxOzrMqE3PxtREaD86AX9KZpYjrKV8Pt3LYrSYPq0td+q
lp+fobtOlbpj5sgbDUrWM0t4DiXonxFX1TcQ7QTzlWPgKteTGVL8rmZFlpVhY+faGNzOMGzbNC9t
sGRakm/m2olHBsPrZ6oJ/+ipo/7F3oSNgpshTv7oTbvIvVpI+hqinGimUzEne+EXmh8J5a5KkJxF
UFNfAg10R4BGKdZ3JtbPuHBN7T3ZVUlre47L0ugmMaf8MHczjRld87UniTjoKNWV2KKMx27LR5kC
pKelGk/OBwTFAGno8QbWqqVmWVEHEcxC4z7/hJapleGOKt+DySTvDpjDXTrQFDSPyAobsCYf6uOf
MvMssh2v0Ac4cZT+WzqHEz6ie2puEINogEXMUoSRT9jyQy+qMU9ii37+c1f17TjdpPDEfRspvv2i
4TJw/8vIJ4Sp8D6Mi7fhvXpegBLD/qI426kadR7eI4r3ExPs/G5ClDcXdYV4Mghjf5gCvVgFHo9o
MlO2lafTH7Xe6iJWgr09EfE+TzanHW5vNklG4jV6o9NlPwfrDluZ/V4kVk1icIbep/9Ve7CP9JsR
kSlLdd+eTKlBvfeI+y0uiajy9rySgdG9/g+vvWPCIQKf4ZaLX03u5se3U5dF0MT0bUTbUPMc90fW
48EKdz3AVzcr5XtHx/kZS7d5/Cwa0hZyhw/zaazyCpo1f86e8kdB76PjqtHnuHGaIUutLRl5TRe+
rhHoT1uaNgeAmz3ftuZGj5K5JEVXefMjYxcOArSQZHawnVHKJCdt2QwUCj2M1ZpZIoXmxSFgtSdf
UZNaMPuDoV4k/PXKDwNBIj6dCqaa4k2agXgPg58mSlJnVicPnfTjbZWOGK4lCX1E8atEv2iYOizz
Vf2+trFmGKPrHfOaKvciOBsYgHF4znlbdrkZmjg7BlBQiXbM+0yUCBVdE8OJEaZdDMXM3NtHMCQq
ClXYdjAfug39KyMcMCNt/ZzEqb/tly3lqbbmi8kh9f91gYJ5OALnKDMPt9AV7UxVcgriqCv8KUhO
ECbCvILxbEk7IlRhd22e4i4/5Sk5dmEb9ysAf6VSOmofzePafNxtTwORe5vAzmJblQVLqr0spiqH
QLoqQ/wzG1Dr4XsEK2pKtcjdAjaZtCF9V2MHFlxiBdH1FLWDwg9iiWOPh0+hBLghbQLdAIv3Hojw
dvFjKDMhCB5quQ4pIreC66tMsiJh1ESSiNBh+8ohzaUvCQTdXBjOLulD9OhoCC9njcEL6xvLjiWA
1+x8EITmIusK+kCMaRw3VyQc1nQuC+2XvTutJarXUsElipwLQa6hzIB48DWVBCg7YMR0JbcTy7la
MtuKrlgKXdDL2emgZMZob9c31ssJUBRH+UIDfRbGOlcVglLKxG5WDzTTntosAIKz5RKwceWJNTAY
6YtPDpFq49miThicCl3I8jevYT3X6rR0xGS2D/MS1uhb5zo7W1LyNmpG00DvrAAEsSrQalTpxSDp
OkgMR2ZVd4CNPXnHZdpftWLSJ3NtSxoWK+XVcPe5wzzu6TTjUGdI0GKwzRk5SrednxZWiSrE49zw
yXbtDkcSY1RyaAbee06CIvH3ySdtGRpI+Uj7OkBn6Z0R4dobyTBcYKbR9C0/WF9mXZ7LvEOsaOhk
U0gJb2eEFAo/fhTa3MK0XSQrBrFA3FyWyDTy1eQ28UJwFGStpEOq7IJCudgvSWEGXfZu118uR2dB
6aaldFTqb09OUmN2J+jl8/eAWIZoaI49wHEHX2EsZJ2Q2Mn1qCEM8onAdTUeNFPGJ+uUWZsuP6T/
l4c7Tp284mjcxL2QKkHZaiQ7wmKahs2ejKyYncag4YxfZBO9m8Vem1BYnbKduuxFOXCNRXJWzUE9
5Z9CnuEZTg4lcyT2TbSpOv9bwjrv0JMcs3hdYu8fnbeDeMsgLxjMqxtC/7W+x//WXnilPg8SntkS
vbSiJT7Mpii+q+HoQe3403S7NLIcJXq1x3dtqZQb8RWqvL3jF6cl4894MH4huIGPbKcndsxD4Xg8
ZPal6xTVnKhIPqQWfbPPJlHOi1mnik9OXIoDaZSlCe1rNs/qxgrwQjTWp4pzs9OVw7lNTnO9Ul2t
a8MM9EWs+Z/mwOGJSmcs2oJhxDc2YoTHXHSviqzaX0esfAc1wXPkT/bA+tUdUAHYpXPljPYmZK7m
6I3wK6bxW3lr2EGoMM75clCl8vh6a4IjpEvglB2HCko4wDp/M/S6GZNYtsNv8ABC23LaVdKi5WtC
6WySP5R29go9gOQRNZr2VDRfxLd3IMrPzNnDi2tOTxKmKDUeT6A839e+Za0VMnB9V5X2s3rAdbI4
T7YOTOW1+iB/exGphRiwHC3vKU7+yn7oUPHZIuvkZAxeVAb1eMLzgxfJ84JO+EMXN2jzkZAieVyF
qJgLmyZL78griZGk66i7Frbn9Vlgcz7ZgPHOLWvAuYR/d4TBXWGb3WpSo8aAR4Mm2jx/bgASUQz3
rRBGrdcAvow/zzxfvUw4mdo/fJ6afqrCsuyGco7vfNWQ48WZVyRwt6VaqvaM08Yjvnh9TSNmmSuc
B77wlouJRahwveMVA9L76x6mqLHY2beqhM3KJW51GIK8/PMCbG5qvc7KhaZh9M41yoMA4XG/nuBe
qgGnPZqP+WaLNRdwoeeqf2XGtA1eilSoGntEcK7xunK7BlEpD5tljkRbf/2u+1yIUx6hVelXm32d
p8COgy+Vpwikl2IDR8/HX41w19PPmMPJdKga7yGnyRM4X9J5SGwX6WaeggXD+sw6RsHT90v7TVzs
bmj/m9ItOpjKdrcekl+/+QwSkdHpVqkxWNnRlUYgVQMkwNiWUnFi9OoLU4YrViDpuH/7sB3fCArU
aKoeXIzcX+LhfI1u8yqjPn451OUmLwF+fd3NXK5/9VjfvxrJRnuUiUAFzV97U8pmnuQC21WAZU+C
VEMtccf5tfzuKB5DtuK6OTK6LDZGlPKPhKnQGVXfF1Bw0ZKtpjVQE+3OtQeK/iUYEcu4BeuZK2N+
uCTowjx+MvcINjuM386dZjzxXqjMaH9rFDrH2HT1QNu8O0Rgt8OIl7gu+DaUbLe1GBkpiATU2RyV
ZlS6Fi0BbjI2Vj3oiaOIQO0ujtZ9zmuJOrg5Fzw6/kZRVu5Dsk/NdqiPyalfzQQXjIXGP1BzSiUB
4c1z1F+6ZaZB2nTv5ocTVmITUUIii6ynN50bv+YqIqXH+OL7lws5nrpsts59Zq+TdBMyhKuoga9r
YXOYgYol4zQJJqGC24dqINLPknW7STsa8chUy6VF/DWDgV9U7oL7pfcrSsXcWon4bn/dDesgM6A2
p9kxeKOZVOrP6YOmkO58ijBFUWW46L6DRmcrIWoFWYQOa/YLxIq2Xz/rwegVxjie8BniuFX36A4K
hPMlZ8FkVhDo+nIL06f0tFJB2gHmJ590RWl/p8XMue3hMqQniRylVkZxZ72d/gADMW6TDzPU9ZnE
TFtOnRkQLsBSFMZLlJhmc+rQO+A6xMe0vcIMAktIWijRtV+UtSq+Hc7xr9GTi/ZammB4ut267h08
3Ofy+M5XPa2+ub7cPcEwqEYkHBjQs8Z4KEPmeKKfE21STTfOImjlqSaGOOniB0D+BP35/GZPs7N3
Io37u1kQBfAXDay9T+I6eMFvq2Qr+VG4/zHRKpQpZszQHdb3lLkGtNz4fuDLIwz/TIqZYTGlZe4w
Bxf2izpCbNvfq7RblW78smyyDHkzD0thcSIMoEoFEQgm8v6OpJRWCtzm7UWw9aGOgmDicgPgt84J
2HguaPzDwTRqDsI6RsnUvgdjvcntbZDY3TLnp27hfEDfHi9mcstArKDc5yvHRHO0ekMcZfvUNEZG
EquepcyFrcy9DSgU+cSeMYyZTBbRClxc2Z73ULFNBAW8sarTtVXWqZJhib62qd3rCkxAGYikatYM
yLOINDIAIXsIwxC2WoLiUeaITycJgp3cthZvFPoOYXxHHTeRp/wsWthPR4xNiZp0IypgOGevlOsJ
UljRiDQ4XdIXu0LOwAs1qIgrrmWkL8hMH3liZvCDSydKYP/BUHAA6Fg4WGU7ZeqMM1RxDR4iQbrN
pXRNuz6xGrEX+PnqE4avHbLy2HF6ds++IcsmoQUmTBHCK6ZO5bNRQg680+ZLmyph/S3VZOKr3625
qGjmCc36khVsiZUH1bu5RTWHI66R/kcFpoEJRTjRg2Sk+woaq+XLgEoqltbReBd1jrupsPAO/cTg
yg4bFb+2qFbC6iLGsWmwxxE+wKLeV2pFQb9ZmoZJNcNHxiAjv8gqp7qga+amylkN+Qnqsqfg1pOv
ytIcWP9sQZHFbZGcFFp3boqKLvxGYH2+Siax0QUTBz8ElHufnM8Bduq5MVQEWMDGMroDyeK8Q661
S3qqRO+m/QQjnllvMqT6nS3Yc0nTvP0S8hAsEXpSpi+D6ypaatLd4URkdnmj+SNgRAxuB1B71UWx
gADvNnD4ZHW0+Q/z2LsCS5byxWn/HaAl27Jp0J/i33XPdSqAKQFXTcUwIYFRmfXmOktuZbV4jzuE
adB8ga7XqVyanhRPymyHFKNkgoKgGqV72Dfk4MEyKtojkDOhaPEo4Fkjoe5GbP/dUHphulZitYth
UewP/o0xcObo24KPEIzBZZy9lMdx4nfaNzWYbBDLsXLqg3zCfmsr9F2Ajv0CiXI81BV2qATI4NwZ
gfUutRmC00Cg2mVCnc4mMsgK6P1cTqv8OMK6wSERr/vFdS23KYmb5JWKCnpVAhoETLX8j9TmXK84
3cBfZ0sANgA7JZEBfG9gen3PsKbbv3+q9FaQfLjgucs8Im+PMhAmLetzUHV4ypcHTeOHzVFyunMm
PwsQmfU+LX3R/34y9s+sHCVsuOJR2DcmHidsx7GylLXEv0RejJqsbzKLHOVPD4E3i4DzmrVi1Phz
EKu2Bi7Bb3U4+risybXkvHdaIP/leJm/a+Diea4At61oJ5JTtLcRtoxBBzetpg1jxrGoKAHr6SAq
QLL/AzMFlDR/QWf4FsckVr2qVHWwZOdIkPg85tzCryspLGsp+Av1JzI/i9QyggFVvZaaqRUZI3Jh
9AR1OgIiyALDZZ66PAySYjBABs8NH7h3yI7ypM0TBaU1neJjHcfXKq5X6EnS44bI9f9DXc7h7khl
pxnNX2Qt/dO/JG0hhslUwenm1ib3jGAdMxJmChqTXB4kFpQ7raVq6liT/q6/txDn/hSHf8JrqxkG
S1Tz86ABVGgKPRdx69ETvjpLzEuSnBBXnTFQOYlLVMyARLJCqHBNhjX6VHqJ6G0Mu0PEplON93D9
HhOnxCB2LAZ09RIivwvcpw8icn74nPu5ZbFUJZdMgdNrIxSJx3D795YEWh5un+8BS1QmP0iIRbBx
E6u1Czme4g6ouqJdJssixuxDsUjUcdLqb6SmKMOcRTFMb8YgqfHt5/Ihxqg2I4BFTBh9B/b7xWpQ
nnhlXH9HikoJ2hC0VQ6b5On8Zs9+r8CXeAQrqlf2spFhJKqrOKthWeHJkyqmDPNq/tL7xPc6pIW4
BhXvvLojBz8sd+bB7SU5zUFhdT4KCg1pKWdZ2VnWzgnw1C3byvbe3iG0SAB6C7n9jwlAxz26C+UZ
bPspQV2E+tv/t1lTx1z3TBw8a458pS9ee8/SauO/lgFA5MUA0TVopye2hnVwQbrxRPHPmklYiXzR
V0b+X/TdwHAntHR685QxylBBy1cdNyd/1ef8J5olqFo3EVz+lnKkzW8kredTrD9gzVEqhExaXjPJ
vrZFHYLbYpflK4FcihzySVe7XNm3VweroqqObMnAc8I/X6+Z3Th7H4GALKQHKANvmcbemn39FU4H
zQFabeU5ANdmBQjPxP+/cQy00ocma/xs2NnVz5fam7D1yiOyu++ZTw1f2qVwlxusVGpj1TdINUTd
s+wK2v9POk13YR8hXZ4I1eLWaHi/EKC3ZRP/NBcw52z3Nhn/upQC6U3NfhPfHAWLUjIwGMwsrUAZ
poM2c7K4gmbmENZuqfK4Wx/9leF4IRiOPMV5+3DFjEOAY4ezPkCaPHcbBKpEPgqK9rvuNRFuSsVH
J+/Wt3dcsBwk3RBzuqvk9/ozGUZUrcLc7c4C2ofH9ZMTmNRrqYfPc4ELPoztgvlUJT9STVF1esYP
PHcMf1hY75QaQyNJp6naGiS6C4um5ijIXv3xSTDyMIVhFTDTH8nCVTsTAF8MMmvO54Th1oE1aM2G
bvHY7O7FkqrrPPImuj4pjwAfOtiftBk3tQfbWACaR5PZF31xAzr0NrK/z+IjAAoKg0SSOD/bt+kT
amhDzUdYfcvIH7IFFHtoMXLLJt+f8Ty/rxne1B5dZ/m3J4js07duSKW1wTrqg5mayMmdnwoNC+YF
SkbBC/6DKVbZb+95P2z8uNIdl9iaZTNgsUdrrDjM8c6Rd8c8FCh5BbveXgsX94u+MrRu7sNqRXTu
dICtxeqTZlE1RsdlipOiO7CH38EqGGVRmhQ6plJ2uW1ZS419F64CKxXQ5F1xPftspH2o9Z8vSY5u
1alaMvGzszyrbJyccr3azDt6oHE70aNMxNuASHF1aiiqdeuOIOtdQOlykvnnVhJKy1R7RhWfOXbH
viE1OE1D5Kh99b0zKchdHDwA5Wuq6Vw+HtyQ47LC4sgc+6ObPPLOEEnPYTTBV5M93LHlMhllczzP
C+xvN1BKCaC/5gR7N1Qic4lraFSswETCFp2TicDe28/s+pqdxaN7N+0PxI9HTjl92Hkv7kTfB7rv
Zc90xF7ioiW0Om3C1E8TfC6KAl7sep/x01P1xipm0Z1URg6wDxPWMpdZ+DVocqA5OmlV+yPOUtZS
6hLtmgdxn11VGgTHf+YP80ZdYfPfvP9nlyqVdTIV9LH/DjxtpFxTl1Q6oGoJDrRye8Ov0zpl4vIe
nlv0BW5WEzYyd3ws+BwQ4v8ImAyrHj+X9B0mMx52RkXeqEJ/UE8kDd2K+PrLO2EqkYm5efhsc75H
HFGritp8TEKYBTW0+tZJAPhHlRTtDT+WUGvT5x24giIMQXXC4yN+NTz+1MNPcEYhKPZl0Vjak5T/
0caRk9E5tk4Nz3W09PBCQF/bNmE5OfL0HtNEWnpEIgRmOYGC0g5mvQH4Yei0wtPdYTVE2Hl8rl2l
2o18AvUb6+C+/tG8hdBhdtTDKQ/fZ/Km5elN1vg3eIsZ7qVxj1n/OdhIc8j7KeCraelMfsn0LIHJ
CbWjXvna3XwPjTh5YvZYs8oylRdyn6F4W/BTpJ3I2bqhAXmrh29xzRz4Y7jj0dDghX7DhV4ftfHA
p/kuAFZ0deUhYUWMDeExS0tHbOjtU/J++FUdXwwiDHkLp5gm17nIp87oEfG+x+ipC15ycE8L1EeF
8MDT9nSJttwy8sDwpn8TerSK2dwDXANVJe2ZOCukIUQOZMHfon9eEYuy/XYDPMzOAUNcVW///C0t
9b4nlfIOfwKgRiY4mwK64G4DxdKQX94buAzVpX8z8JOTsTPKoc1HRP8eD10FfVUrlNDwbjzsdMoE
HxgmuLpYdRuPp4YQLkJGXypMg6LvAbS0+rM+bo048bMCoxDImChCCFEsNO0M7DxduXPhLE3GpJX4
wADOf7fWqgnTcaE5LjeaDIPNjojkzms5SonDbkYrOeCaBmD3fZHvC5Pp7JvFUWuyfiBuNqNiWDGG
6mWCm4cqwRBybmAopq6I5Mt2UYHwOK/mEmf++ZAQ+N5gmOZ10xA7XQhbA1luCrZcdWnb7HbkXxOM
4sPfstGchG7W3aWELYzlUtrTT9u7krM8EQn/bPWmoWol9rg1f4XB04MlKNj6Uso4vcFw6umdqPG4
Mk7VOjdywpS80ifSoUYAIUTfsuBLH6686ShsRcHJBNTVCI9F5ctHcxQZIwda9w5JBES0OmaAnNMU
krBR1r0obToo770mVcVGTI29ooZ+mvzK31420i/O9GMA+93WIJrpvzLlI8gaRO0CTLP5ogzReAHV
lb1OxTUqqKfKjV3JoecQqzKl7NajRuxun5ylcbnksN/pIifkuK99sP8ngUBRyAmMWD3DSkdKNaKf
rGj9bA1bINaW3tCS1d6aRikWQR+9DBIReic5OUR6TBmHnn+q4ekTLPs7UQbUH2xHMFhaGR2JXuZ+
VeUh6h03nnyb9TyKm5c8Ij2oWPY8V9XiwhepUCMWNvnOJBvDqCPVSLwUni9cJJMWDZZ4EA/Hi8WR
JxAnO6CrJItm/eBHS4yfZm/J4Qa7tnyfkX3UxPQ5Dc+BWizEp/o/9Kn2sCnhsmuoECMQwC90XlDV
5YpcZRyOG8/HAHIlqMiDcuupUcCNMfMSnzNUr62hcT79QRwD8Hf7n9WghF8CfVwG+SaVDNI29Ior
lSutxt2v0nRjEU5xpOOnNvM0HtA1Nz60j0CuMe7BkNsOgBv5/5rAK2fvxw9jGOqPJ3eK7mH/Nbey
9g6fGZefuL5VUPylz2lJl4zOEXRNsS9hSSAhZJrI92nqKa2xFicnDLNJMLdKjdzbYk0uLAONNFQc
uc5U5NjKkifYQtUzW/SYC02GAhvi6Wx+qOuaP68El83AqTZgEuACm1QQWlYkQuPcxB3x02U4P89m
gRm7A3k5welxudBsSU4RGrpdcgVcswwdTauEOETydXnNU4rudPf5s+ocLpzKUrMrqCSsXoUgAD4d
A7tcEb7mWcRi9n7kbduNQilViXm94RNquVhrqF+SQEWnpiWnbQ6XAseoZrbQ/fq10XmzrqbmCPcK
LtV+GNzZSGhxrS5F/R71TmB/pPslWP6Hgyj/y82jP4aL4mCtuAYL1cTfin9AIzAkJkAK2HJ3tWne
FeB7daA70jGC456StPNbpwWkLAwtB95GKm2D2V/biBtUYgrMDE3xvwangeOhWjxdNt20RkYsmXp4
IJdROW2ui6axr4a29PmK28PU/JBUZQq1G8wTXG4xIrG9tkH5ECYrfDk7nabh+Z/bJe89RcL8RNAa
N1oWAniG50IcZW28q3KSGINxWSGWd7BtzQ0BGQ+RBtRW5RsOUJMm3e5RUpQuHFlZZ2awXF6fbp+L
eMzI+Dh856Rl+D61GjxLx0PECqyD08j/PYVKlMNa6DfggbpyZMhVNotDSbYSTfSiMcWBjiI60xCX
0YSm1vhnhm9ewqX1EYl6/IsTjOQDg1XHC8ookjhXvuLX/qb+zqlzOpY6oYmZp8Uy3lPxE+619PSW
Pgq8w+HY3YPECs5alAjEHx9q3ij7HenYgPa6pVEVlx48ouVQIsgyXD8WmLORI/wrz0izAfSz6eg0
ofe8AQk9qN0gBSLrgpDBRlbgreRZJmE26HtsD9EZ9M6WProA1egxJ6xZijXu/B3vJiUwkHm0VBkE
vzi7PwFr4tvfEl/diBngwS9jG+CyTlz6xozNEg/XEgW55f3ni8jQhMTa8qkBGTRVXmn+qWYrBkRF
5nAfN/tKHztM/7/m1I9H8oeh6+zmuAu7jTvvWCLD0RF1bV2JORRsLnmjQ0PFzM0JzT0qhOiGlnqG
8gQXMkckM7dHpcVZFRtGmAE6GJRPT6SpgWNjEhnVcZy4khQRkv5C0BEKDCXp4SV+BOfEYF5V8ziT
FJEuuZKIiprDwnsR5yxPSPnSCHFpd5sdzvorwNlHLAulDVxjI58wNWTjgZpnL2lLyKG3Sb9K/J92
B23HJYl1X4Zm0/6QAmOsGAS7wr8p38PgLXK509Zn/g12L36ahwb4NpChRHTYL0lQhkTUPFV9ZuqR
5ppBSjlI2flMT/dR6OCaOpW41QGwuvJ/NhEr1rDyb/qhLn38TXzK/uL6sUDc2rwQlLc/yQEH8t4H
eYqZR+wA+3M9kCVotuFlIlCBuIQyxERV0vPDZhiBVywr0eMpvkQDfDw0yIcqsA+rFQ7Y2THo9mMz
R2IqQ7IfOfkLx4dGSWLc3FrJ01kTnLIEexettnjq0LMLEz8/0G6lp8hr7PA+lF+jafhapJh/1+MJ
UmmThbc9TgWtT9m9U0ff3Ak91oJbwVcirx38w37SCD6HKXxmVpc5il4tbvwOOZplsCeplSPjeNg7
2LKiHpuhAA/T5EH3xuJFDoiT6LmtDTYdSOuHc4UM37MwL+aXN2YV5WyyDiXD0U2RchdP4E0vMcHb
8x9EkhbJT/8fdRL6Tv5yxdEUeXgiiBUfhreSm9u2T2WziuL7aNlx/I6ddCKiM7HEZmaVrAR4Ww5L
7cYoIFLAyXxrncGThZA6BvmI90lXxSRnpQvMOiDvfYCUHTTJvyZEjm9NnoN9ilzn9ks+Lx3JCUTn
1yjuZ8lRqGWZi8bjljS3zR+KAkC5Nit1GxdmJyu436XthrqNHWyAkMfLJAJ8edBxJSq91r1Bk1uP
23hcAvJ/2xvQB5DRmrEi88cN834rtVv1RVbqvpjB5P3Q1YV5MiKWFtFZh5xQRYqvbNT5xzZpT4Fg
zO3S7mfwMx4L8chJ8O45BYLeHPd8nLaQfuBcrrhKUKUiu/x9NIfGJsJ5nImSrWQgStd+gcBvnwM+
3prKJ+kXZMOPStsVaPu+J9ilx7DYGXCepHZSJnKOb1QUAgHMhvoG8Hz4W8pTrfErgzEVH1Yrg8tQ
OOGdNXgs0fWJJpGb6AA6hCkYIfcziIKno8L87VGRdHwmFTwcmq1fRcINB8QBKpY1+mybnqwFFnDQ
xitTtw6p5gWvWLmvq2vGeUVR9EHxAqnlof4XP6O04hBTTju2f9E4VzjI8UoQVdwMOO5FLoFZgkC8
gFYMYt0+idb9Ebxiu1TFU9sly9yLoJh+Mab5yGmzvGGTAOeG+4Wb1LZKLApzR/Egyzj+aNtcxAdg
OykBEzDHznSXH8HK5o2SWqiYAUUPTJ3KRPovJKLI+qcQBCv+YSDp1Hz9Pz2nsEY1uqFbn66bVW7S
L3hX773TUUPkm+5FKkXk2GW9S0yXR4IcCd51qANEd6Wzq5tXgQZI0WcqCQ9tYvJQ5tIDkmqBRoDN
WTbf7oYlrDxhl8aSGwDqNA6vu7gtOoDFN5xQbi7DcXLUSH+EfU4hDhpq6LZX1aSBHGUzRfwfCQrd
HgYTfKz+hS2XiFEMoBH9sW6rgGNiI9TV4rW11KjgIx5LtezNQ82XSsgaUkIRTHTVz3evlw9E6XFz
PtcfE1Zbngne05Y4p6z2lzZnE3en1gNQ2oxzKvIblG7rPzQi3vccTY5UxVnBfbpiQ0ukwiGGzzhG
CONCpWzB8v1JKiVfb0poa1AWU1wUNM+AoQYxCMFQCXIeYn73z+Ra+kY6dxMTlIbrgX3lW13FVLJd
J2sgTMxYvHwRA+UMvKUnWvGL/N7/rmQ8ZjcxPMQJHfnfm/mzySfsgoEakJDR3NCkmaLRO3Xdxc9j
frXOtMOhMW/SesNJ4UxU4wmGb4GuTL3aQVx4rY73Swu2vqjnK8iFCfwAEO21xGlU0C9+H5aYqmO4
K5drzebjXKoX2tPdmxvQB4vQkAfdqHCXVECjmIUpmJu+VV/8Fbm4Ao9uDfcBB1ASk7jnCZqHjyot
p5shi7VI+ey3+sEUC49xpbsj6PrOiLZJG1qSjPQYFG4nAWDI4GGXlNc5CNLCP99SZzdEmaQlRMTr
8OJ1aJS4KroIo48tCToq8TrNIQvrjP+EYS5EKNBhwBSWy607F58UfZrGgEM2hLBF5cRuXzdH7ZxT
NY8il8FKIr5wiodWf+/EGcEXFeIvcR6E3Pc8eZJSC1bThP1jDrv0r7+cPo50ciEofT0MHR32gKnr
DikDDGwyocBcse2OePNI571DHFJ3satusvbWUSiiu5pBWDKrffXXLAaCVTmeH5nhnebdVxsXNfa0
deXV5U/DSu1LOtP++8l3dy75heruLjhTVwnv37j10QVs/qYWSF5b/ZNv/LSg6fzVzqGxG0mfxm/r
2CRrzucebEpfbcdJ6Dq+N6oalhKTQERJEzFJ9q7+fEAP6aDUeILyNEO9KGj4PqUXbvgatfQKGIMG
/0xx0H1vSEfxTbIt5wY1Ih2s9717SfvU5+t+EkobYVhCyyhbaakl4oqv3RlZYWWzsDLrb9NvsP5J
nX3i4yMlj51tixVLvkbiq4oXJf+8seaTGc5uBQ1L41gxAJdyQT6wF/UOiOkB1LMMdAZ+NzzgHVxh
V8Yq/QFwpZOumTLtvvKWKdBtjHh8BChf6w+68BOXeokmfsNjNufBS8jS5YhkH5f/ihqoHYab95sq
Lxv1XSplJsqsBBdx35cqoysVNNyLEZYGdGDdxEC6RRUIRJ9rzxb0xGMOMDnN+LIQDoAYBgOwPom8
fvHvFn0XiUCeM3LQrJzKyMlYIhHwpHfQqXiuMsuoo2/6kAY8kcClLGsFOTqXZykj2HVTqAm8gC5Q
hixMshX7yDv3NSgKyMRUHm0l72SKkLdP5UQdfxncC7iWKkdwivKHXx4RtyC4QoWQlJBXs6oGN1qe
FC2qmcPFtgCNZfrJvVxrV+mWkifMbT/Uyvy7esOoKTCl0hTn5CunovYN0F8KgOhNixnXYriw3uPF
k2A4ItjxORpJ85MKmYzdbTFzUfvRnbytzfUUV0sE9i6PID4gH2iIQrsLVO6ABM958oKA8sCmBFhH
ZTi5NX1ZY8Y+vSuGolZ6E6G0JQvSngTxPbK90B1WjSuTfL0CvyNlJdmv5qxSK9S8xla92IpW0muP
57/BI78MH/fSVp7MBKXUZcDP+Y+K+7AOtQgeanqqgkD48CjaUn/bkMoFMCUzimpzzH2wDzwNC22M
WUloUytFEzOg3XoKi/B3g8U305XgmOsewDVBSS03PyPq7A/mrH5afmHdrlrJyZNlHJjKWJ79CTJ2
7ALsBf8T4DoP1e/A5L4avrI73+7tnoAzPjeuVhx3QjRHYgV6RYEmaPWH//2u4VNXlqNeCl2sN0h0
AJ2uB8v8c1Shiu0CTPQ7qnqjBEassg0rjJKziBBjgMthjlLrqXa0/xHDP0UiZD7eA+OHE4YsA6VG
M05LLE/y5aMud0qmNavgSbxxV7wHwsK/F0U0FhjicB0x0b7sbJAl1TU5n2adcyzz+jUN1uNAAs09
kcFHWbg54qK5CXQt+t5bnF3wMFKoiJy7HaqgS63d/OcvXuAHWX7uKISLrDdZJa1fXXwYIJw+crR2
NCpYUdhbozxJJEG3cglTcTwUq2o/xIynpXe+nWkwDtDVoIxQvya5uQ2K8JUZp4vrD9uZN9wQDwvu
N/f9M/L23JruVBxXq8PBIRCkjMygX2iMkicOSHTOzSVcRavaAHeTbAadc5SHm9ERaMXvaN8mvS+G
vpLyJIk0uMZVRJ54pg2erNCgmesa8BkA65ayIgxQrVe1+1+uvbpH5N9LGxxBrWazVz5DlFSeDzVO
5spnsOwfqt8yTg9SH4pmIrHxcCMQy8196JLchqp0Tk0CueWbg/UkuXpzFmEOo7L+3QColYQgDbZm
RW0Tup1KcsUQp7Jsld+/9r32S0o+q0qPhwbtzlmVizYAy9JUtdyNubZCBJ3c1bAtJ5daVtV1uUS4
yFsMk9Bdz/p8IJRTuOS1eH9y72x6cATXuavfIaEmb47FoOifnOIUJHN9MhH3s7W/FnlzfX8+lFq8
GgGoT0BPKgAB11cG3ujy2BCapfnsAWA4IW1WUg7+i3AW9HO1vg7zrNt+F7B5KXhLjyLXygo6lvaA
lNQ7JjtVSufNJiTbLwY7vf3Uflcqb60dmpCBAP88qmSz2Ll/Y0hRBPrcUJ7505zUwTpCleuXTGx9
REsjGntxz0/U0KL4cpi4uhjGillpSP09Egr+KPr6nvafX3QzDPsX1JKT8KhjMvSL3Igm+UCsYSMh
bcJOc2JasiOn337tmDdfh3HhQIZf+a8u8Ckb1sZ0Ey8m6ja0eLCpBmiuW6wVbWs73PAI4T9WmKy1
g4YbxUbK/lctPPNcOxEJlaXZDY79qNHO3fczF409h44NPilDLs7NqohIjqwj1MV/AChNQZ/NasHT
yMIxVP0vgGjlIJ1j5ffeQXutwTwJN1D5Z1/0CS18FxMp6cMtSLW5q7sjjFDb0p9KsoPTJsTX1sXs
cRehRnqXlmjwjfmZEiANXIUoCXzMD11y5PUe+V8XUh5VxX3uTohunKCZI/EI+5L636ovTVq4Uhmg
uB0xVQOi+0DKLie0z1GGeRrjuXHQLVEJvlmziuBLAf6hsp+AH3KVtlqkGmRDIr/Ju/jlSpMh1CKF
3k/pHjh6G5Dl42yDvTpcqtMIb/d1wzrVLvh4u66IfDAntSB1bjJZPc6MUzFwriAZSgW59jLsRYdU
JEQC4g75iot9uJYSG2TUjObr8mIcUEfdaUG6P6ed5llkrmTXs+VB9nVV9BmZ9zLXYDBIlG0qy2XW
FnxtJX8UI+YmpixCc4XueFTGRvAocmXcBA+jj2fsPvS7YA8fSW0FPTN3zEuRy8UoG6U0QaMi3zvN
Zqpu1t+s7D4XS5cGkUvQALmaKEqS3NU6heADrooIN6aZjy1WLsTjj7pDq0EPkwHFIMifwHaB/vZ8
woc6WSPRVPKxGjyuYLsN1xV2Ha6FL5ZSTqDdjOLPh7uIXhZxAi04mplx4jA4czXB3OU18PHGOXdI
Yxi4OsXP1VpfM7UUtUvH7OSPYOvmOttH//3xG2PsjfleJTtJCOchxXnqbvONJF39A2rHWVNsd+dq
rk8W1ooK9GhuqlDXbur2vg2UT7eJ/puPg6Znef4HN/raNMaD0wbNkvJLwEUPdmMgrg0BPvQ/1sLj
c9RnELijVMwGAvzSS+xjWw4ZmdZaGLi9jTkkGsBU1Y/HALwm5gyg5dcesuWS9WoON9R5T9RtQR7K
dpBfz3BQs/NG1G/Sa8yCdW6GIG+gTX5qDt60H9JDYGAdnw5JlXH8YcCbeu0f9/3vg1AHndKLx8YU
bP0WQq5LAeREzM2WMweazFjgfjW8DA+vZ6Q4M6tFDBM0wRi791Cw4Nx0rxgGPR6y9IxAqRfXh4E4
NvKbb87r5KWiB6DAHbgd6xYvkMPQ/MTz706YUGjrmIsQZSWKPXHdzHjU7cmcr6x0pvAFZfKxq+as
VpgTdFy98/PaIHcXBB515e3EP9CDo30t7aqnrzLAoMszSfH2OwXcnknVlpoAatNjfKFA8sv1NnG9
yXs3dC8owkowvPtPAYZ4+NGw2EDj8xjEKb5P5tePv2oNwerU9C7E+rbLZvPKlk9P+7OX2BU+oruO
t1dPt8yl/wLcsSwsb0xjfItTtpxRCl8Ix8NCmSWDEJ1V0gCfCt99fm1U8hQIkc6rPAhmgYO+NAj+
yb2su+LglgEon4ZmrKK/QqwH8K0X8L0PW19y07vPDhci2MAjXT7WVxNBojfKKOkJXezPz/FBegIz
q+TFnXbknB4OdCUPo2VixSStWfK4hQsgSbWBU7+L+Hl9JHKYQvDO6oZdGlkPtcdyGwhp1eFY+yJo
WPxQ5xdZx4Go47H2GoHbnkbqcako/jPr4baJ3Ztn3EkgtOqdfShr9LtMnerzisSLWKmYr7myfd6L
rj8w/QjjbmdRQJJHJfg+oQtXfDKHMwv2hEdnSLxJ0lKo6UUDd055n54uUGgbQBfPc4hLiTCf1g3S
y55/3zQLdpGzKWfIXXL5BLFzZHVM95kGY++psOmTBaYt1zXwaPesu9OeDNyHNRgWx7Yoy51vu2Xt
vH1pIUrem4OMMddXVOvDICqJb+Mi4UNSuj7EvS83OCCQfCHW7JCn6cl9MeUXfai7Hk/uAW156v7z
cQLWuhEr7xxcOdm/q0deCrM7+PVCFafFOhOdzU5psHkm2K3flFvOooLS+yTyJDH4GyEcen3kPm8I
oJ8fJiubPl2zD6PF3x9Xz/PE8z6De83bRo2FPpkgEQ8v7AyIp55zc/nwsVqxWFqFhmjcGIXXjoV7
nw8mQTqg4sX4jYQUGNn5j08U9rbWoSkhoyKTyWQwep1iVEuA9E3dqWS+UuiT3TyZo//WJTk5hoIO
OYH/k+Iw8u/j17dDEu5V6qQPgtmHtRrtjBgeIUV6lPV+MqQSNrjlhxRCSY1goKRSMSaoQc5BEDmd
BEyTVkm9OBGyr2lV8M5xblymOmWJRx/8Ru5jbOOOw89Es2/jVxrEMV5X5EwlVJgzAom4N09hlgLg
GbQoIbk03Keg3WZ3bKW85ZZm+maeSGJVDDeZ4gLo05F8mW5BVjO1md0UuRcLPrjZfLlnJK5f6lNz
d4JYM3bFtS2rdpl1CBryt2+MYFVO/A8gmIUgAnITp29EoykKSYNkW2tacRpltVai5fnIGlB+BLRj
UE897f80BAQuSBlEcnlwXUCdluwwz2W8iWLfDpSePa78W0RqBm1CIBhWf9kBOxd2y0HS0rjeBOHI
Bf4DDU9ocCubq6NWSzwYeJHHn/aozGfw3MDZqHF1edqVeyvMQgyIegiJ7wqgRTREoDz/4UdP9J81
evEzAsof0GYMyiT+uxplRv2xsbPlHQH2Zk7PH5eu+6UbKSdy9iHbQm1GR2wQJg9bIh+zn/Mc9Qt1
2AzoJ9tAgQB0+LfVO775Z5YPssGrOU+RA7a0pzjXb0EJEzktRR01Gce5WTesD+i0NeJCwuizgySs
8EHtW2nGjuiGfHFaocFu7TelMGxaTH9LnQUIsC2T9gFYsJwr/ipf7fEbyy6CxwoHjHMJtEUT5Ge1
ErwTPltr0vly/XLE7ILA1Y0Xa/w1vW+2JxT7u86WuHNjTLGHuZikuwKzVt8zK/5881cfbHESjE+X
OgduYInPEP373XSw1s5yU48/XLEjLV+idWHX0T7XgVU5muhRX3Vvwz1n6jnKbgMVb0xTq6G03t3w
E6Ael/Pd/P9dWo8HlSdjaFwY6ySRe40CczwWASLIXDG7+AWdVldHak8M3g+vZE7qo10GkGPwGo66
pmkmBOw7NUMk88YZhD8ZNwTNuBIdyyEKI53jrEcgAiTeNkWclENUZKdhX7QPhok5Yi+kQD9keKz0
4ynGS2hizmuLMfyjVALJCaSAREmIzg+Ttd7SO05tBFWgfikuy/WXX8doKxcbLRv2F1suTkNQ1/TY
UrwdF+lMcBgIlcXEpw5Klc4KhLjAeUjl1SjDdWyGPtlNil2Xd7qtZiFbHaVpzn5TD/KEIgF+pBtk
zX6OBg8JYdRq72cnE7Gf+J2h0KGHOjsTHnxYXJDEFa2+6TfMMPP3PJId7vrGx8iigkNv7m5mIH7V
jXVKGFLo7DWBz4gtNcnVKKm6Ahvu/E4uq65uhI6o54ox/3ve7s7emLGDhTuTh1jHEfdOcuFJXN24
vbymgaoOeWiblWm9Wvlz8b6s6lB1FLAhzIcX08sMzFFpiwoMDBVWm+wHtf4m1xRR+eQtaUE7MVF2
U34V97Y5oX6ixi6Cxe1Ci2d976IfmMKOrmZQXgAiL1vsEzDzygND+ErQj4kwxLYVkHQrqSs6iKmG
y7drRMdFHi6XdEE5JpXpkiRYt6w7HliN4T0nPK0vIlvkio8s+TQspf4zI9qbr8xbpKNIRACyy94f
LPFiJtViR2E8utTBI0I4FTB18k9RR74UjpI40NeTHRdU5GzQae3bQiel9ugWo5UZpnyv4qdxfKuv
t8flF4fKEWKDhJVNi8oRmTmla0LkeFgFmh7QPUFLWT0qm3nwHIvJ+R23o2KaiGKwRc5Il1+eT8ur
PwCkJwnTXAUwUDUaxtfAf3f50dZ6+5W7ojGpiu9gzVdQXIUZPKY++5EkNJFc3cJpBo+KxP88sUdu
QS0FHGCh/16Bg3bTvrJJdsms2kYPisHAGr8dqNprpUfDBFjqQcc+me4njhhZdIBXDCMHfV3Pypna
DSRO9W7DW9s83p0H3mRnDe7cxrJ7jZV6lHDKo8G+t311B5q2Rs8h8IQ9QjgrjAGjd+PBB7SAKe83
aaW0TgPE+pmXrUB1dsRqP58qPqDHoFzBcsdOsIN32SyNs06g/rP8YoYha6+DLWDpXDcMCY4xkcxS
eDA7rsJQ/atbrmNEcB7pw5c+DwhLW2uqC6jjn0ODxpr00XnZfRKSJneK+o4s4cEFXUS2CtCfmpNY
eO56RbZB19tvRxXPT/LTp4VbUT/9ttTHx1Rz40t9COzDRSsUg54/HkDvsa9JmUWiviydm8y6xBWc
or4qVHK1tocjdSjZreUP/0LXiM0N/vOi2VmudkcCp/NEUjeC0UQRQMaiEIo5WdOAQty218GlOyJl
1wdQTECpysbbM2W2rn8IbhlH3OhdeUhjphU2Y3BqJ0VvajM6pzkxWpJFbxhJA2iH3DB379q7Ms/d
fmYj4ed38z0L+OtpW05R7ovJIazZwFvdo+M3XySS8zE7xy3eSUcgNOhzoYJFzyWMtX21TH+FTKzq
ckK4P2vuC1mcKUhCmbp7qx5H8PpFtXbcxteYZVWQMzxIcoDlFA8cvesxiP7kDVP6wq7Jsi7Y3Wif
oUbUVUWxn/Tn320cQp84D51i7BMACoqCamUKuakcnta0qaLxj/uO6LaGtJYTd8wPiIvaxVoaMlqe
JT8l/OWNNb6dUhpomO3+GUeknOpNgXg707VA+yevBvVVxy24JBodvY5oTPlE863c4syZhwUasNrm
epKJxwa8btrkAUFF/PUffFdtuWnkaAFErNhSNrCnrKTS7K4PdRLIEF7pOAVj5F3OQ08o5dmWZgHe
kP9Kq4O0A+rn3fqUlJsh/MGin8W2FHXiQf8eyFbnNpYzon2s7RJYO5I1WEL5GVaipluo+6yJiKOT
lAFv+sKVGvWFAD36pWUv75YG5dGJ/Am599eEQbWhlkEl0iopdVNClgBe+fOZt2l4WaaJBstNm/UT
xAU8/mru8tv+OLv1Yku5pwYIUA99JJxL5TkjvP+l9YH7/RHEKWIy70OYUdMB2tkQZipaj4RGHNkY
0ZUQ3eqIWbRvosB4D8Wn0aWp8eCqebVkLXCA9hwGZA+XE8WFnU85PIcLt9XgKfzldD+c/yRA9bVN
Tu7qLFD/obvca1dWXj3lx8fKTV5YXnGmBPtc/U5+5FLRCXvQR5YMv9dUqWb/OqiV4S8U4gukqZ/0
mWAeihsHlvYTsv0+MS4HFv/mQN+D43gcRxxODhkvOKihWB/jI6DxhkwTKWozPRJrbVlYfjXWNXF0
Ivpi3WYKcMTmNAt1KRZz4RHg4eKnn9jp0574Rm6UtaoYYk5NyrW7yjxW+mHjLmaal3722acBzt/2
ppiqfNbVu/6/8z3/FOMwWN1k2BQvi21PK8JM0bNBjl14CmbW80T3qhkoNlgN44NexH4fQGJ+ZaJy
1lPJI55guLxY+dllEyurbHgp8CYbjlVjdBp0bu+tqqPRKhUO8iWP78ZaqyjaIUWP8qfIUbKQeiHc
QMIAEl23VxDijWX7Siiipz0W/h9wB2aAXMIQOIICfxmEWP2/DAigf9KvQxTZKPFztZPFGIee8/Id
BnfoIb5HjRtXO9vdh/QZoSxcy5eOK2eFeR1z53n3l+WO3mEGdg6xVfpzEKT+n6hXhinvFPdDKBTt
GwDVUhnaY1YQADyP+SNbHBgVWRAgQdRkVHdM+Y135d75RhavRV9QDF0oT4gfLJ0Me8/QO6PuAPRT
8XaSYq0aniPYEtnWkMWKwEQwUC7Fz5X65PF9WYOI+Z/B5pSm8UJvypsDNA0SW9O79SA0n7GRMxnt
46J8miJqil5cyfC7sBaw/kcTEjse0jcWEI1qDdECpAkmyw7DvWiS0Ye++FunbtJNr10MR+t+S9oB
8qHNx/ug/yRXpIis/ZxeSO342hjwxywLwmImDU1IHR/tIgq9lPr+Hbdz+l0dr6wp7ObY9fAncwYx
Pap/5ndetZQqqPNesANvY82+/7cgWaqZpAf/rpVfoSNV1SffcQUpyiaYGguZacoP/VZ0bGJoc4n6
rHV2rghchCHYh5a4zMFeE7+IrdWJ898HCwNEz16t9nSuEJ6y8AjoyFDuXGXHTSk8x/9mv6DD0rLG
H2p7vhJM46FOZ3bElg7HTyrITnzOoA6A9ADrf7yJseNZ2y3XDIZ0LZyqGQeRXo5CxLU1NzgGhgg5
DdXkJX5Id+CYyjZE8hfGvpCl/1lMWfjTz/qLh7OOQ+Af1SP8sW/rP2o086K7UD640rpsg+YDleDA
C5K+aPUwGSb+1Sz0NxtMz3WD6sgXNBW6t3aNWY1RyGTnpHlKw0IvQ1ef9+Gj8rBla8na2X5PJaTv
0QMdK3/spBCOZaaE1JgcLYiEpe82hGW12hvNrrVbByhsDM1OJjkcO4ANYkScIu4EGp0bSna9JlL2
KiHLxc7nsHCFeKnR4urL+O6QBd6rPFdsr0QSWU698hT7dXJ4Gf7hSPNBa5RaAt3ECJctE3ZuYuhb
MxwuFKs09AMYnHLtGgbtmRHVF7aubxCEwPqD/hbDMasdW4Xk2J0AFdFZx4P3QNyfLg6YSdLr5Bnp
VQpL8PK/gdWvou2QQA35lX6Cnb2W06wGVy/CkBvNN2SP/M6Tl7ttcxlX1EikUHHkmgw6fzqTqzYK
2mFDi5xwxk8UPjiosYwAOUZBiW+Lbc2V8kyHkH1BHpMp9SCBd6zjVzYtg5myhDBnbdCRVOC2ZD0m
uZkVM3Fv+cUrLtiFfUy7eyMX/+XFevhWChm+kZNT/F0Tin5ZjfsiJYHBcc6g54mRAZyxMbm2RTUB
4a2UxI6DGRtMW9kiLydwRWPpY2n5vT8lSc627iMygA7XufszSiKzKGAf5PXBh8yDJ39uXuET0SDX
D5islDNloxPg7zRYoEFBMAM72wFT2s3ZGrNmUO9UcqG+y4o5eMRmI7u0w1TBHTAYPbErjsH2mLbF
AJ7MQg+m4Txvmg/ccltq97iYG0QKPYgkltigYxd6kx0eMRyfuZaPzpNrw7UsV30vroRYrzUIwCJV
Bg/jzTyiVIj8fgjEbQIHD7CdMG6FuVk/CWkQRn5dKOo+jb+mbk+kEbXObisorh9jacECdrIGumLx
LdpnzQ6MlV/5PUQMFqNojkNLy7mkHQdjfdoHPiRU0R+kCh8dslrDwJtphMS1kFiDJ7NWlqF8L5Or
uEt4qdegKrRvkDk7sADmZd6UbhDv81o7g5O0o9aYyIHSAwz/I58l3J4V/c5fPeby7QomLS8ZS4Es
rELL2BN9Fpangtz5lnK3od0BQLjoZYNn7NBL1XzBSWEEOkOZh8UcPymTMdUAN8oJLRupAvvQ/5Zn
IFI3XFUKIKqtirnWDJzqD8y8b28LwADBGwveaGtQVd2mioGTeqp9qb/cCGhJXgab0w5lRATwa3bQ
h52alTrkYXIGgPUMKk9ETxHAFqjJiMi7Fq/IE9ojXNU4c+TDq4X4/tXcxc2D0ObkJfHXQm2Bryc+
AJ2IFYSeOflRbZf4inbx1HRpJGug+tWRnxMuX0/FIUpfvyHsDd0u0NfBpsgdJHu/CyyA1zJ2cun2
FaX98Piyabk88gkrxFZ0+LOXxnBWCu32LenR3PFaQXRmW7ofoV33GpOWbKi4cLStKFW+qssuE1Oa
MkDzO6+ewjugNv7tOOqNlQcNTi57bx/1+a2+/p3+YjSzSDBNdkPKQKwRBqYNFM30JGpr1WrAi6Ia
7ZpLEyhCKF/W5IDPwZ0lXLThAiIQ36Io7nk/kV9S0giJp38dh/XaCA5rjoE26w3vVBZvX9LIaeBv
qBFZY6CnKv0xtUt34qcBGXa9Xa5FPWV9dtv/4NbngAHKwYg9B6Wvkno4VXDxIQCrLsATSzj1ONkL
Zk4hgqZcNHvYAwP9ZzCfOB1RKYQEGw28HdvliBL3QRxgrCrlTn/Y15PhgOJPb36ZIpXYtxGs7DpQ
imCMgLgiDSCC8D9dTvFHIyBnf/ANZuejd5cd0GODPZpfVpjKDk2CAuIYV6jfrD5/+Y+7G/UlHNaT
LNTizrMwi0G7TZ3z/6ceWj4YLnRNCLB7dRlsAaX6rJT+TE5m+Tlm4nWgmJIi05Si4MOaZrFAofnl
D7yW8LC0TtbGp1emBBaCFGM50uOuAUgQEdL/g1nUW/fT+WfvsTF2PKf/XK9PSTCD3kMC+DnG+Hkn
h36ssol9XQvNgkvX6Mc6QetiaK2IiqS69fUJ4fzQ3H+HYfPPCfquvAEBOStd0vRq0ziketIWbPRY
3msVRtwBDx5I7JyMDMghpW4vXU+m44bvjzYH5AofZu4MwYSOuObZJ5dTcLT4fFZ3f9pJ1fG7/oTs
afQ30k9bLkIJ2znoOCp1M3m8xi94xgRbzboP1GosXTK6zDugxnrcKJZandJeDKPhkzaL4CGxg90X
w040D+I13I7XHthR1/hZYpIiKBG7j41nPMcCJwSTih4f5pNXqZMF6El//8pdA2giQ04n1+zVA0k5
MrnRVu11um++Nu+Cb2V1TrVQ0CxwTZgIiqX1MqrTNkVh8Z9q6xE6LerRTfjlhaKkmr5FS+qKSB9H
3DRIgGAjx1HYBTonxz5hDvORHYLVTBRDgeIrOF8awMxLOPTRA/dsLvw9gVT3GRpmrM4xJpnj0tVy
CWk1Ds+Ql04zXZ1Q2GkapVvlNy1Q4YDJoCUxF/wzUEPJZJYOH0pDIEJe6SLP+ZWKWCojT4TRM76J
guaFrtLsvnhVZ91orsu901tvg8wKarMvQZ7Z0fIzPdc3QXhvQJWoNjACP+rKo9YUvzIGGblRZMRK
dbJvG4J8/FQrRvGwvLntk1Hqar6r2rn0r62xGp1QGv2+kCOLtTY0kclvpK9Yishw0cH/Xv/gC+uu
OrsIQ8XSYgz36v4GW9uFRv4Vy72iQSSY6TVqATT+L124eQVytvgvuQGfJX0XhnPEPnt4kC5sUHXQ
pFnhoM0D3Sbk2kwiy2OZ+4DoMmWzZ7rvOaqCTzvwHZXmn95QAP6ZU8fLUN6BLAxYXAOtBZ+86FCY
t/zzBFbkuSlpvvHfr5Aiu54Cj4JLL/m7mQc778kVfCwPYSlgfdW3cOsgOueEvk5ScMwhXulaXyCi
ljF/nf2MGTk2SGWPfH9C38ZcbBhvAJhd71fWIuGxL+n0JLOm2HftskRTyhdNnd2vjLX1gIB7WvFa
FdF4GXLCMKgkvnhWWnZSp6LNNUBUrk/KVXYtKOjLde0/Y3klYZGEsDLAMPLoyiGZ+qLI3nt+rkgT
J2OlcBGkv6sB1FS2NouJ7Pes+h2gsMKViLtu9Yf67r69czqAFEFsBgT7Q9zCZ2QiDqTsZqBDZc02
sJ9QpmhobT1BE6YuymUKgg+flpwu6xZY03XGCveH3Q/B53/U+F5UM1FST5qV0cN3lp2jxRVFDA9l
wQ7f/iNIcSCTsLxZGHDy+NsZ0px6k0LcfMukQCPwW2RwEArN/reuryt4CYvYwb6FJqYXZHji1R6f
kCapLxZI44lt2ql+KuOQv+bOWxTnKZbVZeTUCsFaw5yRv+rAWZ8mPWJWjG5Mts91568Ljr9m/t47
G3l7zoSP9ZAv/9Tln4RxBhxK3B9Q7fz7lbawCl4q6IVAZ+yACsyOe9ocISwB/prpEV0ryz7YUtqB
TL2xOGw/m04AigAaoOzFkt9aKSDpvWsbUmBkGRbJqXLPJXAnAeisT4prZZ0No2LolZb5H+vObNJP
tBFwWbOTQZKAEJCeb7dWeLomWqAae+r9h7UnL5G63QC1h17/ThnBqEt6IlvBVpx5ca1dh23EqXDp
lxjK4qPdZoF8ZqR/muvu7XlENw6p6MFEdLYKT/bb1TaXh8UZFe7/RzIIM/LLvwY0u8Ec3LTbWaU6
CRJlofTKK1GbRd42QvPeDAPssL0fg9X5VFgHJDnGgOI18EKznHcxxFc+7I13T1Wfi5Ma15KuRHr3
bMs2p5NFlhNqnWRxHwezKaAFrEakvr2TNIfMoQW1nVJ11efDRmnLDblp2Ij9zkoBsI8EtE5pgXzw
d1zLrjAeP8lNVeP3r+R7V6+Tu+PTZsUlxpH0mmOmG6d2D8PYr8nAXzYqgjIrxEG6jNsdAGLqUa9r
M3PNDv48IXBQS+UPUXSNHV1UqoXU6FbfqMT/I4mZ8UIuuA+k+VhpD2DkZ2Xi8Owlfw1e0rd2s5bQ
kb2dtwvMCCceG9taivoC04B0vyK7EWnjiok1bWWhcWbQBdhiYsML6Ly4Txdz00RI3h7ZjJjrvswT
cgWJXWkdraqnImnCA8hZOOzMyLlT5Kl4/Wi4NbEglduDlNTxXWU0GyQ4DBrNiXp6L72cvuNEW2kA
ItnhEwW8rtlnPaD3m/gUUikSe4MNwjWb1rNNS0mCOMh35l0yY/Y/AgmlEApg4SD5N2XXDLKDQFYR
SSW6GH3yU1VENkBRz1tkzlCis2df94av6UWnSBkqOCRiSgh+0E8OS3ok6D1S2SC4yI5f76xdoxDv
WD+1ByGziC6J7fkRMs6L4N/J27Hev8qJoGpxicp/GHwEFtKUdT8MGn/ZoV6wueP1BQa+DLk8/tQg
TebVylFyORjUALPO0EvpUNK8aFbBrVp6tr+FjGSObcjJFu4dHMw7ssKPF9hwZDh7JRny2uNi0rIu
sVZINVEYYvdtdOAjBn2Dh4hd3ouj3GRKLEFaUF+/pV30J77SfAQqnpbOFEHwBGfrCvLdTlnuHkKZ
1C+7BRZfX7lhMY2yxkXhHB10a+I5yRjI58vTF5IPL9O3HK8KYpPi6IH/rpa6a7qJD5COcUDkwq16
rJHQFww+BCfXNCIEcs3cg1UUraanIdhfWyF75X3bxnFJ9JIHkKuUxlEn/DHYpvq9AUVxVVV9GcDq
emR4UYMpn+e2eTVk2j3ouIXu3pdNGrKkWjY6Himgi1dCnIf9odJAtQn+DmpT3z3sqtadLuOht2jv
vx/b/7bRIMi63fkZKL4mUQ4zFLKWKRd8vAMH9KqvSHt1SwesETGSh6TaoCoETcdiyryrqPUhSN6Z
0WqUhZaq0VRWie1GqYzgp4y6XegdgkRlzkRlRIqWBnhHXh8TKAfeyV+CJlz80AKFYoh3KKHtIv/J
eIaufT3OTQoiwnAGVlOK8BKS2VfGbAmUNXF2BwRS+UW1jnxtFk0twPIsk7f+jlTOwCsSU4vC/qAF
Ml6BiFtynnPp6fDaTCmjXvV2QwGIjnzMEm2z90CIDE1I8HaHWJqYaS5/uBqMXyCKpyY67UIJo9mJ
+uQKt1CWAZtimpfP7Oo64gkTOxnWnA3XC4Er5vDmc68G7Z3zhcGrw8eeMfP4zmpLFi1Isz4peV65
pX1O/Qsr5OjOCCcU0gm2nlTiD0TY+Jy/id67pEVnD8IbkaIztvZJi+UP3RLuwa1SimujFpXecE9y
ID15LvpziOIEvl+HUUqZpl4n0+eMn6AjcDkM9J9divog5XrIBAbqcr3vYIL2O6ZUatyrvXXsF4oA
CczIQ9yaSNZlnOD2jm909bCOsSEtOyk9geXNDcO9Xa7xYT4VUOHlxv0WQjgREPbpQYkJ4RQJ6UqF
QC+ovKlmm4kAanU8CUx83UAq4hGCoHiHO9sjsqC5TygOkYV+3/LFMMUXkDyvTCqVzh7FWg3LUV86
OH5IQatpFORblJQdzk8CzZHAegY3wX8hwC2ZqZbewqgrUvPbAA4nY4Y1xnWtuL5hegxRMbWZ99bZ
mxL5wQz3Q1nFL3eFP46bYMUITZzfUJNfHx+1/ybd2Eo9zVcgWRPNpEwydeKbikdNOMnhYcngLggk
Lf9nhcwJbdSWFujsO9Tit2zJlVtGcznGlev4eeYFmJ2fe1eDainn0BPI5KS+JrU67mCqVbXM9DcL
socvIJh0BywVN+E4qjxy/rBCx8aqRope9OxUISj5KT/cTvFJN5ozcKPq/byaDAaiAg2Tgy7f3KYn
dEPBPKx84eoeiyuqDy4wLbTyG+5ikdGcWSdsgsy5cSJclU11eHf/HS28iZuqloO369S4JkDsXMyP
RhUFyQU0NZU2CAfCa0bRFXIoWONiMAskp2rfnMRt7ysjPbvr01+hm12fZbpmp7keyS1rAW9ONNvh
T+WcgC9IpRTmy8TzO2MkUdJcJckTuEBdhA5X/6RZ+Vc4pf8rK6EocHB2JwNytMcMY9DOP6ubC7nL
+TXcchDUdoZfG3c6lJIoyUkoysGu6zX0fklSVhkTBnl84OhhWwoB4YBdHF1HaVyFWMAAKP/E9H31
TmVWBAWxgOkzYFzChTXYi89uWPIpEVp4p1YhVGiuzNg+Ki7DlNj9LQhZ9cVpUY1e6YJQa6YwrxmG
/UDzy6AzTvc/UAPSwM+70Gp1+KVgSnPSMFDd1MXEmhNQuvCaLGGNO0wlHymf4DUQdvtn7VEu3e7Q
zoWOaN6an628I1z3Fssx2ej3ELkHKmEl9aGFPSWymstDBRHBY1/rnZ9AkYUUA4BE3zVwx4V+HfGv
+t07zc2i+ygmcVAAeqTe1zr/nuOloo2TA3JL4UP1jBYxxZhMlDG+ubyyh1oDeADfMTQcHm8HQxQH
qmXD7XFgz5rcEZwAYzvpU79NygPgPUQss+Y2iRbIvS7hQjNKAld12ZkSpUuExSuwF7oCz0iOmuQp
LdGi+nXV3de2F9xuN8b0ylI8uJpsvfhHue13hPXLrAK2+vVvV0zSnG5BW0RjbQao97ZVrWk/Ck7l
GZgygQUnFZSL48dKXRNNBPiXGgz+EjaMwn/qHwHL/HWfPnO9aBzIxPEETdOBvl5vd6oumxWXF2I3
5vKYyGln2SF3rba35gIMDNVztqlfhuv0mlQ6aiwKtMXzArtvAh2VVHtN4uE1RCzqHpPEC4KkTxWu
N34seWZBu3PJHX5vM2tI+X15l7DBPgJLYrB2Z5jVwsKKX6+hdEWzzww5Q0uj9RUsvU8876lJrPrS
iPCU/Yhwzv2qxTVY47ghH85KQTsq6WOOyU7ML4hoOr3wHEgQxQr81rzjJCkkSUBSjQAcMA7OEzvP
G4PgRj3LEYNvWz9aPXrJlf2qMjMB+NEqjbPnA3crh2XpMmOHCDyH3671FhYqA7ec4CkNjbdzic7f
if2RUbshlNusKgzjHljn2gQy3uHkL4l3jqjpqOslX5eEGuWRbYXirojr988wHZ1H/0Gt63YVKJ7B
P4uJPgEM3xDoik4lUKGYOkL6LncMpP2aYm6Da9BvcTG2IaKqnmHYvecKA2QvjJzSw/aS/qlaRt1m
mz+ALWj4l2psk7ycaQNoc31wQKhNNRQc+HAqYy+8JC7/vjgLQPrdtdkldm+NidU9kcLhXg7qvoGG
1XQXtHGnPmd1+dpfLzkk9taXvj+oycIy+PUKvJ3xanpQ/QN2B9E8Uzbvsm9BLlQ3fI58PKkuBgzS
tYOE2sFZeGs2gyczO8CyQsU8GPpmeAhxDmUTZ9G0vhWa4gWJJN2SK7EBJByMl9r1PSmUKFBqhRLC
3r5sDUlza4NLZq1LwV+eGHp2B1bDr1E11Gd19g2DEyKsbuLvbGczSlBFfYGm/8bezfJ5UzsPq9gq
QqUi1f24T0wclZrU0MU4UBluKSICEWixKcXdGwnheh8WMHO59mOClRGrVs0bgVfgcCO1ynzcOQyD
mNfymG5Cu4E9IgrOEPukHRcH9YD9MT6gCIo7FZhbV222lyZ4d/y9j8WSTCK7lAVxk2h4zi3Nqei4
zxG5rowBHnT1GZ31LrsHcy1kme5LkK3SnumwfHE1wgfz24pPaBpwprDbvPvx2hdE7ArAOHKylOtd
GfLzhlvsxInnrxj2Afu8E0tMmIljMpu81Xdwrth01kn2t/BeCSKVRzgwM0zCZbEjjd8UBWS4rkoj
UMfdsNQWBWVpGguhqXK+ulAw/vnfJdISr4Y4hsYpC1dOOgU8EoSyesqLfCTO33lT2/mAI0j3sS3g
4YsuuvFmrI58DhxRY10Zk/krNGU/J+62zfe4+ir65GvhhJNNMHGK92C4BZ8YGHoTtLrZ55FgkkZs
01PWxniYofmeXy2K/uL42Uigld/4888zr5vgOfYTDjRLkdxBRxPN9ozkm+TPe1GKBKtLt8FDmt4J
EHzCF5830OSGkcqiSoCiTNHWMYGZC7sLjawvXqVt7vmalB2Ts+MIP/lOjJL39/lKVNgdJt6gXjMu
oZsJ+Qdr9jz+UVvwEcof4O/GPrEeZnPtSQsrRy9i5WtH63PKdRK1EPY8710B1iKylXIp9uADhi4w
SvuREEuBLFiwHaJh8eiY9n21TXyFU0z5kCmVVjaFTU/6EK1H6jxw4FjWldSAnS0p0OcxYmYMbHUB
4I/r/SF5FOvBltft0LQkWN9lJepIfO/cPKJNolWQkUsef2nszPhaGUkWkI2HSr14dRWM1cOQMSXm
asYzFIXzczVHofzmS8CftO4xfBRB+wxMxmd7Kv4nQ+IVInITn2T/BOXgKGHUCtVnv5ZxqNJWL5zF
AhQWCbc9I0757SmjohydzpOCA5zC7leEXn24vG4kVxWecjfd45jevzg6yeFcYSmUTcElooGqGT8Y
O4+1By/LZhFfq3hgXsvE/wGQUrG/TILxOBaewAJobaS4kFjsWOI5M5lcuUNbN+djOGHA+S25EH14
HACR1lmsOoKGporJQzVkxfC31PaBAihDuQOV0Bt1N5mzf04npY4UOoZznN1Ok57qK2aK14t9fKTW
H5t3KnA10EGq5HG3Uj20ihoA1JuLGwZN3tMvlvQnsX4QOk1/K+rfK2tqIPiWK0DRj19yjINb6cPK
rbwqPaOhcuZT9OdqsSlo4Zv9nKaKI4EAcU0nwU48w4OHkw1u+1SIrqLVGaU8sr3KlqTnNCV1Sp4g
VH4GY150Q00z250J3guH+AsGNJE0HoGFWZAVznEKcSaKwp/T+GiZIurti4aneIZVsbOxmy85r6Uj
0zqPGwtQ698vehLEXhNLKQ0wDGnYlzpeCR73AbDZyK0rLmWJ6i2EeVpPsfN9opCTzvmsSc7ZDiHU
OW3ggcDOk4ZqZgmYy5KK9gqu+1T+rDgzYjEtTFXl5+rkz2+gC4027Nb3h4JrYrvTkE2XkdlQE1Pr
hDPYo09V7Itq2n1JrEmdSSNGUowDiMdwQhCoug0dHP4PLoloaHHNVnhpOv+sBaUkqa/+VBeRRgZn
+jFYF8C4GJhsAW9aKqrVykTaFdOUzvAa79oe1Hm7mZV50Lgk4Na+cOc9y2SyjYb0dOEHSc/paJJ+
6Y5r8RXuNjjuTB6pf6lwoMDo5vpS427KIFFYuIv8r9PdqS+cFGCb+2jv+8O71TfaNCwrlr0B/Rkw
sXmCn23xST0QTXnFD0Nv0IA13Uos0NYYQjbYOwasz5ZwLWIbuPDVLWhYsjTONcjuMhI5KeFhmIAh
HgiYmsaQBomU1FFGR1UKT1M7Qqe4xi34RVmrjJnmnLGRFT/p/3luZmRPkFnvDTxG1A6GfsoQcYrI
pYF8dAaF4/pgIOPXguddyyb09LL7VD2ybTxx8KZbXeSkSR3TF6PgCS1Y69VLKUCXmwnRCTEK/I43
S+Nj2yaGbKS69ZSfoJ72DzVzM756o6TdwLQaShTKcuerfr1pjaVCNZULICbgK98RmWiwKvKpwnKG
Rgria8E+HmVQ56jLVw5WaI+5CIYAkO8W85Y7w8+lT5dzF9OViywZbSCVMsR57cbSIulFFTVtFLlk
X9BKwQ1NyZ7u9AGqPe72ybwT7XYGfMlYl1wHFZ8j16MVIVmF+t5bQbsrwEH+XRC90nDkB8fvxd9q
m3rzVNz8kKRzVoaI4gxHAxA9ShZX9eeC2FXUjEVqk8xMKs7nsPxKc0FkYjjpKMMggnUWGitQpz8v
wUk5rc24MlCRxSpvgZDCzs2PMtkesEglxznMTFFyPs2Z9JIMmA9QHFhftxzLS2mrRKSEzUC9F+Af
X0+9hW7wFT6wwet1x7dr8DOUEwprQQlkJhbAlDmeSYnjajjbsw7dqHNAARHV9BZ1gYOCgLkulEjk
z27W0339HyWhla3Wq5BaqvGp3HQziA0utsZg6caszwmUAW2O8jlXr1KOX6oYVAr3WIOsoGgPGjOW
9fedEi8/WYzdIHQTP1uENr8B+bcGfFkfF1zxX03fzIYm1PfAPuG1sVf0eKOM8WaINvcYWPtghUW6
tZCX/YnFKtQoiA3us/l0fV8FkOljqW1hxLnC90NB/IyrlSlu9tzObsXAso5ZzUFEWPfHuATdOrOl
vHQtaaD1BdfX8HE/N4RpbdaMq2r0Bqy5VgdOTooFWUmgH84icV24vjFmrgz8+7VGaE1H6G8xgk+D
Tyi4JXiHaQNmlNpk0L3UjwwwyofpowO7MJxPK1feHm/9laIuRfW1dOL7g8NSwm0f5D4zhOnFE5YA
+N5A/8E1uhvNkeUzNsK7yPwPAcolWM0dm9PlNREstYMZtY41pW4OzmnCgduJAN1YEGxqQQDnE8Rc
Vx5ka0udHP6uYhkBwDp3UJFXOj5biLOsP0vX+/NSmPxMSsSa1Q8l/eOH2Cin3+fVKn8GzDHaMShp
Y/+sDTFHQMfJ6H8OSFJ8V2BiB+eXXMJyTJHLlWYjBvzvpV78nyMql71UiNEJdIJjB90xYKGK79W6
cByqcnlAYKiRkvCrkhcWak2WwWrpZydaF3S2WaSyajIMjKPoJb0IUrx2m1zz4tukeJw7uCVpa/T1
gH1WMa4PxTfQi23x2KXvmeIjsCqOdiJURQ3aiMHGNnQXSgNiBYjAimEtRD+RiFVqdYBCSBWJime2
JrvNiYEhviQWa6YstUifmTk6tT66e+taiJgFq+Pto3lcsyq0MMv+1XeV0uMsAzcJ2/p/L48UGtQa
XTomc2tpn0zsrIIoEy9NL7yuAEbRmPUBPswaH+rTP3xKxjaG8xYPtQffi0LTBb6iil1plI8eYoMX
/IXmJXic+kjPflYx0MqtnPwSIEZ5cO/h8OKygPSjF7OaE3qhV5P2k7GqT3qwMsV8TM0k1UFOdItB
+ArvaPRb135tbHPyLk6lux2pk58u5aK80gw1iyFIqsl6zeHHh/yRyuV4yRDNsAiyXAoW0pPAgMKn
obuP4KuvFIbb4cxWOsNcGoEwaHAbvWdUd7PVpnyvQXRJQSC5oTSjd24X+KIdV5D4csQ0PVS09iyj
rJA8+qFjnbXHxm2UzsfMU3e7AV0c4SE+HC/gkOJYPB1A5azIrj++g2UuFvxOhAd8av3R3n8sbFvK
z3RUaeqbLptxCTte1IqlB1sOY85BDgh5+1VcyGw9wI6cS/L1UlDcXfRKfCGGyaWDSe6hMVJ/heyV
u1vgTWnjvMoJuzTmasRZr2RVE3NCsFVSvsr9Xvi7ADXJl3tccwiwqHMepWIOt3wtdIlGxwfHA72K
pDZu5nrqFQyTh5z08tcYCDRse55FW59LmuL2R/VxtvHs7vLg//N1FtQTZHfeOK7N1rANqfI/HLKz
uNLsd1EP4aKYKm26bnsZEQDx9mzrYiF6W07PQtYK78HfE0GYwnRpxrORW9OzC+m9BFPIcEEJugf2
dbhqcWtCFGVePAa4N5OAP3k/7PESXN7xWTUDuWzYQ3aTLJp7lwlPCvwS5HVTjmXkRz3iI5E/tlfq
pRqg7E1dIjiRWI0rUbSYOoQuqdXt998PB6XB5f7NUGRxgCr6A4P2VSFqKeozMUGZ309ilw2U15Xo
bFj6hQwRJh/O8TREa3S5b5SWjaw/T/diVNWVtpvfiosTBeyltLCYWUVix+LhVnE6gsNm0efa4T1N
DOk/Her1f8C9X0FSRTGQqRZjNtCrCQjdw7pQuXl/rfr2mf4Ef/X6xe6xonquYcMFxLKmxQN/LbdP
A0xfr/Ai4nkgdFMu+gfC1QkOCZFAUc1emxLJO1HFc7bb9L3vVLuKo87C7z388d8xBwalqiOPKP1K
Xh1yaPTYah13o08vTzIUIubFNjlK8dXHMqA5QQtlYYz30AiR2sVWsN0wD2dJzpZuwO6yKC4eco8u
pdpAnHn8/puXwCOjZn/eZ3+/uQjbJuHCP8PP2NB8jblI6yZjugqf79XBOFdXWUr6o1U5qCKArk+g
JPf6qjcw8Yfb419jFYAF0SMKD7w4lvXTl1jFwS+eGdtvIk45fZV4y13TH6kTOk4z2knyoVqsd++0
UNKKmoHW2lS/pUWHeJL+FJIk1iKKicKN4BnwqOWOFigqq/sRn/mZX9gm4qa+Y/ttSrHX4yrGh4us
f3P81dDT60lUAJvfjtzhYcYUq7hGPMvV+qsoMTH45tEceyCF8cgnoH9c6hWEp5bp863xkSWxLrb/
E2+hthoc0YrzTkhjhgfKh9kCesONaQVgUkASXagIOhbHNP8hM0KRhkiVGHLEMySFOrRBDImC0GSU
T/zG0EUmiRw4ZCPQac/7J/ooIDuZqRDe9ReKvCYnMyx9JtzdcNHjNTgPWwfMZqq8RbHKwDzKRKBV
GPGvEK9Z4Sn/LOT5z0UARTLlpuKnmtOk/xCCoURsY/6g/Q5vYFIYJtgI9CoKOgd+0Kayfw9qanF8
E8KQSK3Wxukjw/ZH22SKjzbwifHoTuVFVT4VR91jXcKEokqaifJo/uDqqI0kh/0F7zw7DaMnH9od
Rhsm6qz8OtaXkXsyaernW+/1ZqFnpaUds7m/HS/DCrvG7psSCpwd/9hOHC7VRAP0vUStuy827+ED
UrJBnwOliMdzIg7Bg5R9UfKTvKdTmqbEj751mPUu5jNn1WjGN2T2RTbOy6Q2ioRujgaXhfyJrPud
EQdNo42LGVWz2kayRhqe1InZlgmwOmAfKTC+Bz5klOxJg73Z/sj+N3/J38itUGJg0VBj0dxsiZSx
JuhOM45t1MFZZQ3eB7nt4QvE1Hl+IpbUmzcpV6Q/4S+YNf1mOtJsuxRsyt8fMorG7Fg+STiEBaR6
blK0XppWq1pA69Y9Jq1L7d2mxLdXJUTpeNE3QivjoT6pD8If5Tt63Jxzby4vNB9PtNTNDcEcMumN
fqwV0OZlZqewBbi3Hpa5OMBiWDL10EJOTJ5EQ3hva0ZlSJj9SDsd5vd0WwYV7A+8dHH+jwZi+KXi
QtXFQJcNN8fnDThxNqDvm+dpIMuXQsP0R5f44Acm/E2LBW+SnM2YkPilIjGta9Vf23paQ+/OyncB
xNCA5OvVQGDk3tduQrkI1wYC9SyqM9sLVn1vBvqpg+i4CuCCJAcQLHn0RXkE4etlYgrJ7MWn1J/b
r9+ECxectE51PxcxpAwAnco6mEXRS8N0lFrUexHgdipBu5xPlcM3v4wRrPcoFlxcbLHyVIV8F5o1
lWZpqJHAHEjuTq6HIv7whLBe0ZHepxXim0SrVkWAa+q3YN+cFHzMsUw7zGiZBSOTqGi9ghNCkt5d
pXpNROZ1BLUKArekJR2PB7XkR4V3UH9ZCmRMJdEGWkpgvGrzlZv/u5C1rb4fe/skmjOhxKDSNaOj
0R84s5PbbGPsG8J7e1Wof+3Xh+761GE1eetfTpkEbSap9SO5v4bg/J6LXOogF4UmQjGnuA75rjoU
yxU/9KEHjQfyv+sZGBoQNzwZzaBzclHQ8IWd/104KDqPsvs9GsEBLoIa1Pa5ErK09vRBbmW1vJH8
ilqqDnJp8sIXKL3mkWRd2nYqfMi/uuysJQAnF3STgQybzbPDfwqiJnq/iCXVsVGwE3iI25e43UIu
28zSLkUNotu5iNaEF4XW9YK/6a1aPXomJznNrTyFPrmpa40WHsLBSTzyAPgUcyP4Czi5knQhVzWu
o2Ot/o0+kuVMaKfpUghgZlMzz/04HhPCGx4o/Aja84kcLNWs2zQy8/6a6hdvKVDD2PopnqEta3yr
2oaD3nn55wov+lyhlQ3BKUWBBqyIPqpsu8zaQ9IuFJiWMaW+QffbwHMtH8RMFo7OyqRvT1FZ2VUq
wJWlwRdzAjTP+DRfeEfKPYYA7rTKwZop1VRSU+Tx8lBwWOZqVtAVLk/dnXN+E0/BEhpoPvNyIsZl
9libtJ4y3nTqST7OtK2l1Dce3AmaOOb9ANxTncEgt+70SQJxburgKvlgmXbqgSjLaj8/DWCpxe3Z
vKmckBogbP8RGLYb1WMm22bCO2XK3/ghla2D6uMH4Muc7feXkVBZU5gxGidyogJ3etXmZgIwRJ1Y
32TgtbgIG+bLMLt2ONpoHSiuNPBbe/Fwnk7u5dUkZOIILQHaRRQYPNpoaJ9rpFJsMRlmb8IaScpE
LSf4C3f7D+hRzk0eLCA8OYmvhmmfmb5Jxc7C1f0dYxr146yaMJAiZLZ/qMVZkPoBPxmc/5nF7HMl
RtIJDRviwKVjzuqjnUWSDJ4zj+yLPoIsCxtiDdx+ZJkCb2RBokcYojrsputfKRuaxhr0BKPy2wdT
XiCpAy6NWC50kbTL1d0zbvUBrNtKpZvDMPUvgkopx6o6JZhmlAyPAFxUGJuXcBX9mLTSSG+Otk0p
v1f2SSx2c5kR+oZL2C8Qsc1Tfj6OQyrSl6Y8HMRioHuXE9eLgRTszSIA6eIWu0pOZi6J54mpuZz1
CmwQZu8eu8VtwOvpsYI+bMHuZ7ACjEUXtFVU2SeihBofYwb1bGf67xhem7VhhZprPR56FDu8H+z8
w38tSUmrN0vuw02G+fHgbL9EL+YK13UiijTYNpaWocQPy4S/7AxFpPaK8q2RBTTlkLuvVCo5n2pm
qzYcfLqEcY71vXqtA16CSOmU0XaenUdUOAulw8yotj5Dos3ADIXANlUZse8d9yXARXXaIzpDnsnp
LHGNe3bNKJwm4j5xu/+jbtGG/h2lO2DIVx+9uo4mkpDRduyvue8tjqn0QfuFjC5Nqlxg7hvNVPkH
9Tj56K4yqeIF5pt4Cnpb0BP7HiGkD+CilrhPOvtQz8ZrOouOOk91i1k1qDj9pCtj6Hw7Qx09rde4
vkIyvM6dZ3v6OC4b40o2llXoz4xsgFtO36mQKHQr+rtA7K4CGZRkAWc/858xeSCZJbth5kPvspvj
fbVr6JzIVGOCDXj9BNXXagliSj4k7fPNbPWRxb/KWfuIixYraBtrOSKssxEB0mXaqL9qq2zstfXA
iM89CWcR8h8y8IzbR80mBxYQ6hyClwpUocTbWeFhXQP4+LfvqtPHPpw/LC/WL9186wI2TC/KErVI
ocKupZ6TP9FjDUhaEw6YYKyy12waYgdX/H3EVpivXop/Aka9W/cFmDCV5GPmBV2O2s/FMrUwLRS2
OhBsKPdMCIIcGyWaxXSja/hP8iBqP1KDMc7uCIZl4plKtMV+Mrr/w7H572tXfk56OojHMkJ4MUhH
JxsG0dcYHYu4mPTJ33r3clvGoBKblzp4kghw6hVEzMbHwvBEVOGrgcWIa354beBydh8WWGBIALk3
YSB+kGfaUizuPC6hx0toj6AkK1ekckZxA/LEwQX4Nzx0DvpHwDdHC0gGrXuGPhwFzeTmxodRj6e0
79XHRUAKcfLCNJjnYY1BzoGpDS7oOzjrNpSh/yHnG7npiiZhEcEAtmqLRpLEYQDgifRQmBKJtbbI
j+Tq9L6WqzzLa2THp+vQ9OU97ZeE/acPBOFxgmiZk5f4DeZOCf0BJJWWnfPnpF6IChB6xC8OhKro
guNhATyMKsRBQF49wTDZ+UTbzLOWVBOaOhD+V1fnBAyfGP9PTZQjII4mlgkOpb0InQW6rS1kZFhm
rBeVHWp3e64Q1JeRKw9bHbARhj6qZDXU8jIHPUB0N2sSMY+trR9VcD35GoQcX6cr2nr6gdOM3gk1
0r1WmbXiCNolSUiub0yDh4rWEXXO0qLQyzw6EgPB9A1Lf36dZr6wOKc7FX/3jiItkCSnGibsNY5d
dUK0m5vWK4hcymPrRC49BtGuJg872JyovYeXkxvgHOsKbx3B6/pkYj8OaQf9usDYptOzGq0MbV32
wR2h2rgN3vz5JMzRhtyZ2323Y5MI75GDHbliY4aJV2SLRJPwJvwo4hQA52Ads+/BaC1Z7r4cl3LA
5PcsA7LuQRA17a2pAcuCllV6X26ryCpwPcyKf5+YNnzDewFVGVvKg0OvbeFMYJipYHf97xulE7xc
Y4XA1R06YXme6ptiYbZZD4YJBTLCagIyj5sMSZ5wBKY8aUAMyEGKdZtqmaXcJJX/gv8Nlpn9gN22
4VvVyz8XZKKbwCLoE21rBtvXL4PeP08PGpp6HNsnqtMMSjLvD9DCT8Kr6rFB2VSLfpMWnIT6W4Gx
7Nq/M6g1ceGZX+8xeL+IObuhxHIkyMHFDaALearIAV1d80r/GSeuOw7XxMpbWaoGsbOZ4eoNRqzZ
X/Jb6QudfVQDTDjyZBVLQnK5NtWeI0e/ChpgYuXzUVnQNaHzkn4zF+da0JaEGIz+Syv21TyMzUI0
1oTxK+8AbTyYoj5w8ookoklOE2uxtRhM0RydSki5YRpv6Vjf5nWNYLwOGdybiR39HbkLvCeugOes
K/E0dobiJRb+rDc5KNtGjJqu72nrXwat/TzuqY4oJ5oWULQfRwxWg7Vsc4423O9qU6eYY9l1zTEs
CmGGQgbGrm6Z5VoOUSnqPxMrS7D7RP5NlXfKdGt621gZCz3MhwiSK/nrW7voYHODZZLET3PPsnYd
W3Hf9060t/RrxzeMlbwBA0PtTA7o7Ld8h3Gd4i9Rbg28r+RhUkpzM4PWnMnFXy2v2sTlxR3M9JWl
DYDtaa7BYFBiY4XCd2x2duP5SFe/wngyn5nuXEM4gFXn/0weo/M9gCRwpjFS+4uYNtgFbS7uj9Yd
QpTd3IUtiwQYRlhhnN5X2Z6c/4t+N4yfWzR3jD4YkekBmUL+YjRIikGBYEZsZcUxdygF2SvDQRgR
Qbu7GmD5K1rFJTYI4HU7bUf50iUnC458MUGRKZaP1XIkulrepswpz3M3O0ny0vQ5DzviKq0djLxf
pP/SYA62g+VCVVng2ca7P6SIvIYtPmW66EjhzVvcyxrr8gRgi1Ra4ZKjoScLAfYZqDOv2ro8aG17
aozSLhDOuWOqJmyxfEVjLW85g5+ucFKSkAjf4JYm51c9vOsC0IWf5/k5Bb8XdSHN+bXG/+/irRD/
FEQ8dbitV2SB88MQA6ZYWXb59Y1X6fuoqomqTuYcGd5igM2vh//3zJNs5tffohcDY8KpKa2FKfNM
4XmWUxA1n1Q8fV3dOQyM2sE23aqYatWbIWOQPTEjgEW2M74htWaD0gAcIuiD+2Rsv1dohLKNnrxO
NceU1UmCvPjMTo3+2eDeBKuWwSM8B33yrneVacgRgZd/Z9/PmscqTbB+6Ff8/sGJxF85Q8kejHVU
MT4BQ0onpU0ZB/0KdQp5gKsAT5KyO42XXZPf2AYbG9S0SvDdsJjv0b0X/2Zt7ISmmSTPqnwOmVmv
IPxvtjryRnwO9l8eRo8tc0KwLAQdHulifr3ZaNSRnNOFfUNzlwKl8PoSMpkVsDIGNP5aQT8ShYEB
mG2BGMOblRC8r1bCmzuLyuadUWMI4v0gcwqYXoxwPXogZvBxlObOO0sAMvyML0IYm7sfqXQHEmmI
sv5J74SwP3NGLKXDxneIEFiRZppmiS3ZJ03QWkxYNN41I02I6sPpWIetU5CUViFiU1y5cPyIQygS
SjvtXrFs9kNMPlEghkYP2FaDVEJQjgJJyrt7y72iVD4gl8Vt0+aVKemRZ4fcTvjXqoZYvY+77fYn
aSjTdZ+wOsUskEheFKYz7ooy8lh5TX9Y65P5x5kVK6Acmg71EhcaDvMCgMrcBQmqcvKew49g2OIu
HX03InZ+B6/nQpNcFKE16uYj9hyuqcaFZAZoWfX5OIkCn1ICMVjX9UQE9r6Ly7Xp917R8qACNw8D
63rGQwj4tMfIrRYWQxBUsBG9bYqPyV3QYfRW16n5WeVitjjqdT1qKpe9yd4aOzGqfJvMYqUnGXrc
9g45t2KrR0ZbgdIGYaUNHtEsoab5Q+gedzxyNKOAVjmjFjmTCWwwGDVmihVB8HBgkyLMDnkptjjL
xlsZKtBHdtsh4IgGN1ipyr86mr7rAsl2I07Fin1ADeki/D1b+XoDNk+mQhHe1xFfI2CoEjh1MEME
m60kQftSA56tlx7u5yzeitVrGh4Y+NQEmb+W8YbeglDTrkXIGnEI+eoal7oH1wjKDEESXMepxFgg
VLCpOOoBGm+3Vrc7FQCmd5LOTYWPhryT1rrZikiqLLmvwjuX/8sSodqfseJE5s2MXAOB2EFEhLGE
1mJwbakjZjFW6qOeHU5GVIoD0DtHqZ8W0D5DAuaNr9/5KqtvMMXI1mg/2Z2YO0IK0mBQZ4Vvlmc6
3Fwdd93H11rLojLWrUiY+gpUnuokN7Xay9SjLhDryQaVAXbb085lNA/mQo3t7vORJ3N369xkSfJ/
teMO4Zc5AHCjMkQ+qSw3dvuWonUd44tZpvu9w9okLCVXtuLyfcmYMnG5+iEibLBnDO2Jg8Xe6kQg
ggkTMdoV3IC1eozQ6ac0/kONpVJeOFl4xjNX6pRiyjG3nFCtcBB6ZuFfBfvNx+7EZFIGJm02xn2q
L2rtCyhQtEk+WjUc8Z2YGtWbLDT6UPKVMFosQQ9m3LjaiGWEsYAbxRUUUhbHligrdsZt/tl3A87R
FtY7AMqE/JEubaAdtC0dSbQZFiAlnsA2kUIBjOBCsUeNhNeAvMk9/Lf9Lnu5ZSGZBjbdvvf22NT2
/XYh14oc1OoeDQamSbxTLnDeHLXcsivOi+WJ9EiaQoppSV8l6d9A9Pa/BQH5XZI0XQATsfY3ZU3x
8IuBjGshxfiXs3ropzE8NCCQw6Vm4fTe8Ixd9OPIXunn+2VXv9zAsQv1pQxI29OueY1xCazokLC5
pQ5jeYA5XDGXovHDRJ2qciuAX9aVbRof8+aK3aYmtJCKZsXLImwMG+rG5tyhx81/kDDCIjESv2bw
kByO1wmjbgJUWxx3ZuZVYZStfgvkvNaWCj2fkwBj/6YDaamzxjRLcKmnBSALpHQbgx6C4LVmeTs2
OOVjVzQ6kh8Ud3BlASLfV0icLCNVQ6aUwRyPLm9+7SoLSg09I97Z45H0ert1C8ZiYGd4Yz1iaH/I
slBn1j0ODuPW0lZH3AsraEJ4uC0U1TiNkLyR5Pxrrf6nemWaRLXnONsERLWMFoQYlQXSW7GYBojX
vKEzTQ+0aCLHuXRJ9ZUMe+VTHmcizHmeBEwS/5aAf5PzoeQf/bsdh+di3KiEBR/Vlo7u5jdph8/N
B6Y/l1BFvEJpZZl5P2VclxCoU/ThZVbdn78uqghdHHybqNYW4n+RLGGWYD5b15/gBI9SJSsZbC40
xjV35auVKdarq0ZDi6Ury/9SAjeWU/MKs8q3+HUIzF86boz0PB8vVz+5EWrCfTPtU5nMHMuTBRnt
Jl2xeqGLvPEtMlS9CuL46gNdf+hAEBmNVUGnbE0Gzv5KiImJHktRAM9Av/kM8p16oQo1ey3QgWg9
WOO2B+u6thTn0f1ucObVdQkFCSYGi4BO51/QChzs18ZDj5tLDYUMN2HgLFz/de9OnkIPgPiL7+lz
hgVgXJNpIO0L/4v1+XOCc/PhKOLnPav97BAyh/RI+CpwcjKDVWURUjFKXCEFddejruQWga9LS7Pf
gDjtdU4dHgvn8dUW9uWzv+fr9z1sRA2WgoyAimHRQ4Tn9eGZuq1p/wCx+H/NN64XT4mShMi2Mwlx
+2I6Y87DsWe9t2AoBNMV/nawixOh92sGWXbKs9U5l1AHUtOKq1+ABQDJxul5X2HS5+0yVVaaoGd5
5cEVRZiYE1PLEfhgKFjrXMQ2SJ3+a9Vbu46SiM8I0IYKgTEXa6WqGoVXwUIFJulRosZNqE6qK/m6
Lqn9RTivrc92NCoNzsTjqLcDPSAD2604GIA53eBonf+UOl1MhZa+1rEKvlQqtOvPZXSOroVxC8Uq
Xifd7b4Gjan56roy+9mDThUDgO2a2SN6ZkCIAceD3OSEGT/0RZkpBdQCs+LT/RTzsX6PgclffAVy
XvGewikYkQoDl+Z/+0MQcdFhLUGHF8ptz1A6xgRefUmNJA9RRZcGM+SGNO8gZ6Cc1/mcLqVU2GSX
fvXaSo07+bnjOaPBgzWlBXvBXE2+9VVRJeJWX2n8k4E0/QoHDLZsYhtSHp7Hs8LO+2NSWLjAjM/R
NUm35zWrFGYLzj+8ZPiends2Dgr7703RQ1V2dUBUW3nENljcVTVBOCGD+rt5C4g8jkcf7rHgO3HX
YuVLWColU64S00K+ejc9sVcqa+D6wdJ2LA3LonJM+O3sdBASVk0PYORItMOBJZtL420AE9HIKeDT
CZ63njmQY1hTVrjifRcbNyhGv/476/57FahMrVeslMHH+nutdjauGEXbThj7XLI6grGDvYlPDWgc
VqAng+sImv2fXUsnzeozbBMr6VWIQvh5rUJ79o7wC33BNkww1W2LbD10FfYlMfeZAEx6r71GzOKw
UlqE0XKze5RUiRBw7Kv3VYkZglixhp8RBFluwHd07DbTlKNrcOjgaRunWOGesmgBQvFn5qYy3U6G
vaXBGjpIpaTNgL/0BhsOSfiTXZy5PvDtxTPufnYBlHd+5VX0Hym49N+Gc4ZgaFhotAYsdiwDwR78
MKqAPhnc7puRRbdsw4bIeTOBoVtrk9/PANV2ERq0oKB5t1H6eZRfl7PIqdQkMJPBhkFZFmElbjI4
satjiiATckdc7uvTiQZsjeNzGEOwvZN0Y6jJ+S1uMBZnNDHjilAcJe/br59fT5hA0foxjAbQ/IbV
9B7HIAA5aO6rLVWpHRs2aNtkElV8PCbi/0+KWa489kniq39wBi1JaASzNKsFy/fsBFnL9iQHCPow
NPGqMIl5wyEZexEggEJZsV6mDJStQxzkwDsBM+ZrcvBuKKkChgOakn8mFEbQ13OjrjrfgNsEmflW
qyhVXpl5pAMw09hRfOh3f8N+lWoxKJrFzmxQGCnFre3lDnq/Zz4nsnv9GQfWCfuSPbxfRJObnzAU
4CpGLIrWNvFSnNoED8D5UDDCrAMuSBXFtW9W1IU+/Da22MG7xGpJ8bT78zIcjDf8i7EPzmEAQu0C
yuqSDr45GB2XqOyg/oZ+kKEGl2Vj8Ga47i9UDcsZHllV08Urz8z2dYS6zLaipf2hHHZxdWBGYt5n
7FgFYFUxmNWyVw91m4sUQLlkHRfuTD65Dv0DZyxzW38Vs1dgbcRFx0m0ILaql1zxlbFk83VpWjkQ
Sr9ql4Mf8otN0PQJNSkVaoeOIF+iP6Z7vTajym9dnFE1gpmyisuwqeYEEFA5KtADDgDUTqO6NqKJ
eVYAixnDOlRGlp0Q52QBoPMciB+WB6ONL/v+Zf7U+2HJVgEMwKFcZIaqYG0CJhwHwGR7igA43VQY
wmgn7qFydQ6kzHQSjmTR7VPv7HYL8dLvgYk8NS2Zri4cEcWQXZtbNjNWvQyEZ125zSeYS/+tDo0r
yEyT5oAatmxiTxRVqFHo/UouTFfGbBUOIBQubd+H8eI6JECZ5yzK5LGFVaSsX/PZe2v+tDBDDRuh
1WJCFod8C6G+9XTuJojjRjNsC/bWKtGq7JJk8KGwu8p74ZnTgdgwhbWEp9GVlgOIPGOttxCyR5EF
K2wj9JAP6a/P3viM9kjvjZUMIO4l0r63yVo/GPWWYYbXeeZgtG6i6F2a9qwphzTuepQJAmRL4gBS
NYZDiOYXtSUfzcqK+c1o/pxeeH9/X/BhShaQaaQmbNnBddFJbcC9ZD4FVbSoV/mJNBoZ8hbd3rhQ
ogBF6ueV2ntyId/2aQZjyKDhYyWvt0WcFqs2cTasCE54N7ey9iA0oKbHdfB/Un7RSVm2A8+2jVdx
DiApEgzMayRjU8kLm6VCHjtOyWnGvy4wPI2CD6RedPwtCtAvIeHHMbdmuQd3xloAQDkijTASKm8O
ZIMwTQN2Fw/uS2pzh8GK/LxkHRLwEsd/z2PoXj8JHNGIz2Eiz002R9GbtRtU+BP/SSphQhZiT/VO
h4ZmlZ8M3Mzo7ADTRv8GsPQlOEmbSm5LorWYmQIOiBFVIDZdOLNNrQvYZSt7c9TzNzgiDhBk1KwW
uHcctGhUdIx3+RTEvrFUcuYSmYfnbP+NF6QHLfpg+wrWuWCRihHENHRRX6kGLi22fGQPJ6U/zXes
3WZvKu2gG0MAZ9bD5tqU62Nxnyl7Wkr6wi1tYYfZFzfvs3DTkDbJIAoOPQKY2s/fHhVailSGsldp
XEdp4Fj1/sngM5FHdgzRXosZsPPDBnxGt+EaY1XctMPzOO93S9OtTbVd+EfrEK7tpyatSusiRXhG
+RatZ7sTcVVRvvrlxRbSZa/LuwOv6L9I7utJm2ZBFC+U6ey5mOwFaJG0jW/MVoVmqHEmWt4fSx6E
uQTbKXgEqegunlYdpov5tdsGQadq3ZxWyvi+TIkUU1CN2KdVf7BalRyEkwopIfGdBCXn2xZNQgsz
3OYzYiv8/7fIdK7ukHVFJ0q5nWiVEs7cHonjGdMWwvXpqaT3w5LQLFjKt0fw21fY7Qw+JzXhIRLV
C+1Oms+LAn4vcecHpamhTTkwmwpkREKBqAjRjRwC7JaLHhVfEmOiMI3ZJO8O3ZnwmP/b0bAHtabR
mLP8NAz06tOSGZQiJ/ShOTfXxxWpcD9ts/vszILRXvZbAbE5nw8M75OCjBMvkxq1nzBlB5eMaC4+
uOQMvVyDzfRmy1SAbWAVZEVptdq3JdAXtg66zaGqHiqbhOpONxpMsjqR+XERTBnwPVkEkiaVeA8N
I+f3YxnqSzCXDyMbGKDhyCZHhSoKwxx5xFp/ToV7zFCLIRaEqVbEU9WB5p/cKQKpkOD2Wty7cSlM
b4+rlR/40/kAJaskQEiOQ3wZqqTbYUmgvm2KXEzS6mKmWZKmTVPrvlFxtCQhOFgPhgFc6TYFovsi
rbMDGB/QL8KVs8JNTuKakzrhEpZ7mNmQsTHlbKzLiYPa/+YcuTR1HDuQkdjhopRl9OowpxF7qo/z
6yKiOPYeMIrIQxUM5L+GrnnTWJIdpsoXF3aYVlBMEcOHV75+GlGAK6PZnyZAJulWXPlzL/2wmsgU
Xa6mHFW9/ObpXdp9akpRwSQsa25Z1Hx07wel6Ew7byjVzFJ0VCL1jzt2Oe6PykRi8suQ2HvrZWpV
LtXor3l8Pq6jdLBA0bz15AjRngR/v0lJtt2L8hCY48b4kdJTg/wHR6S3/OwZXEAvh97k/dPdNMU+
LPqsLfuT0oMSBSWkzJOFH0xVKN2Oaz82sjg2zonuhRO6jxJfwn8+ib4KVqISasQKWNpf7NGNxFuY
AzmnxEDaBeHQBwS7QPkNWn8pxHjBNKUSJeyOyzikYyVkT07X04hbNtkbtKV5ACbaShvSFk2RSbx9
Y58ttoYc1+MqZoGGaqTG29H8Qwju+uRfU3NXgeY+/Ues1ofCv+PmFnRp975CoAfO7UKdu2TTxDR9
O6ko6x/bkZ3N1rgvMxXO1Rqu2SeS99XluuR99eemzuPXF2Ll+S0NeB5vW2798d+DYqHxFN2TAka0
6Xr9CUUqufL2/gWGQDzivHok02HLL7c2eUUMO7yxd5XqEIYdacNqn7g0R8MyH3u9Phcpl2o0AeMA
3aXbsyVAvFraPNDoYcbI6pcYOwSWx4JDmXYgT3OYWPmrosJl0dk2HLSul+aB7+HrLm6EQLau2/gc
tyzc1awds3Wfq55cI4fqcjMnwFrsq+YzcPRMa4j653St5ukuqRUu9aG3vPZvat3EtthiTVJCTGsS
uY3WMIh2XYSkzdHUE4rFItWRnm9YK5gDLvzNcnC82DwXt2cyWSp4bjU/h5Q2nvSRryUD6Ks2a4Kb
oaNgEylJnmBcKIPBM31RpWECSfZ3KTPUuQyPNiDdFFQVqVC/CPmdWN0E+L28NUkpjPTRkDzPtww3
Ti9G1vsWZQGKEyYoqac2K9f4PiyBNos0mzSsKzJJkiq/B8mstx0oKVUMhmQXLYS/eLxsniQz5naE
IIB/E1P4id/SZ0hm3A6QB5cTkSgH9Fs733vYm9KOvDj1uo4o+mDWPNyOR/h4E+qJXzoSSsOn4jb/
uhTp+65ptTmOVDf2OoBMmV1TXlTjzJJC+Udbu086tGU2EqoYCE4bS57aQ16Rqzn9QC0jnrzSh/Eg
DWTVgI/bNjO/Z8WH0GLBpQHs0gc0/i9heSVWDjPGTVWJewV5jqa6oDmglfeOq2AEgaPsSZMIQ0MS
B9ThrNcUyvjmm6T0l+pQgGcJ/ozxl2JPHTUn7NwYhGOfwwgYHGfVU8crAbq7N9WYeiPNejaQ5wC/
xrGwJATJl0b1MiR5Qx100Z86BePTjtLirSO32GtkxBgIWqCrjg3BTTn4dbmUfdB/i4eipYCT59ER
oyiCaW8bM5BsqPLrEhDvk3IDOvGp7vIFC5Ptog5LdafQf/1Y8nUjv9CHQQEAqx8lp+lKbdKHHwTr
18UN2QIapCNrmRUFmBrMW/RMADwI9dAB33s2LKrRtflquukWn+dLd5COEXh2mahkExactXYWby/s
1Qt9yVLsqFkxiNp3//Ci6C4tis1Y4QJASh4G68FFjGktO32tqBkA6cQfmJrNc43FqI7Efi6XDyLj
3ZjGRuFxxIbA/oXKrDqqHC5nG9Ozr8d69xF2z/3lBkwOgAYGPKN9FlKEy4nSNWCdN6uv5pQnGH28
WQg7xoWLX77zg/6hO4Qw+5kqu5KBe4M7cf3duJxnChnsXS6+afsup6RtF2HL360dlt2LenaTfc6S
mohcN4BMaKzvHKXwSuiz2kwDkMi3Ny0BO4+HlAiarKFJb+xnqqCmVNBakmFgSAEmlpdCHMjsxFwh
YxzIFaeBf7S6UhQwA4T+f2As9Tlo5tR7SSYQQaUkuMEdWD9H4XZvEyPtWeHo/C2dbkcKKY6YP0o0
lFK6fcvMWaww1rIEPfh4OL6fFZp0bFvYwBBKPbXboCH6iVhxm4WCpq7tesnzv7ml2LWmu6XSl96/
DxC9ZAp6AtOK1dB+MO69MTldvxpU6bog6M78ojsHW/1L/0C+Vugaf7DJ2ClrmZe4CBOCMq4Pa/h9
A8lSR7IIlBdrtBjOqnoBpe7Uo3K+jvvadCP5c8kr/cby2MW6C7It+QO+JAfw0ZP3b8ZBjLNzfUHN
Z11jkYq8WafCIXZlCHuK56MCcYzFs+k/a9yxfJVN9bQ/l1adDwULQ7Czrm/xpMivFZGB1PV2Pl9q
ez1Nzwot8Nw/ebVyzWN/cmncdmYmnh5Raep8jWdA1+O6Uh45ehss2VSWb4QbTOY9bYDTRFshMQY1
PaKKZBnil5mKwcoTlyhWi7ffFiD3NHjqSYsEtavMaI6DHd0PeI/NWvTI0ywlGTuw3bt9QjEG7Pjd
tVExfd2xMFVUW9rkPsfAKTnAZ91INtA1tR4LF3f9KVjmcO6CubGniq1FYe0LE+zbsCugJi/iUjI8
CI12HVRf8KbYxL/YloTkn8w7F2ng+/iN49axr6zWWViaEP8U6A5qqNNPc1dq167Gnc8bAGOmSDSw
rBzmUE7X1TXx5Fg5s6KzlVaVXkR4hxhxmmC+iWL713EumQF9gimAE73ZUXo5MPWe8yYfMXytuFYV
aGEzovRsv8Gtpt8t5awJVsjak9V9cpFa1xrrGbKKnLtV8HfB8aXw+d/u5M63eEelNlfGovWmjOjW
O7iV1V0H4lx6VUhJE6nOvYpW0ZIefrE+Oy9IKRb//KWQgZ7PAg3R3Z1rN0gCoqSjfMoJkNy9CnhH
tFyQ7CBgXFoQ03cofGmt2ADqHYF1IktBABdzWh/wECqEeeq2jh2Telv240Q1Cx0g+rQPldHaoBC0
rLaF7/lr4sqWpvAIE/nPTCsIyzFynomHisXPLRnawAXLUxGN73kq50HydOK0Wo6VY853r45X1vCg
MA64jCnbUpMIgxPmdchb2iSRBKVgkem6+SmGCaGh5GPd0c1hiMB+zCN03j1wWDQJYTwjLQZiJaEO
3k49yv2pn/j47MtivUD2rB2dU915ftU2f9GOq2qOzeV9oGBeSZM9uW6Q+lCnbQH6SHd4sW3wCROg
oT9ed2VDesryhJR6Z5BcuPE1w1+KGTpKqKo5rL69y9jMRCM1XbYnPm1oTradyh6KIyyC+A6kFHcn
JiBdJO0blVb2T1Mi64/s0lPx+PRxgsrab+it51ugD6xIrDHjbGi6Xb7Dm929fBNAtL2ovKAabDXM
BGYR+VDsh42+nMZcaiGk8shtFEcEFKcyrT/0RoErhpPCMwaiiZQy1YVS1QuDgXsMTNWEn2vkuOMn
Vf2wW574xxL0DOM2r6Kmlm7eCtyR6u1JwqC/EB8Y0yqA91lMJ+aco33LgH2lqbJij6f1dhZufqlY
lnlY5xvrPRcYGC7Fe7wzFquNoEHSQaeElZj5rj/PbKUATg5oXg/ORGCPK2hNY7TiXR6eagLMd9mx
yfrL+UthooMCx/nf5BvaV+1fhSqzfXZJZquOikFZlDSFxNXQk7/0DEdkwR35I6LWKUHEOdNEwWj+
PM/DPTk/8jxxXuiehj400lMl04COjOAEPLWmYL7AX7ek0hltCmpnFwJQ1fzvWcj2eukuRDXk+Z8M
lCW69PGRst7LtdMwjM5Ut4orbOSvNuG7D6AcrvO9U3UV0fK/K11ERv1LKFI6NbHEHdNJn1/AL9A0
kMACEst+vPiWnW0RseqmwK4G7BU2PaNUM13bZIXr3srZWFRnBvCJL2bhcw2wx9clM5d7Hs6iSQi7
H7Lqdpa19qZA95ukt0ckbRFOXC/H2ZtK6PeNH8tUTdS2tdViDgPdlAx2Fq36d6iX1Nf4pr6jgRn1
RJuCoPt3PGUf/9I4mVOWQX8cwynJi3CwMIjbPRu8ico0jJ283KETtPTwVnujY3j4Rqmw3tNQM5MI
FlDcVeknXa5H8ANBGHSwyfROAESxzctUF3bENpxPUh2yaz7EA9yrrdikLR2T+Fpqm7bX1f0H/cti
yhSUjDWPYNvqEEI/AehuKXAvYGtwvpC15/RXKWo4rxtpfNRwnExkp7rsdMaqgZKpp8YgIL3RImNH
dmwHOEOFtZmeGn7+EgXa1MKIV7lzqx6q75HhkCIP2IX96MJEMqqhQXyTxdRMcoLpcbQge31z6dko
1FM4R4uon8YjFjgF000bP4Zka6ApHwM/DjHmOAWWjfB2bAq9PjEnUFdk/s9jf+rgx/RtVw5lZ/9X
upSLCGeczaRWYEYdinEh0uTlFaYjJSDlPDq5rN+Oab1D5POueTc+51FkB9sKavqA7sxevmOAzAfh
Iyn7fk6/dw7WaNCE9dhkesZDuZIA5AZPraDH6mEc1t0F+v0AudcYKkejf+crZCM6ig99OVXc6C4s
YYyF6EZ+ioovUMxW5tin66OnSBhRKP1u9VJpSEKXaGKL6n4zXJDRg67EuzxD6zZVj7cToZTdEJcQ
s+nMQ68xZpQIRLh5CIEJWz5Vr5Ya4yU1Ro7YTyyyswvjRR/0cqbzeu2RCuYAxxmBGcbN96Q1rEhd
+DGlzZoYRz7goADfcbbYRBPFLxndwRb/shMkPyPh2YA/jEcQkTmbqWUUB8c3CVijjKtk+O2Pzlja
Fb0NzxiS1AwaM3zaLg+JUNurqq+Ee8LSWSxe2VZOteKhETg2QQ01jQs/8JA4VSt3Jjsb/PdrHsJl
i6svKC2/Tc6f3eAb40wHkfEAg4zKz9gS5VjTr7PHQZwtxM6JGwbRLsIQCitRC8WbPLL1GHIdgQB8
fuOsfNYam3a2VlnEreZK4bT6KvjxpfNAyTLeVUUiWxwsw96MCReNiZY0goLb+H+8R3x15YdMIJGf
52SDHQYa4sNTH2SurDZO1pocv+hvCTDsa4/cuzcQ5o09rgjgLyObLpPjTON93/fXZkkrvX5/W1MB
ygDS3lIB7ZcxiTz3xzc7rJLfM+T7nroKtnt0lghVe1xPZnE/8l1auR/UfNv4mnT1BFfGgBIj4/91
FeaZGGVwKLfDlGtKcYPC+m304+swTDiItaV7mMLcq7vjtGl7Azx24kRDeMwU1FmnqIxnNI8RqRvi
T+WjGW35M0FACxuY8wK/ApBXYYGA58OTiMdxbxtXxlLqqQUxO/4H5wjq6laFWK6j4HnIz0AHQm1A
trMgyIjBLX99BDsy5ait/YA0ClV3sJZS5ZdmwjW4K/45WfGFphTpau3YfOuKxBot0bgw6Rsmrf3Z
sEgFzJ7ioSyFQVv+67SedlWjDWwMIvqo4ofTWsticCscZtFYux1wRWGCmcSF9pPc5ysvNLbVasGP
xLu6pWNrpYWqTruO8G2ZxXJD8xOSkjomYXP6P2DQ7iWkHVf81k/EY9x56xVVwBde41rb6y8K3SGS
VA7VtzGZu2J9Bvx5yJg2RRUhCCP8wb6sJ1Kwe0oWIZGkXh0fSq1tOM0M5IfQoJi16zakscc15DRN
Wy1cXZtoba5T7vbtJNBm/0eZ8WSqkYG7FnRaDN2BjKDwNMpulHwRBiB/FmQulhf3MRvl7JXcTMso
BtAscE1JLiMlsNyij8Wh/sEKYAI2N/6otRkCjtWT0Q2WHDgHVf14aBDn8N8EKpa77tRYnabK8L2T
+/bNP0R2+E3FEwk+fRR6rnhN8rbrk+h4GcwW2v8hRf4G0g9f2da/jqwXjxBaoqdUVImuFD9cCbJj
SeMaLon4WuOt1cBzcbh/9v1B/FJcIgBMfh0PDJjcKhfHw/IME4NpRMETtu2+r3F+RijSw/9SVEqI
hMe2qyLv8AuspR+8BpQPob1W8lMDB3MfuJucqcycfu5hz6N6ysz1ykbVkMd2fkC6rZK7rGgiqREo
K+UvXZ2nXz4caCD+oxW/h5csZEfebZ6bzfZHAOJaWPIS/QIhN9G/xx+TrNfFxTURqkm3bChLmmFJ
WxiN+WO2iXlu7woxBtT4uSMxc/7czQu5RgsfPS8bt9PYKeCAeJeG2F5Pejz5MBdSIb34EyEVTdyy
ZoxG+p6Mi5x2p4eMvgNyQhkr1HqJ9BJWhTzn2DBTSE9nmj5w1iyNJTB+4pXkM4bMKx2xBSAuREv2
vXjBpnEkzQT5++lrfSmluVagE2lulxCi5iBeUbCcu8vZSf6cUlIQXP8u+2afaCRHhM+iLmuLpIx+
lHsweDc3a+pT7jEFb5/bV5Hqdt95Mtwqxxf5bK16XsM7DGvkztcB77ABTo+Ly5oN9WOjv0IoRDGg
QpTBhWl3CYAvWm4Rd0K/JIfGGwPDkSzQHVa0eQEiXBJ7vOZNfr9FKUKFlY1u5eIVyj+iBKnX2/Qx
Kp4DYBsSi7AQiEhbQELXIeAPRRD7bZz0nAZQ4iZwsf8XJalUyVi5K4a8OAMUvvxRvps0Hp6bn4jD
QXEQqTG0sKJiBgemt/RHs3DdWnmvkexLrmDb5TCC3/298lRdoCvNmw26CQMLNqtod4giQ7R2APmQ
VIZS5SZMFm9ERjDhCqYylwo6AtYPKc0DztJybFywx4Q64iO3mabvIRRtcz9OlLPWvEnQoFwXaewt
vPqnUHqPtijUqaTTg6WufIX57cd3ikhXdU0UKCk11ws3pfbRPSkUoHyIrJeIJzDsw9GX4SIwGbdp
ewrRFRDloqR2PJxsC4yYrSN0peIKeabKx4nMQum2G+Ks/JpbJKXcXh64ZCCAIjYmL8QNh9c13+XH
ElWS1b7QEGoUCJGKBlT5IoCawrDUcn5WISLoTv7+G3yozKyZNVLt5tBsBBgkBgPWTvBuVfnQLCLO
iLuSeTStAMPmmHMtagzstSfBiu/VOilvriscRLtP6hw2l9TZCnF7XTzbkJZT6kZXdvJHlYFMHE9U
9jt5BvuID32EC4GzxCr6e2VYrGqf1H9/De8vRDzBTe7HJskKINodlxkv7X0AfPlRyRI4T+78IOkI
xoFmYaGT+YJjlKSeH2pRdVRBD5jKzYgHUpYFKOLjGgc0crHCHkGMVJ6mQ5mk/SXsJeHNg2idZbk1
Yf65jF0gKfzC7NFSUFPzyb0pmrjzXyOVAhlR9Etjr4o/j1cTnrnuabNf5NOYkmo6HIZwuk1eKBTp
k16h/0gf3y0+tCgqQDmpZ4SVt/nm1evbusgWmwDRJPDo2u3eBlmmpze2FaUe92Fexly8U8pC8Ktd
qpNKOuPdQvEZ+IKsMgdYoE+pVdO7b4Qu3PU59JiefukWxnx7ZKVQmXsp7eM2yBUC7PK8j+8ic6qo
od+Y5WGJWadRFxFXkbCBoZoncUOu3CZ8YnwYn5kwLFjfzb/Pm7yZuXe7PC0PHt2InZIhooQWMApC
S+YdzdtdxklEtLZPM53Op1fiU6aWMG7wBJLiJjWsDQEIarg5TlL63PiLbwrAV+l/1j9kWvedjcfq
+1EWxbk4qzMFAtEQIJ6aztkZqazSnEn+JFJ8y32hDILjMxWokUhBZZNcOAK58gbm89PWT9uvX42B
S4HDforLvYJrddsmiMbGR6XGRgo0LOF6IFnd75XBGh1pgkVLkZ/9BExLzQZnWXcI1kfNGqgxDTbS
FAQFg83Loe8Hq4x4oKqYJefaRzrfecjNRuKHLhr39G7JzptsldGDxPXh2IV9o9Tnj02uEY1EaTvE
pxOpHkGqyKmFFOSm1plUmtfWLbA9bSqfbp9HUg8Sad+EQIXLnc/J7wqEGyYw3ZK/MVM0Jw2qs5ZR
iUqnKIQQ/MNAoZnoFXgH5VTG6cymn/ZJdy5V8rxr6KPHQSJUxrMC6Jl39PmM/17JzxXjdLHyHdAD
fPxXJIa3zSTg7Gac/Hct4ihKXoe6rXAo3KDKbze94R3Rxf4H4iZpMzYDDY4GBJmgiOdVjnu+pjBN
AIVUK6IdXHqLwN13MhwvvhZ3tUvT/co/hlUHTX6sTnrQhYtn8UWQELQZZYA/Wbt/hikbi4mbplLb
mmfwbwxSOSirCYGMXFiaceaGjhotRn2sJ/uyT6/B+pn2MAO7c/tThivxoFmyIAvzkdzKrvb82Q8F
B1hekLzmujYNKiBR4mewWBhCBDdQAe2j27NG0ZKD9mUk2CaULwaFjskQ2/JKjmQ4LF6IV3FjQt5g
GOVDbuw8ACj0TYt2KZ6m4DG2Xk7/IClVyipMXnH0K6gim9AlUpIKIlHfvEi+K3SANUiHSE0T8jJd
5KuTCmeINZ527gpEApEwKYslK48ax76Qo2DITZeR7P7YpCM0b8fcjLlgxaTghczydCv5gaCT0FOs
vfnwxyiyIZGl3X5sGE5RYnkxDA2Js1TL6hANOXW+ptom/Ew6JpF17MBztFivo5L7DzZ8BUt1FQCF
mJmSKS0O+V1/yK0Z9qolH0Bkd+jmbXvXSAw3qeff7pt1Xf5NQ/14q7lPHDf/+hFBksCVE9DkbKrK
EGn1GoMOJ1I8zkxVfe5IqYwPjcjj3XbtRusXWu1T/qTZMKHUWuXBFLtzjZxKwiObt736ieJ+z7xg
zodFIroKGiPn5H2aGk+U3bRvPX13h0r8hG+0+3Xhli9S5JOe/8URjWmuCA/nhUpVg2Z0NNzsPIRf
fsGCFpbKzDo7OEpwR59RDrSUogW2OVQSFe+2tisobF/vbWPS51oo2vly4BNTK2CrXeEbIGeGxC5x
4E5xnPgW39Z3xUlXXPf/sHS6lTAsNIZm1vROjLNKzlE27qrP4SBz7KEDYeCcP0MqUhSSrAHiaFMz
gtz9VN1+5Boel1LpV5JNfcNCrULVSE4cV/vjPWWO0er894nL95Fzm/T6UtczDdwjE9yaoTKVwxhF
C5u0IO5EA6CynztDOUV542i8QHeDWrsD0ZDHtkWtg626cuWtSBqIKzqqmuZOcT1IcDhZKRmvj1EJ
aK7loWdCCWIwqSi1axqe55QGwwkarjrVSQo7YAuYFuVDYr2wdvq0syrQZxZQtYgHE8Jg8KaQrkkS
23IJ1b4rIZQcbYMfwFmSg5oBkPboh2aXsvep5Xs7CHOuTd6FTvXld4H2DqempvPJKKXOZ6NYVRj0
1KSqdrC3zbuQeotmPnJpnTRaKt1TpLe5J6vpSlj2p90Hcd+wBmd00Z5HWVcXsipJvYUGV6BmKTum
dWLn5SLqv0LI86rgvgd55PDTuTVgdNC2tKkJqynGY28mZm4pwgVuzOIbivTBOkpF9tAQovindf1q
gaXilUBp7gPSSLPr9nWd3AmySVkpjQvxhh7PnCNLJJ5MTE5i/dxxMyCl+Ef7efDdaSv/czjxLED4
1HGokjiyZawUFa5tat/y5GZO6TPVMch35A2PMNQI0giVFGfAnCYWU5ZZRS8ffsum4o8kTrPrcfCe
SgVgx1Ou6VkpnjPU4sPJ4sWU/4azvQ+cEGdWmpY5PJg113yWF/D5GR0WASLVZu6JPu8OekNbxu61
iaHFDRzP29NwSl9nAGgTPllnZUO/FNI7j58DknIoQFhWiV9oQGFUCL5XsDONPUo7OM+mNxWZ/MRJ
UZb920ux9YZkgxa4WtGvZrimxspvw2Px3BodOrPrWBSrMftT1PRJsymSZOSdas7AEHy4fMgAHTo+
MppkmDqzUVktuf5/r+h2DXhNtwFDNA2AnmjyC7W0XSM/jog2TLyVSTF4PCFdDqTpDJzErlzrQi8l
YVu9mqWWbaI4affnMPg0EwUlPVrTCMTde+qOJzcoMiE1zmc/G02LulJN+dB7dZy88KgeghIqsHxt
Kpv0IkEI4fX0kEbjJ0caIN5CEv3Scj7aapzyWQEaBg/bLgdinYuxBg8fqerQ3Je07/951bGTr8Dh
dd6BZ7VTx4Io6Pyv7MumneWXHEDNGLtUtf3GwvbUam3Hayadfr96jvssqaGU6OMUGGllSvpPq16s
MQOhnSxIfcuUbSC/rA7xrD0eqJt+P+ZxHH6JbT6IhhaMyLkKM5fyCK7ohuu/gykg0de8LU8B0t4V
ytHG57zjZD8H8aVuOvzLeNelbaVIF6kgcDawZlumBzAhEtQWrPwbfxjmI/h1zBHdLCkbXtZBexMW
gbMN5PBbLUH5t0a39XZhhQYL8oFQfqoV4o4NbDOnVd45FHlfW0kO9ZJnPhaupGqbx7sCSQu3xSNt
W4OOopzIHQC+o7ST3RmeyWgUeOcwyOOgNf4g8fXSqRr2uWGZf16Ir8MQWSNN32WPeB2BUup+gJZr
FHBAn6HhHv3vqMhfV5pLsNbmXyY+v6iMuZX0I3WL4HflNL/0KcsNqY6oYQzPX3qpRogyLX3ad64T
Jb/0rcZLpDZe+elbr2qKVCKjP9w3tl+85RNk7dJLCZyWq2Uzn/T/jyQeLNiDL0DZ/mqfVxTyK5A2
B7Xzs8G/25uJtFNoChjMGYHbkNGC8k0TCHXGzL4nCYb0gJ6POzWonfRO5ZcFiNuqS5kRF5Q57GNs
eoMB9LXWgWdxpn74mhux186KKuSExU6RloOk41Mgm+Zt4O1lvhdrI6W62awSpe7dsCk1rY46QNbm
zNSvtebCvC85R+U5edPuGyM98UOYZV6HTttSTwbC7LOs/9mfAmJ+vGQrjnjnu4d+BNgRtxTTCeK6
tncNGfqAVr6H3pbAuq3kcA2ht+Z8D161oFEZylU9c8LYtgQH9Uqfhnbbzxar/lI93YyUjTTcCJlt
alFsItuLXuDRqeRTOxeG7l55tz0fajf9ukH8lhFH21e65bLWr2qs+31vTL1RstJJ8HuigSRplscn
ITIN/FYUG7VeOYF1dwwEZfF7EjFHaRXC+jlh6zh9Ydnw1VKjG0CZDw1hh2iPJ7RE/y9qNxZbC5vU
MM8npe3XiPqPIBqjM2Jh1IP88pO9xptxOU4LRw9xw22iIv0j2rf6zwPT5xeeTVTh3Wu4dOfssOCk
4d/Q9d87mdcU94PvbaUz758DtRcHzbLhFlJP1mGdrqhfHirN7U0kkhwkarGQwAhlUCaYFAkZOLVn
t56s8ETwmLmGU9/xproipYr0kDFOUdKiWZZd06j0W3t15Kjm9AqNSyNuPoYmgMEiGGGJTp4uzFE6
pkohvxblNT4/ScjYUl0mz7bVx6syaoOArNoHVp+A06h+crgMcD+HOT3VoQ/otfsbdmYTCb5VinZk
iiDL60J/mgHk8MiMtHD1oyGTQpM1EUJDYccci5qWgg+gpFYwHm80mw1VGNimkUtLursTllEOoFCk
c5sU0b6UPjRO5wtFx9nDMNE/hNwpxZnWcqJhdVGndAeU61700QxnmJLA3nuQ50dard0/+jL9nDya
NNJ3gonhnNGIGIOEOHM+TTv0fR2b8+F7O4stwyW5oq/AN23nhrJXclhYTI/2AgS0d2rqNM77+VtY
6Y5ACjDF5/p59yzd37IFoRLu51wtcUZx5TenekcUr5wAxcHqZ1pOITJSWHUDsVO4WCs3gA6XiBj3
CgUVOJlJyfyg/QtkuVvPlbg4fyZ2ArmVXFDvUezS27G4YqGLbL1+R6hBFx6XmVvg4iKorsxPR1TF
4MGoAO3dLHrhhqOeoJ1kJ2tfVQt3sO2/OSyDkKD1IFU81nPWTM0lYKdUHU8vZ6N+jyQ7CLbEg2NE
zYnPGy2CbStbhDJm8+j5yXMeSGcjA53Ly+bMSyvvpKJqjT2FppdhE9srttOnXMetpuW9JiX4XQSw
oYZzWCNsjRYi3elVeUZg5Re70gm3exVYBDXBNOuOWg3BIolf8Jqm05pZDydoTi73FRcT1l+l/V9B
9GmtVLvZ1hFJ2U1sUExJrjop3BIqyG+TPh5m/CxW/jDW8knh0iAopRire4V/sj+YhoaLdi9gDWK7
ZuIsfbCKOjxbrVwtAZzt+AMZX1Q+p6JfFGWlgmEx3PzFXyVVgtdUsAYF7/WhaYqhOK2PG5WNy5c4
xyyTeQL5EOajFQLUxs7AMIfl7PinqeM3s3Wr0Gt+dmYm5G2HY4nobgq+BCGt5FvhU7z0E5l+p/MP
NGeffKQl+EORDrJb6IS/yAakZ29HJHxWu8OfkXS5gl9eSFMp07nGgy5Wg8z4QCxYZkjj3cU4kpJ4
fn+fnQm6WGVQbbOV4ukqYTpDtDJwx4YAB+5DFpUFlf3u0MOS0eO7obHMrhsKkaiVHG2/A0ZVye/e
9BzSydFCA9VJ1ghlez97UJ2a3lv30+4EzNEdnnNBAO5j5BNLyWY+zLMxuyWEDda8KZUAfy3xySNK
9lfqTpn0meirD8w9WZPKaj8H+WBDyGye9cVD4DdYy5s7b9ViSAXsAII36O0Nw0ZmxxZ26zxL5a/V
fLRfTe7XbfMujd4j+Yb9Ty8BtZVEzwdidDDmnmCwx2+flwSb9cEz7tW+yrhGRZ2HwGZ+0McC47Br
37JdmFyXjuT4LUiYr0lHJbIkQd4QIkOWxxOm+sfMaSX+dPL5/r5Nu5ECjSoD5ozhafMqzEUTCnKq
Qxfo/BoE/np1lvNBu+VSsHUebia6SN8qoxjHaMPrcP8DOOeRf9ccB0UIW2NM9+r6dlZB9bnZ0lk2
mfw27RXnsDPf3HJlKo2EE9w5t3jlKspeIb6H7oIJ0ImsmRC7FvpMxQsXyVgmYrVB0od7bkgZjiZM
nRB90fjZjd+fgqSn3YSNqJpfI0I20Xnid2vI1qKtNiHPZvqFaWaupgMPmcFqxDr5LPSCG4m5cwHl
kvkdLkNGodNnBOpHJ7BR8pXI0g/MdNQhviI4bgtdenuGISAP2zCjG0YAcM8lEfLJqZtkThRlULai
qwg2jmVGjlkN3WT2k6fe90so61GMkouvsFfOQBFi4kW/BbLhs76+fmjYWd/4tnuKsFcAv1NQUunc
HA2T8Q8pcQ0QmG9CdnuW1Q6eo7TjElB6zeoIsDBNZuq34pknR0q/vGlIWaH8AGjbXP2siPkJIPzB
qVMvGi+sShVBvAAxbJi4b2pXf7ww0R8O1gcjckbs4S7ZQpUX5msPAmTUUknB12o9R0dRgmo4lkHe
UZPIRVjE21ssavuNvm4Mtcv3PGZ7amY4ZI8x4yckHVizNQZBcThKCwO8W3krsg+ZyvAuQlnFrD6j
oEKf4wsidwstshhHrP3fUU8IHfug86zLVeCT+iM+05xLGYjuRicK0nbSyPDPbhKzNk+z3BkMBwL3
kzMOU1aCuY4AicBuCxsAc3ZxjrDAz2cgeJ6C9fFgeIGsfbZimkY+6TVoMI6S5CRsmq9BGb1AShY7
p+aP+Aho3IT8H1tBaK12IzIWFjwvYmdjx9O69t5fMq6jbaY+rxYGJTtz+JYFG6L3d++KhTImsHDf
uDPBXbH29vYKzOwJNx8v8Qzmy33KXdWxsq9rqwFOUiiR+t+SmVO15zF3L1HR9kSa9Ic9o7WfXXqD
LMQ2cGLbiSena7SHKdkqmfQ5lvcFeii53w1OUew5vD4Gqd7y5pS/DS1ptoxrlwZlNqnXHgP07CnL
kw9qrawXERaKwydGqERGWC51n40ftSYEcZml/awC8HJOtAfchmsGSwJPjBisfiOTrIoN6nhMtAHj
6Q4UieDn0rF9w8z2PSygHnQ3O2R3iOhZ8jhR6+cGuBFmBoyiHXrynkMC3/CPspV11OaIwX6wf0eU
7bik8GhXmj6gbAoD9SVLe9P2gFFcss4f0BEZYvd4U2SCw6M4iMQ0mU0OLnUvvzJka+8I+zwaPb4P
u/3gTgsffJouEGeCmOwm2A3vM7McmH9tkZ0HaNhItEFlKMSjAZZ0eZT9X0reUZHk3mfp0aGTSnwH
vdHuWr06Qa2I5oVxjvnthv/Nc5JdQUz+oTfKB+5YDOAPDtALZSSNJlDl8KnmKQDMLdnNsUak6k2G
RhC5SBm+BGwper51g0GcpqozhLGEjxlDWQVen1osgbSzOrWHXfQLukSSFEwcS3bXDYnMQbuDl3r0
JYFGrQN9YQRl/GtCTdBk3uVFhP9nsNd8j1pMvqR0XlA/jaUJeuBLEWdz1+8vYIum61zV8Bw9d9vK
nDxvJbteNHyZ/l9lXvozfn4MggGaLSX6gQjtWlpKIA5TqV34xo3MMjdzWegz5iFVPfpeSP/iTM4A
CpAcq2AN8tPfh3Wn2Cw+DIU+jK5RV2joK4LakWhWUpjt31gsRUNWMsRis9QAICu37bhnEJvP734O
s+Q4wh2RSkMU1Mkk29Nb+MX+BYbuc3bgj7k03dHjD3DA3C6x05VPsYhji/qyMWbUjNxUObBbFMT2
cz2RxDuMu+Y3FDQc8Lj3WqLLqXxrS3foivTy8VR7EZePoKAKYCz7MnoQnUSMg+6mmvN+nQrPknuF
jeA8uySBQ8gz2SiRu2tX6OOthW405CjNS8n2xvyM4BbG3da64v3eCg306criC5Avi86ZAl0Shz0G
R16aYaV01CPX7mcgIRAZvHmvEQSlQBKGegdCZC2sjH2wT+rrqILx+ObN0os6ZFyLxtk5vPSyk0TU
sLIuzLfgSlot6cZSrpBczWCsNszpOtM3zkV1RYtib1sNMasUv7XVxzbWTqqubPpYzKbU7w2VVrh5
SdQgtisQfCsGVeAHeXSbsBt2svECaU3/ACURjpkhyxQMyqcTybAPb4H6MEeh1HRNsi6dj7vMFVRE
5tbn0CiD1llR5/lpPdq7/Lw/VBlfIH/aLfBhlJt/BAEGkNrA8B9dwWKG0IyKYJ1badtuJovLXc92
EEAjSrwQB3bOvqdb4TOz+68f7oXnZJ1K5bF0wJ4X2C55yuVlg67wou8PIjXh3Y8nHMb3RdfcWDo5
EY+rH0W9Fsez+ZFlFjS5PVB8NMLMtClBt+ulKRbgoUi8IPuMnRLYS4Mz657VvLOPcRnjC0CxjR/U
6BOAiQC2WmQoTbiJZmaO1SSiAs378sBCelz3ald1fps90xnunAZtyvz89TiVhXznUAJncpAqk/xq
tRPh+/j8CyQUvnQ59uRASRzYiD5MxNDZMKKoC+TmWWhz7F0cMT5oN4L8qZ9S/Y+fEEXZvAzyf7ko
QJX1F6c/NYwZbkL3izLguxHrNXUep+RZTzAdxz78KTdBP5+6DRZx/HaE1340yNzJSI2z9JU/nguJ
dC+azPZvKrE1C33ynA9T0f+S2/sCtWru167fBv+++MQ1WDHgqlI+ouGhRn5AiEzs4sfm34+Pbvxf
HUXzUKy2XjrZofikK4RYPSYbT5ec5IcoDIAPyaJeg42UloQsedTFHsOL85/W4t3YbLkdCTBVkkFg
tVXdPeJgp6wTjlDg6AgTSbdRny/7ahY0Hh8LCd65TR0yUOOpzbN966XmJgy+SfVKFUSdbbODRoI3
6/gKL5bI8MVj+Ote+1KSx6LfdBgjNdH3IIb+A6Y2Vd+Bd+R/4txnMrzTFB+wJ3WOZp4qvWNhY/DQ
5hH56xCfd0u4ywT5HAyUQUjZ9ru69iAnR0X4MlAvxjlvU9h7PzxA4RMZ4J5rV6j8W7scrgxKvYlO
sYhef/1BgKKoyFcz2Fr6qn5DB8YIoYYyX9Oya/bRWsnzmWda45eSogq3cKtxOjNb6Vw+xsPtA95O
uYFr7JGM1Ic+pwc80/5rSUa8IUAT1lDNXi633uUl65K8kZwx1SF9nedSYuFE63Yp7UuyxfU0Yfqe
KXEaUuClP1ycREm/H33EDtChK8W3EoWFS7hplJEJotOsEml5uT5aE9oVUtVkvfU8r6KBmw+2Og93
LtnTw/x5E7ZUakZC2LfdbHeNIhFaylzQwX/g+WvT+yS3YE9qzA+RnZeslbYoYyqS72WP6RC9uFZi
yggV8VmOP/4rAc6y+iD0ca1CQL1awHBxIMpwYFYTYjIkenmBaJG+EsKYmDBuG4T/w9KzJAeaHSh1
rER8s1Jchq03CtK7TxV1DQDlFpRrujb5PR7arMTegRnZurymu1jAW/E+KHlbd39mX9tX8iN1ifpq
DIyG3ak75DSiits/JoCyl5EX+v+q458BfSsJzm2L8RttWEnvBPQmE2ch0q7hGSC/NPsVRS6FdKrd
FWxZj4cIp9wtBFD1TXduCdPGZW39pcoTt8n1iAR69RsAiVDRYP81WHgnFHqGCqwd7GoWh/DpObv8
+zAnZby8GTVTa/v7nqrCx1/HVOaabX/m+LBDba5wXXCgrKqdZMiziEWtdTp6QJJWDPJcghQnAQ+8
ZL13i6GBnn1wm8cgK310AnhXKQYq1u1qBNwTglrXLu7UkcXbSLxndwX0SLyJ6C9aMnn7RdyNALbB
/nRqDy5sV2NuS6Eh9TEu4O3yVgNzn/PulDnRnNvqoUFlGtOeK0PslthXQxwWtNSn/5aUU76VXMDI
dNyk/wDBblTmc/5XcH5REkP24LOlw0bme0VxIlxVdtPmGKTPSswYp5E4rLhorFlPeE+frYCeVrfB
aB+fmayPNosCBCFBxZk3rMszOxNVvbeXv+sG8J16OgXDrzxgplu9vz8Z2bS+L8RmQcdssUkxP81D
C0fhflWDiVo2xY5XZraCbp62pi5hdvG5OCp1CugUAycXWv0MFHcL0JVVqzER27Jc/jiR0lqKnekp
ng3ivpMoaslfZ/5MCIBEVilzliR2jgg8XsauFwwDq4Ls0Fufkq+t9pz0QTPMj+qmH5q0ByhXnu9n
GupC97bWXxHfMHOilCgwK692cebOBy0E9IQ8rwJ7G5BW5A/7PSOfjuU/wo1KOwviPj9jiBw2AIBL
/qmlAQnBRiqCyHJD4v/60YN+OAn3HLtS37WlYvlLhzbO+2sNe4705JTEI16FPVrLkVLUUa1dj1mL
OI0aBnLqeRaqGf0Vw3YrhFXSG9RJUCkQ4DdaSdYyXAPURoBgmimj6eBmKP/I/zvGGGbUzMnCVq9M
XQw53LeLHLKpAr3wuhmHLOKmpcuLTF6AWwltQwtphMKo8muQepYjiVmHMk6vs2Hir5WWW2TzbX7t
H7qN6dssO05+JlKtpuDRq18xCTVWzgsauMiB74VEoxEx4nTJ5ltddvAq3NhMfkPr+dNnfhLPxqYz
mhyWlwmo0PhYMZp1/Q56N1CI+Yvbumdk0ox9z67+0PCmHQ/2IUkNinWSY7m4JQAYO6/d2cj+3e00
jGavjwqquUJ9v/9hMSh6p1Cp9iYXG35aoYKCuG+9NQvFKNnyDhBQs+qWV9NRJ+zr7eVYnVjJcsXd
Nnh0nPnvQwS0naM0dAUS69hLpO8DOXwH7q9J4fSsHX9YzHfxuc/14G2Blc85BfRCveffH1NYtS/N
aLflZpe4J9epQ4thBfs7FlCvshV09k/27D+IESvjtZQbF0pbDTw9mCwtqOqBW+Nh7xDcHVcC4K6T
PKC51RVzE++oTIeHMH3JSzv0WPtAZe49YcudolSsMa2dtoI5df9dfuPJuqbzALyCg/FO+YO/ZO+d
5nuWDz9bEfGv7YF5w+/GsPR19nOK6BAqDR+PHxIsNS0D8DkNHelBBFpkiL5wvczWLcX3xsKemFhj
0xOUyVlx1WuP3FDWnGB/ZK4BGvb8DUd6Mrc8j2RdzH1/dzd+Asy4vGKKRaVLJtoNc7CSAp/k4Kmn
azlheFkG8/4HeGZu4pMZHYqS8wkoBaYEROHOYDvlmMI/5lf4Q7fr/yG0bYgYXMXyyWOBWQxW4b0+
6ZTKXfoXQfWYMGnUG8tNUmVyOSh8ojV8nWnNhntiU/B2dwo76DfFzK1Ycham6emZWp1D/9vgOnqr
WljR23AtVTirYAJxjrv4+xhMLPLlRKvhkJ/Nx4pHHppQ7Zwf9+9KIr6FnqFt4WDHT2l7rv/lbW9d
WPsLAvOwGloIfr9Zsf0cfQT0Lgj9ihZ/0zs4KQvzpruQy0f+EtjQVsFduG3F/pOQ8VI7TTdb4TqP
D8kB45XpgbKqoHRiWIm3zTUjNrTQdxc73Xz4lnX2LOprRpBqQHxVnYvcx4enUdGcHwQv2D5NNueG
SmqAJisPNSP/QXGHEor/PFAfj7y4/Z3PU91pBPfdaOXo0q7OD31JmmrFPn4+ox3LAnHwY6tL7gv0
n6A24xT3gwn21I8ffToYGgmLr9uAV60KfjCLcqEbjjwmysA7QJB/9WPDSpELu3+yGpYl/i4NHrc/
p6d94b7f6rBDN9HzQTQXAcFsejMPNtagnKz/SwuGr5VJv/HQ7SavQCiuowxQTp5B8mxZ10QwrVfZ
TWLVAUzBgQM0mS1xhPpjYUQ+4j3EX2DNG8A+QkGloPJaZ0BRkY8dCAw8Qyy5BZrKghsom4tQLCLn
s0NYq3MBJnmtigI6qQ12iOqKkE98ss0dIgNEn1/2MxQW1OHfeoxvv8hx7XyyCgec3aYiHNSZEPzw
XM3k4qpkkwhibCeannxvNZA9KTWBVkaC0i/s8wLyspcHWVGfO/iNsYHuC574UoUmnSP5J7xrDjN1
/vNnpLzDikjQdJYYMzxYnN25pC9rWF5E2w3F7zxUJ4G7ptdTAYbON8fYrgoTsRn6TntZyNlk+q1z
jePlhGi4pQtbZxTrlzq7z1pvpItVA45EXqljc/jq5z4uprFkeAa+0GCXtuEYEZWh5Yke4OoElw4P
7vTC158u9189suxUAp6IfWmwGckCWiOmT1SPLVwhn39qKEEhJIMHgogQiaEyiRHwZ3C2wBAqtbAJ
sFZaI7VgfOUjbSwxEJikhraC36ZRTOyGtho9X9t3ACc2EXWgp85+ZBMoSEesvl0wJl/9pFlY4fWJ
Hj9DniNpKltEHh8tVtBdpxv8t5rvSfXiB3H7/AUV5/5obtZ5hc9RYYOuajiFM6fpWB0CDpbSUFWK
xFiMm2XYo7zvV+VKsmAGTJlseZX+AZ4QLNysp81uju9aCMqwUzCjgR0+qfu+uCWpw7oMKq6B24Ts
LQcOul+Q9Xr9qCF/RGsuGc5/bIbBJaeyj02e6wtW6MI8/s7V9aftOf8J89q0lSSuAGxeyEv5kaCO
ZsOXSrgB10+ZdYT87ErKrtDlq2PyMdioH4yKSEPu+wiIYNSWL6eXfRwVHdbsaewCMVyxCdKDnzAJ
eRq5BsdyM10vCXT9Qorxje3fcjYplcf0dkmCWcGB47Qsh5tKlmq4KGKJXlzmIiCGCYQKBfoilQsL
ZRBVk9mSaO7SdsfCNxz2frl2Kfk+2GFWQP8sDnonz4qwbcvO/i2QJ50F/hqsdkzeyzbEP30RdDwl
stFIZwusl4vC1Y+atI9BzB9oLJjilWcRtrWuWXPymkN3eAIMWNSg02SDeJlXVuH8tgbsyYTFPsZz
tlgtlZACvjaOK5oRbnETO35GfZVG4Pjiys3vFRZDBoxWq6DZsQHlOt259HiJPwLW3Wu56o58g+zJ
blTDZRjx44RCQRg0Iav/0Ehnq7WX7hqWxEjY+9IJDvGdvLLWfpw77BGWJVDaIJX/qZ2oGXPUQgoE
KXhWmFfw7FCxoseQ0NNTzUKpqaRoredye5PV07dXsIjc9/6TsRkzaDM2Jqeyw2U2mhfX2Z29P+CS
pp8t54+J57PPzmVs9EpS0p8m1W1zhl2oW3NFB1M4jHdgTQt7XGaRj0i7h7CApnbVT8aIKXryHPId
s54SoFbC13FrCApC2aZwr7dwfE9zXPPArt1CmWnCPmsHdynBd3D9Stvrgi8aO0J9XIKGSNna/aPU
LoNFYw17si3EKJkl5jAZwUJ5sQL7G0Up2hLcK5j7o2yxiapV9RmSLOBijdCfvToZY6qBQom2Y6zM
edUsDywuGyf9GA58mpNpfrrsqWdYxgPrEZzosXrBehpXIjY5ucNlGgYs174j8ccIgRuV/hquatzX
UjmoY2mAABENyu+XTWQaRLXDUoW0CRTxlY/u5oCsjusMn8/seMM9zkhAQwpk07WPkyZrZMetcMW4
fJhaQPZtOM+WoTbLxrmeeBg44j0Lw6uuy763E8uMovFxpW2mOrQeE43nMKlA67eEVoWrDysR/pLY
QRQfl9zpwtP7Tb+fRp5Ca6hYHrchAvdl13B6PyYre9DeRK/kjoDv4PXaCpC+uolmJ+xQNnt95gWH
oN6MY8gVYLzNqHSb+yACxLUiyvvB02dU4CvRGjLYOYAz2Ni2aT9J8BkVOglYdn5zEwJyDufPcKgR
BA+oJllQhyAFfox5cMLEvSFuk2x052dySQRXu35+Sy86zmO8Ky/B+j/hCOSqAEIt4MOiLe3HP6dp
9zPcBnxGQbLSxM4wPq3n8lwaCeMzgXgKhBL5cQQOgLwXCV4vlr/m+e9ftyukq+0VKdb6+Ip8XtHK
eYYblekyAU5bRqDkHl4w30MULHt6RzZzmkzDEDL5dei+wIihhHgHnd+uTboy7EfdXmIqoiAl+t19
nRUG//6dumZSWZFRoQ1YiGLkCZuI2atGApQkFPETRdTE77tCFpM1hrE5kftK3VIQTPeaOtJiM7p2
/gSEWygG2/AUbM9S7S68Em0rVIlVtmFDiNIJgR2AZ1zkfo+xeShMttniSTXRIG5urwe6ygYKXbrp
C6dEwk8rI96JuhdLR+I3qAp0MVX8y+DpxwboubE7iCvIkbmoCPNY0ByYCOMok3hzmwjt3HcrHo1K
HOSjfHUh9gruRbIT1AyWgfIiDnVcnzi1tJX3BXvMteSNzp4EmG8tuqGBMiUq2hHRvQXQciNZ8GLF
qBWU4qU0nXaGQCSARuvywTvSDv3ffFCFSjxzYGqhWFtrHAavQExyA9VgX8ZejCY7pcCQhPek7IY0
devmnYjG1+Kv96X3ueQDtNK33DPArW+MJMwO/8UkKnSZ3461ZjupJnSoBtsg3HDISdW8iFPuTcF0
tKaDwT5TrtCaDmyglKkNmntz2+s1+xevxzcNWsYPqQN6wpqc+oJ9xrZqa0174eTaafw27BmPfW61
XRneOoMtGYsOMM7EBFsSVM7r89hYsnM9BRxa9rBB39p1+9TbuRrY8oxXLVZ3SZq+dqsQUk8AMUCL
vfn+l+RobWbvbHfHcWJqRFxo+BYNjdNIjxaqbBRAZISR9+Eqv5tb5KfZ6OLVtmOvHtYZYCy/Y0Wd
U0QePgVW4W4wNU/0zU16QuZyobx78I8XzpdHPoVDspEmTw2x0iHuvqB+qUZGCiFBxLtRtotPi2J7
nLNjSw38aahSghQ4sfILZm/XWFSMe33WDS+TYUwgt3gGzp4aY3Ev8EX0gBGGzGLjoYsczNEo4tTr
TglQrtmhFuRqmtJZ1jjjIbB4rI7TFfAsmtAfB2OUx1IUo981xCS1XQQ+IDuCM+X7O+lAD30zSC29
MmviUQ0iO5x9q286wVa/a6faG51/3v1NbIOT8Ee1dFKpV77cK1x1Bu132AOKztMc3KQi2/3HxyTI
pU9AO2w2K6xYOz+EKy6iprNXaheuys7cVwCJUMv2rd9Bb4bYGGCtyJM1Z8nYKU87huwHLQ9g3gd6
+WCRT6icqojy0ms7N+lrjUBN5Lm+a7Fzfc8cUoG0dVDH3Z6H8mr8ZcYZbwurD2VRRPFVwVX1r5Qr
Cm/kNMLSVU0nGpxdyRPgpdzlOh3PRKMr0po1XfPSO5+gfZ6apbXt26zgGoPFPlzPrdfTKo20eI1z
YW7zwAz9HOssXSttZMkYET7g6mjpn+D1M3nFEPLdGxpF3PDFE5eAnYgAFsZbLAbKNDbWDg0BglD0
qFiymL01JPtJM3ojYo4qfz5Bsd99IfFO5KjJabKspzyjGcbnwPA+0LsmfK5dqmq+vuTERRZWk5Cx
bC+QkIsg5sMp5eudarE8ARoo0nYIsSN8YCTDq9J7k7yqLXQmLaiFrDWRva4Sw8V0i+YWsg4pNNtk
k3+snAtN2LNo0cyDbRnDW5IMoiezZszAd3hiQPM5W7SrHCIt7Xnh38vpeJrE/rSpRng+g7Jz9jp5
m2GE78IDhaRh+p3OxGOWI0aVl38LVQ6M8dC/mzMluqbCPts448HemQusf2HMM3gdNHGtVq+Hkrsw
8YdAEIjhSu/Yjd2FVf3doxu+fnTlI0jAxm+jm/V/rhXrZ3Q6rAX0QXtbSzOTNSLGAjVAjvlZWkOq
VryZ8fr23Nt8REf1DEZzyP03zuvSHdk2cnHdKsc3pRIqXYGwfhk6n8q79GZY+PDeddq7EN6xWeWX
XILoIOyfow1RqMrYcsdZXOJ2t4Z/GF6abSQ66q8Q04Xmn/r44K01OagaOT6GipAS0HQuwTImoZzG
CLsnrc9mzpptlT/Fc8LnRLPwrcXhVW2jgVkRIFrNEugQhGCuxMaMQoY3wht2eKfr/Fn8VCdtg7K1
OvHwvKyXuOUfuBNBpmifOTU7wNTgw44mv2ypM4PdCi3znFwlEzWX10Js7Q6NYvOr+sUKpVqIw0+g
PrN65DqI4L8ZtAcaQucbrzA9GSLzJ4mLdcFSJ69QXcUdGDPirkkxJs5hmMmiXhpQaC4PpIghZJXT
YwSAdIn5SJGwO/pGcwhSYYstgH13pfj7ys1hQOrL1scYZvfDdNOBdbTmPfZ0h7/Ch7BLkp5ZPju5
4fb2YVjT340bptcRAEAV5+MXsxq+xvMicoL2hgxcAYJH7btud7HlIy2i5sSTxl3XK5oV32Com7HP
/tsx/8qPdyumhhF9OI1MP+HVrWtuPabn6RBDFsxHKzoNi1UYiqudicsSw+1cYfvbXPBNGCWdtsFo
EjC7p4DWyr5cURKldUr4oQ0HOOjhF8Z7ki6VCZ0rFDM4hqWxzn6Z3ow5eo9ctEDVJKLKjChX3MSh
eUkZXwpw60FfIFY8UJChFfhC8oquOy8i1cPQwa5SPtNWlEgZPO1gXKFZzSn8HfbsFKxKvAghEMPy
jhQvb5A5QkwIcvzevg9XzmXoaQNjfG3FGbuoh4IRUA8QdYByPP0SIrXQj+fGP3IQ/T2movnBYbKA
8Kx2btXuJO0oxXa4zbcoH31j2uKjWRbnBp7TMupcrkUYYc9ujwhgr00WxAvfTWxYuwPoVwpyRooM
PKq68ZsYPZ0otQi3z3ODr3JYj+87lp+oMAIehYd32F2D1sQ+P4ygaaR0Kv2rLfWrd2Pzu9ehb4ZQ
XimCkVa17yPNvnfSQ+pYbkE7YR+lXCT9PevtbHxo+5Be9N+sSFEfXzCbnRSrxY9zP5yGak6+dvGw
eVkAGRf9fFgVBI4F+j33MZDCNuvwO6ak4HwTr+4U/DPnRBvmbZmxb0KJyzvLMezVXJOknrqaH9b5
hRP2LJd8sxbNELtSeG7rlrDzSaw7wpbSN8AMzLhPLRnnIChY6Na+QRvMw4j0madGX9ztTnKZyt23
93Q3DBo3y3IQ1+WDo4l0KCVOtHY2CSu4wVfpVFrpYJP8PXI+Dt4gXM/wFRc6jcMN3weqssjh9c6L
m1Kck9J065C24wlvLpaNMi/Ui9Df11p8OmIHYUOcDKto80PQnwitnN7SbaWt/lS/7HUxSAmV4IXt
6e7T2z2HycZS1TDV/U38QLXRVBvxhKiZGFkDROd3Ma+mc4FiHGjdfnQA5pA348wQWQ3Xjsu52Rtg
qFtuUwFpfMVPVEdgb9glY+Zt58DGvVvUai+GVteC3pRVvky73IfYa5MPQ/0zf5VRcwdXW19qL/37
yLq88dEFPYWRtF3BK1g6J+XydmzC8a7nLv0j3JtCbUTQj/UKDZQh2JLFVnEpstBjgVMmpbtZqeSE
GH2Vl82hHBubfAE11fZARPBgWpkjESsBNyFcgi0J/fUG5oKm+ppln8H8MFlXs6YNR5T9cZ1OFaip
I45dhuqV4vNUJZHRUTkXm1ZJtFl8sLJts/Ks1nd9LX5W6yYkPFlFOlzSoPd6ekav32WslPlXHot+
IVPVDdIUiyLR8VKsbfZ96dqTasFGQam/Xh/Ihxg7TOoPdlHHlpPMUtYhrk5tkHziS8AKon9I5JjZ
11MtbcB4aq6bbllZDCYZpWleNQZcEpuxOVaRxt8McIyCN0glvu0/dU5bAhBEi0YLrWB7YS7GZN54
GBXsKidtySysqePysiY/Mprf4XrN5ktIhfeXdAGX7c6vfcd64ss3KoldHCDjIj+mEXbjeXqMQR5k
NFbizmDLsqLHp3piLMAx8DLjybePjd65cYPCRnbqwis/QvyIvULP1qbZIJCvHdkaFpjZdy7SAAkF
C85GXSLAPWOCqn/7DATZzsscTY1aJ48tCOzWFqBdHi/9ojEYG0BfFjDC1wK9Xn0TscpIDN3riV6R
K2JD7TrqNQfVp+yvRkTenhM0pSk4/kkD4x2uXeF5dLk9qtz73JP0pZWhpoGAhtIaKKdLMq2pnai1
rtfD6e1T2zG9qlsOtvS4k0cQWHiZukftJHGvg7lkOwz0eApaQ87DDxikmAY93uc3pNQiQosYnFB4
X/srr6p1Ntzxu/HCjLgMmnMSsEc3Nokre2nBKQk2hipPO5Ge4vAubusFpJLd39sEDioNeZOCCzKL
3I1pUCP25KWlZpNStajEB78RPB9MKyu3QvtfnLnX87QTm/1dxG5axMIAnFaLdfEuOP92RGepe/nb
1JlTjdRghaR4eNt6HS3lABXtid/sOy2QVSfYa0jHT9zrAXRlY3ov5GgKP0vhb7LSKzzhyEaMEhWy
RfC4ue+58VwNYakc++QpsF9z95mlUXzYIGPSvW9BFnHY5+QA3iZ3oqEO5xigI6ICA+mv70Eiewuv
688EzqvEZ8ZX805gjyhz6YXQR6Lfw08RIkp56PHY4bswh7Gfj84rEXDN4aaNYBMpOLgk1VNtiA6M
19iDIAWnGvn9EqSJR12WexNN8ezMEc3ak2MumWu3hHdKnUUl0JTg0m9ozLrcQ0+fqGxcjFA0QdLA
TBDLEzutOKJnDUyp2gBNGobGlCj0CJ3KDwMzAQ5UiazQAls0qcsTFCKaJd7TeejabkAXs/RhBZde
6vdhfu1z/Tet5CJxS6ulMfKAovd4n+B02++neKFA/N5JA2dSvpHVDoYIFDD9L1dJ5/kclcN+N3eB
xXd2ZbP5C4IzX3i8Ck4JGY8ETRsGmOSaAEhqaeEdKj7Yyt1FB7klusMBUeEwONNTR5lV43W2XlYP
gFxo6q4wpBh25ZpctFUDwvjYGUq1dCnhui9iI55bZrnuWyAKnNPmDGsVSOi780Tn6MAlPIgxFxCD
ZrAdkxG89HOkmMgRkHcmdpDkphRWbhmcGBL0jyxsnRJ3Gj5BAP2MF33rDR8SxYSKp4pfAHt2NbXx
6g7A2WOQsmwHCZuxBHk4r+n1WRxpp7t/EbpvUnZoYKZdzCyXOfszgH+yxvjoPzt1h3d2PMQS5ds6
oKM1vN3ZHsqF+7eIOvwdZkaUuFI/rQpbODyiXjnxpXIw+vg5X62wP5t20JbxYk6ZV5SO6G3odi+J
4o4mCnuErl2t8TXyD2gL8utTH0/DqcgAVBbKl9VPfmOUvolZRnzv3tNP4tUi97eEUeDtXG8myAq2
9FAzSUy0+AmLAbYDivXK2NG5om+sA/l5KEAHjKb6bPlOgIm01LEtvUPNaOp/8DgZCefuyv42TZ2I
IuPShWyL6+rRPfEnzp/kiQSngyOG2nOvxdUAGotBAJr56zJ3LKwvvz13zQOYK5JiN64056ojZy6y
fuLVTqQl05VXdpoTmfQNr5wApil17NvH7V+bH9cGKoFSSn2XSHeJamVspUk7XDBmk2QdIHqStkwD
nb4Kxs+ixwuPuWyqxJs6jlbWYimqCyYMedeWz/1yMsm+2CPvzhi8nuGxbPJWPungbwSbHkALqH63
v+Msf+BPKgFUISPHyPSvkpsZYygSBncy489GbdWh6IHBSVLyskZM80bsNr5+5dymjQyfbpbxhc4f
eh4Ou+Jz30J1q6/rWPzIP+GdlrnksPdyaboIjSSqGYBgx6DDDVaPmoyazyTOdW5zNyDceklPFTe6
k/HoEovytqwGwYrKjYqneVVFSbeuCmu8d8lKEvWoIuOIbpThBi8IRcJ9UqZ1lnKWiyNjLXpAePJY
E97JVArcBRdTofsYB6I8sIq4tF2O6v19CbOD7g+BKPumdTr8P7td7k3MKBMbdgNEf0RKNsR0J7pc
ZC6t+xLNG9bGXlDFsAJ5Iv6HVj/4XRDHb5UqxlLVB8A/ICyN6YZn6EXUHuK8vnro4DT+z2IluKqq
Vy/NF0Uw+yex8+HiNacAoq87UzDsoyIc9mYSDtyRx3ZNVhYWtwNwbc+XifhRpaeYGr8WUf+gOlh9
GzwIQA6rjVbs1mPxpcZsiX/C3wBg7ygwcaMdWoXUQNHiyzChWoXAtqnx2DOcyo/5PfOvVTVYIsau
ZMgFBEeRGPEhnEhAFr50Y5CfL+Is8JxOxs60lqeRqg25PRRdJbilKJUw9JpRir05q9yDFeUgZDx0
76huG9VilCIShEV7Wfs9APbzj0pYZ7EFV72f12BjNjgVuTfMBBKs8gzgsNn6fLABxJJ1ESIuRkXK
k+uJd8Z+DagysFvJg6EIcbCIO/gakzqgbKNEFU+hr/qov6HW1HIstRbIXxDg3iPKQNncZ28DfnZB
XaI/42qCzh1uR2Yr3K1FNcTkDMQuzbX3XSCTSJ3a0Pq5dJPJATXEUHPYtlG9MWhI5VBRc5LBsswl
zqpMXvItg8vK3rnjsIUhIar42t4AleJIfB7Jfc6daYiceEhc+c5dLmhRPj7eFN2vVH8wDCI5QokE
wPQjFYG1js5xBxsefM24NoRbssuu76NvyI3alTAoND6WeJQRNEpgrdQ6sfWLV31sJRaeBh2EFISY
RtQe/zqdpQMoTBhezsMz32fne8mpcBLQVspK6Gz9i8VW3PMP+hT3WolhMoLIUfYH17l7IMHmdqOl
DIXpzj8k3YhfWUxhzcB9EjfJprkRminVNXmD5RYxxT87RVF1Piiv5vg2ko+vk5WdvAwgEH87Nf9g
3dCj7GEUIr72RgFhd/l1FdZR52nIz1XOlTb4A87eqEp55K5xZiLnLmM6D9lEbwfqxWKU9k7Irr6Q
R2vCuFJjGTjQJzyn30YGQR6fSWdf100TWkadmD0X40Su35X1CKh8QQaAuAP9dbhnQ2p+9ujiUH67
O2oNbdoWGvHXt6BQDWwRFJhs+Z2MUFD08bG60W8/eMTG3pLwJjaTMMomNT7fcbrscLiywMO7MoPR
jvZWor7WMJ3grZr3Pb4mjNuu2/DRmnGJSqXxUQ9Yi8QAkPiydhNtlqeYLrh+JQN5LTUaOzHhzt3N
WN+lYsSOMCQf6JjiiVCGJM1Ff4oh+KVjkZJTjjCAwmFrQLXg4dghd7HJb3PK5XWpF1GUo7Xz8j0L
frYRY0VAIo/U0wGydZvjrFPK5yH9mAm7dgw1CdW0xGIh/q/8LdIGgJQ450cNwSMN/SMfM5KgbkXJ
mE2z35ambMHvPGgt0bQO0M4GPoIlgJDk3PiAabqE8Dwm/T2chs03pXLhKPG7hUDGDJe86vy+wAlN
iXwbWMu4Tj5nqfiTxL5iEv0wbCqF0WImHImHiuBso/MvxXsPej5U9vTaSFj7d/mMkPAAS5it5mon
iX/JfwM5M2ENYgH21MP0ePFHTprOnsqtMFIYisspt9VspGyrfAsS6ZRCp5s+ynnto1hpNPhcKZfa
M3KaJ3nYiNjX89djlmFUpCntxDnLXbYzobo2IjMJOpXgBFiGrec4gjd2w9CDrjrLYTkY4yHw6yNH
+m4r5eVg2POcXhhdiBa+GzOeGB5yi52kevI/MrlD/rvQbXCaUDeQq8vIP/eYnm5SsclFwcAm1EYP
I3Ib5I5u+hvbEWSAA5m/swe+U4zOfS8ZgebXiEAwVoYk1YQUn+ysbivQspcjW4Y2Vz16+WQItTbE
nZzgvpW54VC/Dovm2vmCPTkgSVBYkJ8czkxKw9ZupO9dMW/5HewOa39rBlLyKe6IeA4O/KoP6ymz
2jgP4s8a4awE+Qu3frQcjWA30n6VUvME+6sP8JF2Ejpp7fiXOJKMIRd/W9/7RCgcGwKWIim4IjJB
j0nX15US2n/9oAMD0AtTJZUuVZp0UNJVPx8l8eh2BdizUuMDe2MHWTNs0RYj478FI9IW/EFQLIBW
GLxbwF2BCLOfOUY+ft9Mth0oGzyfr2cdpdLenXkXtCcLFjVrortBWNhF/OZvCYvBEFZHAK2MYcvW
vpDIKXPRx9Tt0DktD2CAZn7jqc1lwnaZRt9jJsWxgcJR1PwAcXHDZGRru/r5ED9wPOh6WJsXpBrl
Q1V3dnc5JTXZuJUrPYPfpMeDk3/zbaDFquRUlN7pER2EAQWGpCI8AHQko2p/VC1a99XEnt6kwvoX
09trCClEep0qdjmpRTtQM3PTe9tOY6SCN7bGyiImfI0bXfSdzPKZBKsSUCl3XkXKwYhnlZuTeSj/
3b8FRJrylQx3LMZyrMOS3tnycnACAUjqpT3vhKVB6FEE0Nc/SgOVNbO9ikkC/iWRcGMofyWq+2Zg
MPo2+oms2M32piqxxWd3RmFyGRUzvdIz2EYkFBVJrCXLA9QWfH3cLfI87re4KlceJsUBN+jMM/Hg
bKbZjlmpiWtoLAkUGoLYDfTsmA7kS1TfxeiKVjU/SscUG+TDKYFws7SgvRavsyY79X+uQmYQZgzj
HhzXBP+mzQZGg9ut4nHeQcFg8w6RXfRWZG9Siij8IxNoxPxr7Yt2sRI2y7Zl0HYBWm1EUMOWaVt4
OCr9Wr9byaKXg26githBxBW4hamHwhIgsaJIhYxnYp2f2BRK9SUxoNXoc+tBnYatVXOFw79x8RXt
bdvtnkXUY3rcP7uP2ZeU7bvzAw85bOZ9WHVTBVhwv6gCNursb9Ldcw9BKoBEwVixSLv+CGPFsvVG
1S3x6nh2+WqqBd0n7NH4MFCJF4Tz9S0mEnBNZGAopqsE5S7kOKQhlJeazmiZvswPqhcHzmfUZwme
Ib6ekoGYP/5ZQJWSZ0K8JbyLv0gDWVyp3oPjUzmApKpNeXtj1tuv9P0/qu7+xkoXKmZ+tORHFEp/
91aevzNQj/rbU+xu5g70lMwtTf4tsoH1GGuvqQwB+pdL2YrK4kDu3X9nBSCWCL3QeEIFODVaJchY
qUdAPncLzSzLsNg3ynHGoPTdXlDDptbEgbLxI1vPlQ9qu7Ntw8vlBLmfz3tN8jBTsXW70I8rckFA
ucmCLOiLpt5+mpfrizN7MZ4qWAJk27hzSmD5XT4wyWAeQkEtzuMa34GSIumPr7eqxUzrf74QLj5R
FBQTQAnQnj3T6quxziNKzuemzeoDmP2Bz2p3/2tcJqa+RiMm0zQgzAawwjXu1uPvcrLFDz4X293o
kvZdpZpMSSThR8YYIcapxepp7YhLdJaINpwkhWVV22E8ad/+zZDZbAvFadnAiW+PlovuaCyLQNA6
1zmW74mcs+d4Gd8K9ZnpnnbDFeIMUWvyNxkI5aF5CeP+CBYmXiIyXy9gb1IKjIEb3nmz5q2aNYXo
gPyABYUzCAX5d2UYJeiMhtd6l5lxx6Kxrl6BqYn5+XI/OutV06wjG5hT3TxTUB9q9+jLhnXGvHn1
7nvyjHijxtsGsKkLQLSJaALE2mX1bW9eYNzsWIr8XykXdnxypMZ9tco2n2M9zHKwSix5h2e+5hVV
nTHpqlZ03T2rLxsz/VIb3gmG0w8s7Hh3JM45cBArRZkASjKVubVyE7ZLNwjFrfqe3wazrLL390oW
mIxa9qCK2n3dk+wXEMGwwuv7YaaI7JhrBWQYM+CIklIhhmQ2SAkiK8zVsAiqCy66+JuSgtH1e7o9
93PY722L9mA6IMRcDavqeoDg316fgc6zNBQ5P308BKxIRsMzDOxiQzu7aVZjdh/zOXH6UhIdBGa4
iy1EvH9VczF99vapAluOj2beKVssmdWD7rw/qT8aj+UgWK45pP+Ik4GyqRzFAE5pCk0O7mbTilEv
DAp4yHM/JB6qT5Sz9qRr7JBig39cZxynbRF8fdAi7nHsIh0lj7D209rRb6+bLm2ur/u/vwMLLSVq
AseeHQUIezXTzaE7Vqg4IFRiC31J/bxgtX28xN9ZuaQnzqSzHu9SY5TnnaCjKuxmzA51ATK2P5yE
KXk5uVA7Z6J4tbQJxZky7Bm/BUbl/4cQ+jP9CUH++jJTQ6WSNk/Ne1nCb1b6WI+eia1jEXQVRYiA
jLcNHG0FLFb/rNicEl6LaGB2KRfhMsu/O99XEOoh1WBlfYZSemG0JWUMhNgFOAQ3z/iAKsyOR81U
+F/NQHg2YS4H7VDvsUfR9Q1DK+fbavl1kMWsqpqW2rDxD/HGa/A4HpwT28Yxog2Sc4G4Gd70lzA0
Kr0t2vZeHOMuACFdcU11lleYJl4MYiRnV4rxbApF8SiQbcw9Pyv/Nh5lJSGYxzEbN7//G1yTfbtJ
DdgicUFDXE4ZrEjlHIDs0JIhtsX++AVSbFcoZhs5J3ctQOos72TF+5MottmNN5ntDiMsHBg/1bah
fXUOusw7+JzGNLDDzmTEkKggZ63F2nXJQLOE4g7znB9kixMTHfQ22JzcKuToay07p0nJkE/kq2Rt
6kte7FJexXE6LQPPSb5SBTRaAD368/aTlBBm/dPZzhplm8pxLjcfpZLQog7fcc6CaI3zkE96Msik
UW1fslmXjA8RfiXySFIm0tMpxVUt6IanerrW0ykALWOFSZc7gDO0Gfl+geRxk4SpJv680OzedZcm
Xmm5KaDYtAWtk1xVsaDTVD1TxMuhC9zcpDfGgYy8CIZwwvbvD9Kungu+i4bR/ocjgoJf6Dg/qJP2
ZmClwNtBw/7W14zI+JYU1fcNZCnKmABf/yDpfM2ac5k91e2l2Qf3VFcGlXevhCEUQrljELAKjT6E
nX14qOEnozRxtSBZ9VDtm4L3zQTSvj21ZNGdCL3SfUmbAuxekL9edjhcOYYM/4u9s32ld0f3p5Mr
6IaprKBF3ZdufxdrbfnxPX3AiRpix++EB+8H4BSR+wc2qWiWQZx/BKRfLYXcCI5sEvNgUu1MeMI7
8ZZ5klNydgHUvYzdlA3NDcbF+hsrwtWW/pHMC2fsMPnwV5B9So98nWqWJ6zKAgxWa8Ao24B6SFr5
I2K+cYvLmKsUdoCz7quzGnRst44rMvtoWWcQxbLwcbwVlQCuT3kg7aVmUwU9ErqyF1pIRE6cOjdo
ueO0s7c31LcrDwPj0tVWxm7brezUiUeO+zWkGB70XpvverITkIyLpAa+hBzPrFOlxt3EW3cAbFIK
HKUd9HMNzKyh6xRvfdNzPw1Uy/6uFsFPzjQlAnQgi2nBgEn2JeTqu+1ZyrTmvF5RRgF6vdYsBr33
SEB66CpItTMSx6khA1nDmG04SNkGY30U92vwoXFLnGKypBHJderYAljX055TIvaqDlAzYPe0gE9i
9qyDeUSx6wRnotIuuK9xaoj0aLjFExR2Ep1kk9UfAHdS8qG1knZFCUshSDYVlDwgJA3HNSSMbe2G
cGub68YWb907GfHUMSiq1z2nX2IO45OaZTMu6N538Ve46zLtHbK+/q+JEZXlYAgmLhbe5MmRrYW2
6ENMLmVLNSV3cpRZUTTkY/vhjGbZjhm7LQ82DCQy33DzQ0cJskhVKOUU2Zq0wiVilyP2bZ6harFh
DJsZltoejDgvyVnRDSGvXHTSBSlmpEruVTMuqdyzHTg5lhNKH1hpz93evErtDW15qjfNfSBbtcJO
MvKBObl/QdkvtOQaxx+zpfHS5RJ4UGKBSXaE/Iroq+t2TbfrYMkmBp5P4XbGGU6diXEfqPtgYvma
nvB4RSYnJRm7RMcZ1EVdlSCW1ldljx1A1yq9Z8E3s9Th1nK/jVqQGMUj/p2/XbtipRCf9tEX9UrD
be38fgigmj2NnSiDbJ2kdHdmX6cfAZNvGgIQa5u+a7DGA4mZM4RGX26ydz1F14NU6Z0uhHCYnXMQ
HFINeE3znmwzhSxAzCnOo9Qno4+iynrPrJsQjqGnu92fSGzYSjS7d5kJZ4c9UJQ/tIVx/p5dtkuM
5a5neLCzzj52kQsTMqVtBWA5JhwqZ3uXJmxWSFcfIgGn5ALfaPyg58s2HUGWwb/gcZeYAIgl8Cs9
ugVGRzJpD9jbwUmFuFFnnmBi5d20YpwXqf4Ju/5Ir8onnuTUzsMdkfNF9y4sOkxy/D1FhVvABk07
gnn8980r7nP/WgMB9sKL2iNcAYEC++ebAc2prfGdLgpBfCbL62chOegE0djvWcueZjZhCfCdOibi
mKd4P4v4kn0cgL1ujQ950lpDdjP1HgeJWgj+0nMT2c8eXM6YHkvc7qcxWzh5vIm2Ws0gB2muhUsh
/XlaBZ+dhuZKjTnGDdlOMuM7dIYkdMq9umwiNppcFh3S2gRNYM+xjL2w6iXkkmEPvB13ZgvOz+GQ
pRCXvQ+X8orHEnMe6WxsGHWAhNivYMzPxRgNBMzwnqa5CC04V5+YkH3uE5NVQFjg7qTuUzoy0fO0
pqVmvBxQtP4cSplpt6bUtOLcfJoO+Nlhl/LQdFbNPHnUr4oS4nN8NHn/U1ti0K7gPH0bQik5xzK9
LRkeVIlYr+zSwui09fPiNVfCHlxCvrbHXbH1zfOz8gQRefu11iHbf6RqSzjh2Kogg6RROPejcSQf
lWEkfj91KjvR8fFbnUK0xjtHKHUaSUSGPeMtd+P8Pu8Sc/ev4KWOfM5V0zk3J5lDbu6DzvlFOmOZ
wNplNnh25CDHlKxrzRSgSBdfeJ9iJ47b9Mx0xgM2/gWNE8Ls9sfrjt2KvyQfBajSzh95xemE1ID7
vEmSNOmkzraPf84gt4Sl9FzPFwxt9CuR/hAS48z+zaBntwhDpYwYcdH4J/ReZxPrIVYr/XH1vcAY
gpHQTA0wAaJDSCqkfmX9pqSGdD/rLMkprhR9ro63jl757fCUrZzRuPwQ2k7a3QQrBezzZSJm8Fvk
E3lXjLtiF5nBs9Uu/YeKog4TKs8t+O7HI60zyha/q6wRs67GYv9np7NVlPA9Rc0sHHgHX1j5lA2Y
AqtYE1P4M3SroBlGbLOPHEPojfsleHnqxKgXevnkZRrSZ/QOugpCn+bE/ClnbZoZgs8R5CQt28LP
KFOt4O3Y+6yYlvSMsnQO0cun5sR64VUc7g7dfSTJ/PTVqImBQFO7cysxlB7ED0rcIr3kMkJVBrYZ
lYKZhZFnDHPRO8BDBsnUX6uFPoApNAfS/soJf5XFRV6sTCyvfZC46nyR2sKjzHFz+/rdkSll89RX
fII+ENS+053/v3jg5lwRJA9fAbTH0QKJHtGR+DFCQl/zSta3HSywp3A6D1EChEVVKB2FQ6OX5nh7
qPpFytI/shNaBjNDMh6oQIimn9OWkwck4sptO8WrvaBHVEYm7JrwbnUEt5I2N63ITfBlbO2RIZMe
NiRPJNqvgzMNfhDnOShzQ5N5n1ABGCupPE098UqqujS6JFIxVtGLfHjxENZ7sJkBH6bjgwi4Ku0T
12r9i/2tVktNxWICQDYd4Tgwi4t3cGMYhGpmiWLUOn3w/4G4hjv2uOC4WNL3nLgurkB/L2lM4Kt1
gtBqPH6pVIW0rDmXKcPzwoW1PqEswM+61MYLcsGr+ZYdLxUGojVCkS3yVwb9oSaEVMZIyUEiCMcP
qD5ADYUGikmMbt8xQWBN/vh+dxczS2pZcBEc8GP+0gYFhuvcK8QUwKi0KdQ74ZNaGS31Dwcem3pB
k+TIxaLRwrFiaTkORhQxItMbTfBbpQ1zQmdnORfC2DAZp/FBlRo1EvMEu/RnrX8Qd9v3a1HSzJ3M
sRrgRKDl1KxdAkRqK6H4o0FjhykFJ7/+SewuFbcXcC83kMdEQjguCPL6wbLH/jo1N5lrXLwAIlnu
SUz7lI6dZJ4wUsIDBhRpNZ/wp7Izc2RVz1VLpvAL97+mGxr+Vb7HI/xwonjH+3xZatqr+QuECW8r
zDvn/ofDGm0jgi52n8OwwqZA2QNbFPeMzXRtld1lOQNHCFemaTXcCrbaCKIeJuH1GS2iCvngQ1Ix
lOwEHJyTxdQBPJVC4G1+O7UiNDl9at9swEUTjWg+PVZ69zbqip910tntGpHVlz5o24YULotmLq78
TfeYFoNd4hxPowsFsZgvxzhJ3tr9EVVswx8PSKW/GeTmKqRUYggyImb5BJsrAq53ZzHmWHeOzWv+
ObED/rx1Jz3JMSjk26Dw5JsYpzSX3rHrVbSzIybTuSseDHcnn3rbuDQ/PqTAqHN9YxzOtHLA/+Vz
ODAUdWCg4eFR/bZRglLnMB3L88TrokKOpE4KW0di7yWeSKZcAkNE6mOjN2lWKPGpujjww18PJGln
69Ke8JiIniRSrk/r7vSskH16sKm0hmwg8CxOMKM04wg5l9QwFovBCbzWb4yJVWPBzqrCoUCrh5WU
1yzMwVV4Bg7ZPTldJrzICrHyuUSvk9Z09wbGnX2jPBIdoFi/2BeojbRil0rGojsV0EmXSEGTFSPe
J6ybIq6A1TNAamtbrDP2K8gfT3TwkNGcFwr7zR+httstXOMVdRXiWN7snxLVLNP3a8NRPE/0pbjQ
JG+Y9jFrlbgFfE6OUP16C8nHBpQt2HtCamClqdOG9R5V93u9XIzlqqxiAOEKrO9FoDkGiVEU/vzG
QloUsObQMP9JoP986zBGFSy8Ad0ep0HCvLYDNi07wxwG4VjdHNgYg6DEyScUf0gFypLrtpy0QYou
1Rab8XMkj5wPKnavumkHPfAUjMth+DAoAgReO9slMEAKqw5J6vI9/6X9nI7DjfJz1B1JzzABLS1z
EsdrUBmfiyh1YjGzPISHZ4WUXyVmC4q6ot9u+LeacrY+5vO/I7i396XbUi4NtVcPgM8K09m+nnXP
Vm/jL+myaVqAnD26uXpBTqiXast4H9d0jus6LTHuA0E7MjbzBHkiuII6GWbbpKedemXlHUogPoig
cHM4R8Ege/QLPI4Z+quXSx1lt9d0XwhEWnPp62YudF4RdHPJ1aL5UhzV2mg1SEd82gCZ3wKGNKjh
ii2ild8KIqyWc2t28SS7mltjBTmDVjNGIBrpQIufwRxHvIHmeYnILJB8VQIzhVru7SqBLuIVcouq
5Sz6sKgyMpDfQ/SFWuNhjNoPiEsi/cmPTqiFg4hBGh9FuSAO2YEReVCfo882r1UbNvyAdzhIsGQK
3RctWIUtIoYTjtDTqTMtncsRiJXuegSQPCaCEiQCXy7xXdfvr0P6EVlVpVDuSKoNR1Gs1XMF14TC
kAFYgAWmKSfAKi7vnWNLimYMvLVw0l82I84ESSoqmgZYJu+32rHRH/XG4XMCnWy+1Q2TUnoUzzuO
TIdxI76hQGFOTb/p8Dkb1h6wyRTEthCH+xyeCSet7p0SHrE9d+Fpc5SnjSm3mc28uEPan78Wuujw
SIUYO2NdYK72mWH+7FYcFa5qka1coAaOHGsvidtPdjQF+4yL4AodJIxomc7l5ZWYAylL1Obwr41u
rUhBMcEAL0vQsd+iKK13F79iPBnkfwlVHuEUjfi4vxQSHLu7NOLmh8/bXlaHK4MgFHe4YqmaDGR0
iFKxcEM3/oWwR+mVcbpfVtfHQHagAycesf6CvjIwhzXwViju+Aq9nzwP2sVWRkRYJ8zOb+CURjAh
sAtmVOHgKSFTOBu0rTfqOr5i0uc5+xo90YSpK6hyiJ+97ZP5MRl89fWSJTWZYLsmdjaOvjASjjMk
25gtRb4OcfCwN1D/spczVxJS1x3ZR2zTfDlogoN77lOmonLOP+/W56kJO7RMDfwpL2NSPSL1gmr+
abrH+4x6cZ4N8jPgPqHti6WNZRP4cqepnYaotB8sgUxV5hfugvI4iQWNZiPeRdv0tWXeE7toTSBW
YdmKAB8akQRBx2zczPmzbKw551m2CFBtRzkL4N0NH6g+RluS1akjGYQ4ZqtvRRGVCkpdHpBBpwl4
kyKkpkD2xObmOkNQwKJDA/plRt43VgmjucWaDS4Zm8sComLSgsi0U8xVgWt7Rx1F4eKBMOar7CYv
0hep/6UQfGaZ88yExj/bNTRw2p6dqTLmWygZaXjy6HGDY/BhJgtZrstbrwjWX/yWoDdx+EcXH8He
v0f8V0/l+wGQOhpvlgjaudm3TwAyzlWpw0nPBKs0UeDWw4eFAIVkobIrjmeVS5BJj1zh5CzAHOSJ
tLUl4l16urpJYy8CjVb0c0NCK1EOSNrbIQ3GNtH7NKF2+O/v+reCMLHNjORQT+040oJwlzIn4mUM
Ro8s8V/ERqmyC4fDbgMnuZElBoBCA8YK5qcNSQYIfVd5FWyNjVfS0ofVOOBsSLdzape6vC3SBCAw
r+dvysD46xQmc3zmsyIOEmjx4KWzcA7vwbtGkkDy9eS3RMuLTEjT5Ypy7HkLfiCrWyn8lhvAY7tU
ahxNFRHnVbDcF0SGMKQF+nznWgRwTq66l9ikdPu/vvY5sizMV4qvrmu0eyXEB/f7leIUzpjNXLDv
M4GnVMuY/TP4Qox3vGShHYHj5pa9DucSiKm4XPsI44JKRfIhSJjoZZ51ZcDanF9TtkyRuANRZTg+
pxoXig1jSj3xnd20dyC3D61qw2vQoUHIV1TkeUczqd4vumLrJ0m9sBkaBWbEZUfGaL4hMdmLnKR6
+UfJ439U0P6xKbRNjveb/8nde6OFAPhTwFCJVnF6XpV605U57hVV5CDRlJ9lASAiJ0xcaQc/wtRa
E4uJMcP3y3VFOaxNKfJdi3VKz3q0l7g9NoyWZWVZtaqAC6sX48deoV0MTw6q8sPuTvZia90W1qyG
yCBD4WWqFq8mxf5EXqm9k/htcM5WWgLF++S2vUPI8+0g8cufk0iSwp10z/3RVjp1x6rZYtT5vt4I
BfB4XOXYAJdyyTS7h9VQXqUBu0a/s3ZR3DrZHoe+CMDHRljQtV1p6TM6UEmLt91jAnjkz/0fEK5F
TbwI4P/xqz5IEnr85IADME2saCuQf9xcZQGowFD5RsivZiCgERJNitrWacIsevqZlJYnp+A3AS5k
yrJUZcj1G0Xek+vzcBLvslWiaNNU/Jy+H6Z7vhzSCzY+wj6uly3XqyI2uNPHI8Dno+8Z/o9SgQLn
kCXwKxab2LTVv8FaDG6Aj66eRu4aRXXuFtKlVQUMxrirIlEKXdH6ntrt134+DovGTDk6qQGYkp0+
hAkQ9JlEUpqKGEAMpjZ12R7bTP+43D8PnI41rWWrAeHe8QzmNeE/Pki4U2s4RYJwzEMfxKRukYQ2
jx09G6nDU0VG3Xs0zqVE6UvnF+IvJiuRbICZVO4rCBvDB5wszgs62XQrBYje5ofpnzBujmX5UgiJ
m3FMigDqd0N/gqBXltSb0Y4VAcHmujTmxTQXVgsbXaJvyTSPmdFvcp7L8HOP7n0QR0bMoTStjQyi
C06TsXW6tL3j4ojyGQdKXQSmrmQafcNztwNa58R8KIeFmrTIoreHo3OPBWfxLFqL2dPFPJ8g6okH
f1Wh9sLt6ZGzvSFJiP/nNsv//ZpPid07s0asmlp6GJHEKukOfvjYiuB9nszyHgpblgzIs80V+b3n
L2W6co2m62qEgo9gRSHrDMQRw2SOlDa513zKaR/2A3uQEBFQIAiDHZtzYBAIrKG5beg+z99Q+zNI
/kFhcfcI/QC6LlQqVh/NAct9GUAlX+iUIkPnoSeMryxmA0MESFrXU0xbsqVQbK9ti2uT33Y2ySdS
RRdpZzPgQRf3pwbZOcnFfBrK1iEfFb5VP/uLLK0EDleuiN8tJRpEhZMpWnLHH6HFLUJzdsClfEwY
IcKEnf4UhUHQr1PZRlxIrPQ5qhoPMSOxVU9iOW4m2bw2WOiL0Qs60gm8pWfD62+ntLnsG81vrc9x
SZc4kg9T2OkjsgE/wQ9CFKeU8MRviQgANtFwQYhTdaDXqHfPYarKvcnWOHbTQWx1RG+TeoNUE10t
hUd6gMjn4qpVWQlqbkwHNpcG1l3ZN94lje9pPlxLTycdfgu0IKd2mvErOuNqDpbS4ILirm0uKVJx
TDxiKcu57+z2j7556iQisK57nx45409Yh9+pfNiLZWy65u0bRl3a3avt0czSkaW8ez+JmYUF14B5
1L0sXpBKBvCxJGDD+OXutnYtxwam4PShMuxxQd72srWc31+X4s+UjrlQrdBmZzFxYhDRuS3qN+4A
0x3skqStOVXwDzP5RENK93eMhGVqQK1VXHiq74obFPiQja/dR47vRDx0FOgTIP8kZT2UBg2MLW6F
1hRJieGXwnLJSVEpdS7pgFyzGaB9SeaGRvRkzHifpse80k//qcbhsfY1xl+6REaW7YHFhMibLWoC
vz94In/aw2+dqoKmd9pikijxyI8GlO2fVMLdChVbxLYvF4jB7tVpjIrajBOPWGDvMpBI9R6THRk0
Jr5TfdRqkBn3uZMTJF6ioIrehlG8sAVyVmuAw4SW8pahZsGFCfSy/J8lur9xlDwtAPh8Zv7C7lrr
I/kq4hd3jBVBEN/iDdpwVLxJHOzUS/FZYE7gxB2yC8taza1q9QkACQBypKzwSeCWLfvZA7XgqNDo
wtgsCnw0S9AQh9VHYNMwBt/S2OZ6Mraq13Ck00ix4LKzBwjHLPMMwn+NgcA26YTD1lubBFo3LFEu
JL2D2IcYO9xS5Cd2FCLJjRVmoIHFNObxVBOEkRcgVlY22GLg7gR0mHxwNdpFyCYXYvNZZ/ujz1it
XDiMoqy2wiRb/e608RIiHNbkq3Q6znQziNSGFsEvf1EbndMxX64nH0HJmfdO+GJ18bQP+UrukwHw
Ranu7Y3CaCS6nrz5J8d+RVwe4GkpJRtvJmcjV0q4J+ooafR9HxR5Mt1ziZn+Q2lu594612FQxb7E
GsGZXf629YdP5kTAr1Guy4k/7Ke9C2KkN7lFxbw8bP5IVLj0p8NVvkM6ecTR/x43coJaOn5lHluy
os3i7yEwtdZtIcYZsegoOC7/7eYqOsRON+e4OhZuLY5qvpW8gfPKHozeOSLTjnqzeOQk0luhL8RR
SPg5PLsK8k6W/wuTmRfqvj7rntjr0dwLjdGqLWAXC2SSAetrGvPwfytbvVQt8QMiQO1YS9Iv9arX
vE6RElIK9gWQetGW50OZ4S682rRyUm4KX8QwYij2ylraV1O5W+Bl+KZIh/Dy2g2r5fTWPfjAHi8r
ZNNU0DfmDpu1RRgPzb+Gxs52rhIvfk9LXk4ZhSJ9qSkvWzINEeUX7of3vEY8++xo7y7qzxmECp6i
vgA/uGQd3jt3BggecJrTK5DbN6vSLDOsQUuwwZqSXqEfH7xzFP30efhHxeb1VQJ1T0/XkJWatZaW
M615+RWE7W6QnKTHuYDGC0PrBWRbZVFK7lFoUPd4npLMWaFuqoS8+wBTUIO7cma5Nhms5cUH7Qz7
xMIeS/hU+uGeBg7x6sk/fB1qn3hXqpVxO6k7u+R2Y994BK27VkaPGmx9mf0wOvP05Ziy1dxCYdXn
iiUc6trT2E7zhlujNnaSGF+ONwvbOkiR89krgESfSxjNnY9Y1ACEuEcHSbTUtVgau0ldnIsbhIed
1Bqart4tywd8+uLBHnBSkxRtn8UjXiZc0+Pno/NBgy7TKin+F9OQpP8WqwxeIrCeuybe+ELqo0RI
YYNqbuGhXMOb9wpEHTDa3wcJwAhdkZANZQyTdrQR8Z9gunWqD6R9Mf/XGxt0JsOkTtuKipXvn4GO
YGUTmB73J3sfGKxIzmxT+eiOyCnVoTON+43d3psxcE4JvwUuqIm9UStwV+xgsKovQBhp3bjtxAU+
/61GgkSVFzVHWP4ISecBqtCLx+kqdPlj/WjAfqeYPBG1V60H6PEbmqfp8/Aag1wupq6DC1oOIKwr
XzjzRAxS770MNvrrqQRgX/S4K4LZAFT2+wIx1gKiB1C/AX5zFkDhuAQ5F0tiwbiveoshiYtqHPn7
wNMYKEy128zunHjRb9Opum2lW9zhRKJM343H7OU6sZ2/XNCHGMvVA/2MJFwMYMoBj+Tem+WWPUIe
3X4wHd4BpHbCCDjLq/uZzYzcOWh4zc9pAhCTweqJJ1I4cBO3OY5ZP6jIzDsfpjs4nvCHm8TBfMGW
kfAek29B/pPQVcJPv1TonMLn/6UVNE98ybd2buuP/ecfyCkjGW1CKhIk2gsEfKaiT1y+L1ZsF6GM
+ddJkrAWZH0FLneZZViyv807U9ForWgygtL4Q76RqKUdeDqUjyBk3ixj0magkQHWoJhc+xO8y53Q
mBvJPVm8BJrM3lilxOxh/67fpL/Y3SNC4VCuZmgCVlKRDz31cjQjV4udlXABXesIXqVP4ssceHZO
dtzB14OVW8uuH74ufYOXJVlghRmkoJX8oju1H2Dwp2nqjkB4QGNzwz03TNKKblJt8u/WbJbq5HT+
SMlv8edwFdoNNq1M7YiGhOzjfg9juC9/H+J0OLnwFZ2dhHR9bOXy9LpnJOMoB2pUlgqHHneA3U9N
Ca4PEss/XwcWWLx3/FSSzfGFdnXLhR3gbDvEGjEtQoU1W9lg+wSa/mKerBuFVKUGOrWkZCj2Po70
DsqQUIcL9P+rBsFrrkcPvq/a95KnGoX0DWkBNkLA8OhNc1gF7IknzAuSlwjd0VjK00rLwkhaEdWw
ZAGUJ/hTYLXsnoBxPbg97NI7WfhYbFOPObp92QJ9u3Hy/GUsMZRYfQQzjbxnNlB92z00KV0aZta+
JbzrGn2ig/131wYN7F6hbw9/VCzNLJJ1UAyejg5ooxi327CoMF+PhjefIBCD/+7Nr8iUOWgOpJXo
3Y2uHJMLJgzWGwgh6ZoV2FQKEhY4y1Gxx+KLgExUGhZpfpvcjUgsmqCY/4pr73vQSMKTnyVeXjup
yLAmv7c2VfFGkQufriEFCEt9uGG2UwstOPp03GkptRfnB/e9xsjP+SNfBg0PO/vc8fID5/p+xHrr
vfthlsuqNKUivXt/CV/T1EjmX7t4VX1Fj4XKYDNe3cx0QsPZHw08C9ND0/3HGcE3oP/G8v0+F+Ld
rQFapg7GvtRysQ3OeAO1/+HPGf4u+mAtYQfg7KjxeSY1nj3z01PEMZp26F73/T9pGDAKOzdTnLEl
83vEz9p12+cB63im+knLpT14C7DubIV8CQ2xT/y+6XQTFeCqC9bigawu+0hByrQrq37tE3STAEYc
LZvqcOn5nKpDalrPgqC8solbozRDIrIaUsX9xC1e3cvMwMzX/qTz7MvWvEGS6I8Hgt27lYYuGqqf
yjXs82uzdjhXa+sIZR5VV6xNlMuX+AVgMGA0eWGZC5MdcRbgN293+8/N7cz5PaKXb8HNxK0xBNxT
vcZuRQwxMyJGSUvr+CEjWDfcEWzTRhPDCU5FLgGdU5bDKOwfrgTT0pa2IMBy5flRFdBnLXhr+d9f
AUHaoSaNMsjVt8iiiKccoU9lQUFfMT4nI0F3V9oYktZCBk6hciUZUpQxpC1WjMkkogEg7pdwsXqL
St8/2D3Xs1LfhssmHO9EHBfKZ6FbOSWnI2P7mQ47ptqp1/2kxvxW1rlWH9AB5cYED7u4nYEnA5//
FW3pPwY4c7z8uoMJGR/HhKSger19sUbbSFqzjweUPTvSbfrBIj8kdgcGR00+z2hwy7kHXNZ5Ei3y
87DlX3rumnYPEY/QS8B/imwFsElhBzN3lMRLrBQ/NCDgGLzc1q7ydh30LUgrO2n8z41/9h0OQ/0H
/cg1f/Z7OBnAvIEIdQP60UCxZVo4az5nHf+Ad0IixPEow6oz/HVK5E1PireVcsE5ZHSCx3sKHR1K
sT60qJ+jNVFdqnQh9jg7+0FZF7/m/Rjli/OdN3bUMJvps4aBps3iYHSNufXMMaQggxtFSRdKz8YR
m7Tb5gto9aTvaeHWtdMm7seuXFh6JZfERUDxSzmt7EUuCNkUU+qFsS+1Mq2BamFlrGHsDRDil/Rz
EPqDmml3PZYiGea2aLLyP538/yELsn9LDzBtzSi3A80fNIVWhbUxp9MQicoyp1EKio9G6HeOugoD
4RaavOhxrVID9m2SydkirqhZ16wTboLsUFX0hNnP4vU9LW/r/bzB5zxeR9VCoGOTrEQW0T6siq/V
q4FapqVPOYqQgyRd8FhFehpumj8AWG7NuQsLH+GItilk9Sizdto10UMHdLIH1fIQC8pdJU16vX9d
GotblHF1//Hn03xR3JX5sv4CsYRrkYqZbwGueodUGOQpztFw+agJPJCuY8m58ycYoEUdxPfJlBJe
lFVgQxze0Es5ekkKRLvzt4OIh9s/d1VZRY/DFVHjD8xO75bfTLcloXCu9svGD3gq25r0T3NYEa91
ZeoK5HpgfTr1C+jXfzQ+f4ahuM/3njhrHR0uVR3p/231azhS80yNh7CG62uXN9Xd4VCL8vceh0C7
VSBUQFVSPKS1dzC4y3eIzoTpAjAskUActEsV6nwbSW8dYyaFPvt+Tc3aN8DsH+lB2AjvqkQmZKbU
778fFR9+EAAbNepHh126Quyhbryo/ttAlcDrxl6hUD8of75Mw76yujsd2oCYL0DLI/0ZxyUezUru
k9ytgw1nFV89l32cGK5nfwqNTOP6WQu1Q/C6ZcExZlvJhEk6qhvDyoJJGxRvR7O5OLS+i+jk+iUl
J8atM39c3AwrIMMMTzW8me9oc+6b5ka3bvhcQDRfLdrPbI/mvTVpBb3DDQjCE6sxd/N9homG3Eup
xV2974gLqeBxJvqkneRZyP8cV4nFcDK/ELu2lZUvK4yUckTRDJWON1o7Bt/ggZGUR3hbaKyKOzjB
sfQkB72fWF2DeuQe+VpS0xJd7sPbtpRoLikw7CDBK5jQak4xQ6zyeVZxzGzTx/u5ddC2B92hj1rB
CXAIR71UG+tPVh3WtHfx4udWGoPUhN9yeAZtH5RwgYbLRcaN4G0arGmSeFJfQkqy6inNsslc5fET
CKAlwPap1njWFcUn0n7W+LLPg1lmcb6WPm3/UlhwMUsLLYv1szp10FyVMzULwDcpOeokMAsmHRHe
uL/J2VjkxHdH/u8Fra0ut65IyabTbmYOfy17Udy1STktDDkbYxwhOnJnolGcL+1/FFfOwnTR51Wi
/sFAcVOcRf9GRI9JJpgD+hO7JdfvrG1Zi/YYofG8GYBqit0LNFizNvQoRzEW8XynrUgRJtlmSc9J
j85Oxfm57uoG7OmVCjLq5B/M0KqNptXxmhevoWU/bRJrsS+owbOZ6t3A0w1jCJGu5Qd/LxO0stD6
KCnNrOgBE1Ut9D6G+10s21yab5IKo/+hau2GDJ+Z+Uvg0S5JLLOLbrp00HNL/sZ01aX+v9tZlKil
4qTZjYs3DGpzsGZhYHAg58uErfbhrE1io7hUM3Scq6Y3znnmMJwY71nPzrDv5cXDJnhv/dS6Ai0M
xMw9lKU2Zr7Ft2zsUlMSrOMPaIy8/b1TWiCvhK/NG/oKPtJGCgO8kpUiw6NP5ve/KtUtAlo4Tcry
q8IwK26C0oSXB3bmjmqCuDzlY7/LzrXtuaQK7PcK8UXw/mhas8YmT6UKj32s9LNlTB85zO3OnQyv
ui5ktvoUrmH1W0EQGl7ICIJOmVxnjbx5+EV7HmNtzVayn8zbawoqV0dpBapC0Hon0YmZbnmVobwl
L4Xt0lbSS7VGZJT8cYC51gxkVV7PpeEIwzDPdO+c9w70Opd/9As8oH5DH5obP16/kEzNo0+PTPXN
J6ibZ+c5YX7hjmwbLgqBouHUFw9XLxBCTt5wtY/x1+2Lh0J2OxcN2MG302TiLJXF9ml2ablrON+D
kSX9D+QwpsO1mtg3yGbPhz/fBNzHe3fsacnlGef/1c7Y1KA+ZkLlnUI2J243kz8IFjOBWEvoO3OU
D+7M51wBE5Nx9m6+ORLxlmL+JKdBvx3fjm17QErXKbeSo3BDd0Pwext3af6py6xREQj+tq3HS20D
xtNBbPQFIRX5zZvdgcBJVH3ke7oKIG5nWO9LDQZHPdLY7P7YYo+IIR9RnqOJIYvltGxdKxUlmY80
yNP31LaeavRquHKO9/HP9QZt2JDR1nin6oEUjMB2P7l3TjkvaxDyqeBhYiMnCTM8d2WyE8nOJ+up
S5vF/0zN/VDCWsKBEpDBD38KAwfpiCa15BYC61HJReVwGUshaIBRLYlfXCPd/NCsTVgJaqAMDiF8
pQNE9121tVXiInlEOUeYcfwIhAP7VBSKcw/gDySl44v1BVzAy4p7FIrOjIf/K8sqamhX3FMxzuWE
L4+19cp3LJAlCLuS8hhzHxu0jv+MptxjiyOaPcuAwfMXDo/fEQy3lFbr3nvOfh8RHmsihUjNhPCX
ytHWQVqc3WVyWYceyy8GLJ/JiRrJfwn1ZJlwEEnjVxSip1zm2YIbf9MRrdUxloV2T67IGxZJJJ2k
TM9I2NWfx1VBzic0GPqs0bF6tm1cXPhHMJANkQ8wpx6YExmNtPgrfFIITFSX0y8c8McJFC51PuPk
o+a77akqSGKnsz4XhrcXra+qMw5Xe8iu7x7WKKjbY91j4iEYN1Ns3j5uaFFDsKwwjB3AhZYrujh6
h7+KkyaSOToW+NACkHihCGRMNBj953VqgpLcFNng2luvYnb3FsfG4D071ij12uba9XiSr6/t/Xw+
yw0+3CTBXPTh3VeN5S+uI8mHyTcvzhIRn6uW944GHGY+uipk9bcUyO5+Hk9Np1dptKZhoFKbvKWR
4v+qP0l+5eiFQImINtecns9PvwZ5FvtDsGd0fhdG4CyxXiVq+6iE/x3Ym9FSlGUjLKE87bnEEN87
S3OaVwbp1VXhgLzjHbeVk5XJzNGXNujGtyn7pCwHMbv5GSUztnVF3hTje721xk4GyzS3CMD+nH5w
y5bM8UfmvemQgVTVAVqs+Snt9jMEF/REqcxZg4MCXakQL9amy6kqlPDRXnaVIAuX+CWdNbmd0mU1
0bngy9baprUmYKfdYxAlA4lEZhcgnkr+tceWWjitIon4f+YoESme0FcB6T8tTf86mK61n7OR/BPp
S9YNIEwYsAapBSnWWT9HKBUhN7RHOdMjNXBagbrhYOpqGDcdls2GLNWF4EPrNFgIbpzUUsx+6ce0
8mF5qtfah9PnCO6tXiLSLzaDKdW/Ii+CQBPeliPSMFa1eYtI1A6KEMwZCzrN3nw5PQ/Z5T2EIa+c
suVf6jBXGeSM60khN9gzJ2khYhHQ9AAcpBqizBUvxEPYx6aJ21nXF9OHSIqumJ3+fyRqdJEqDMYN
6lTE2suJdQeB+MK3O0FEKe2JazNcffFpxy4b8JNwZ69JEPlLPdgH2xz2Vdb+2XkKbUNcVrVeJT0B
XwiMihoy81VdA03LFW7pLopjcFd8U+yuD5GQW2cLAoL3VdG/3DPv0HANwqmfs+JrG6SP/6hkUR9h
EThimtYUljIoD1TXNaMR1e4VUCC9m7EjO7nD2Envcztj3wyNF1wWIV8CbtdIJOjeujQJQSNZeN6L
0MOZuG/gDFT6Wbl/VrhxjnVl/8d6M1NW60eBtzmUB3uL3XGPbK/579zWnXLerb7ZbaaG8wwXx31z
EglWu3xG3+TE9xqFcjTITEDOwn6jSF4NNlcKNplaFlbloegykBHwQa40QLDdU3rMMLxJRPkers4+
Qdgc9GT3qgdnVi46h9gQVLV2l9UJ8XHEESjJl10sRPzvZF0/q/kEqaOnJJEYxUOnfhlOziOsn07W
fWR2ZkKLwg93oqbwLUB3L4B3cb6P1yQBYJYFUCAdLsCYko1Wej4mdu/72YCZaRQhK8OhdM/mhsBv
PywO5SxYs0pKE8/uCp7yvg90ZkISS6ymrtpFgzbrexHmb2JrC1yIBhbVubv7xAePjPERi1inGRvs
nifraBCRE5KHaenHt5+fMWJwwVad3ps1PgxxRBSpMPnOTtvTPh7blrENbNsiZrPV1VDZhgLGQYyc
ba/IyINVPlg9aGbg62zHPPiMbZfTH6F14400BBs1uVcbpopW/HVPUxwrRxzOaVxFqJwfxhufhO5P
AXxj1CHll+OpXv9lKMiC2goaQGd1mM2tFsvrkEs1GCF5ABsZJ4K1tHTlOaymGxMtKSFyaLwyYQmU
EzjTUCZarzIxS7ZyYw7SVG1ppFAzb138/AjVvjkcAoi8tUPwUdDnn7ULiSSGY2fHP4GKaz4hHGnA
mcs6kAcPclzAy+fmnvUp8mJGXnrVv6qMz0KMRewMrEi/kOZq9dUUqP5A7WzZ4J3LCbhgYn+3BgZd
xKLz8JO+Cn2g3a5F8f+vmlC0PYftNFk/Rgwu2a0lpHHYIRoMszgIfvldz03rgesDzkg4YdxZIeP+
JMlInI0yunaCGIJLQQgOGktW7DsUPLRB86DdPvv5bN51TGZmlGJWB8r30Y9U35pxhvrbb0KeHb1+
20zqAPpxSFdfHU0NNt73hpX9WJmV6JW8WP1ErtOb+/yNTLI5j1fN9tTVSiN1Cw7a7KMtw5rtPKT8
Rhmza1fJdiMYIaIt9OoQk2sZClQfu8sG5H1sVWUYF8fHgZmsCfHhLH6jA1TS2MxUVPtebm/uWxuB
RglwXowineVGmGK619FuXFxutXhhPhgxVm5In05LSnfgmajCFAsHb+HRtl2SivYE8tjPlFIz6+OX
zZ3jKGQZo1CJBMHdbDD6SaHYVU0Oherfhz/7c+3aX4kT2IzGxBbaIguE8JARHlVohVT/gr/+bcY7
BSfpgYLwUTs2ZPiNwnUCljLowLsMt+XJsmmd/ekX8GRQV7Yum3RKWIF2gJsXkasCVZ+ngppdn3S0
5/MLyfLjOAxDQf4Rx/2J3CfB/IH03y6mNq1+j84DJEg4QqwhiwJTn0cAJ8la+S9LPn6AYzmKvju+
977UwpLm3+IWiTaFf6Fwm9lmp89R1udiU2vxNxpgaakcP7hzhaYEypl/TKOV7eYVQoRhfW8GVvzL
604vNNDZejmWxrpX+fxGaK32p+x+FXNx8SB8RTEA81b3BSls1bZoxRJt4mTTpzvoLzzjyDMZCcVP
r7kuMUCR8u4B1fN+t8yeVMRcotAQElmBbgkAZG9XPaPCrzJWoolXw/twJVOpcIJIS3gW67+8VHVs
9Hz5QLQEicrYSeUDwC3JeuJPq+kGwOiIC42IfChJNByj46iDAXQFoBbwX4S6a0rbucPQb/LtlKgP
oLi4gl38k6aoYHR/zlrzgR8J02aICtNV2pyA9XIBBiQ1VtuCY3FDpUhS5STpOl9Cz0PSwTkwN0rm
yfAZEuRiy/HnecF7yYXwW8rKkhB72Ww+Dui0PebMH0yoKp2D5URKBEwBJe+8jTlAE7JIZ3qC3DIS
pjx0KSwzSTQnSyfdAImznVvOS0XCvXr5JIZRn1D5MmF8couQN9eCt4y9IAIuyyDVKFP1t0iOpYsE
Dwla76jFOlZj+vQj8EPFMmii0ePEiXZ4MRi8Ae1P1BVRZf3OLC9FuHAwx0L1uUg2u98ZHhFCI3uN
VkrxIAnxyLLLctho/it9MCmdMdIl0+GDI/d/12D/1Fj8dOivNMOwjUYsHKycp3y0q7k9eG5oo7o/
iRmI6j8IESkBBk8rhMjfDq0Rq5YblXwMc78R4gcydnjgpikv6CpCZKpgaoj7uJxjXaQOyNCDcIvD
k8U52X5M+bSGFmbdMm5v5xy/mfIZiJa6TtJvilPTeB0rtQ2dxA4NJqftJOS6JgfE0exkZLCRU+Rf
BH5GcNHSIDcPhFvAUQISF6MN1Ud0hrI7tvpijIP1Tc5OuucXLup8FwKb92WZAmKHKL8B4RjlQ+wv
2JGuee8nIkKLmW1/kXRY0gpCRkJetJXtjAjWEJezMadfU01c7sxnLLlwpPIHUwl1aaqq1HwTDi7U
nvazfqRBcvGxbcZ3MxIN62eRhbagLvqTA3VQ9c+4CPvF1GA0gQ5GmdhCSs3NfwnPlrg1ceVAKsGx
MooBdA2Bw31q7RVkFRQY5FfgsezdGt5EAmFo5cSi9MXwkxTtlqmmfjKsslVhkKtiI1WPzfj5G9CZ
kxoxxSZJ5IhBbLxlo20jKBj3sCQW0DKn6Ib7NRzzCbhEKrOkS0lbe325n7xhrI/eCLuYr6KlywbJ
LfjJmNsmHUS7FthjEHCFvi92ACkUWLIQ1hPDQzEHgVvG5Wm8q5IwtSnNNFys+7zJALxjH+3vB5XU
5QNMXZtIYhTX68SmQH0/ytql3amvCeJWQXVkmBpMZhyQ4mdm4Gra7IQ3RXln2izNFXjXRoo6bJcR
CuGk8T9og4ezOkhYvYHhr8UInoKLz8gpacd3a4+N5opXoBcO+FLhRAGz7wnVi/NOIt4CiYW/w4zF
l5maarwRB+aHpTnaFY82JDGmSHZn91w01JKraWukQlIaR8VWoq9rhE0mM4jk/9BkfO7sRM15UsEG
WEb0PbUidQRO9YiyYjzTrHfPqM+AbcXAHImyxUnXRklCQfF+s3ASXAPRjxcCiAImYbkqFb78aXQQ
4s7qyMJEtafHynvlP+lbJ2A+/ku/lfEaz6g1Eyv01ncOYoLUJGh/uAn0bvZVsC6yUlyuy6qfMJJg
om9YECqwTIRWvJO0ftB5+P2rbrNMZeEk1YVpV9z0zbfB3hFHozKpF18UGelDhGwHEr/VEqB/QAsh
6U1lOZsToojlL2W8m5uuQqnyE5nHC8FSSXbHvzp8Zlc7X5dM2Gt71g9Xk0Sd8SIbJzdIcGUHdKW5
6f8deyh63fKDggzI951wSsj4hn0lPTdssi5QRio+PjzQqTCDINNTiVY3HNCrVoXwC2MGtu4rrQKW
SIgOL9PGj2JyWpBHlO6Bw/MLOJuq3PU9ZJkvOwYctGI2FZ6mxx9j8KNYVJB9Wbp1uToe+3kbix7f
xX+QFrYlkpyH4K8yx/0MfFBlYY+LrVj5KVQ0rLfVxMOApHcPlxdauKteMjwX4Z8Slplb6+e70OmR
Mf9SQrOlIAXTanwdFz4TdRsF+mC9MDQM5WdPnJ3vnt848HQEQm0PrI4iSUcjRv8AolkGBI5D93k/
rSHRgN5IaS8eynKhPpmQxUJftaiRU4hM0gVHno3wJOpWRuoTu5E3f1ndb6jME7gpG4+R5+Yfe6Pd
FkqBm2iu7yZyg0YHqHxAp+snqaoMuzk/bPa1XF5DQrfgZ6nU13KiPb2+R9IPWD2mLITWn3ALDHZH
ZZmP0XWqVUnv53IPPylQIdZIDmv9Ehb56AlYN2WUlN7Trrm0ztWS7Wa0WuoCNhxRP1N8JeigYjjf
kDm2fa3GRtS6cFEpg4VZYnBmDgyO9E10ODPXrzoyBnGkygp3uhKxjKwtCiEnms5CKyMKKh/plXyX
Lb4f02I6heS3uJ9r2G7/t8Sfhd2ozmAe8vO99KgNA1SPySGg45VRdOiKtAe68T0w0K30RyOlJ7Oj
A0sgz+gbDTujUvbxHiEuWYB+nO68G8s33O1DtWMIZsxeC6yV9BeJ3t+qdRYm/CafNjgyJ3Z/ZW1H
Vr0vU8A0SV9FcucWOKQCRz99lBlwOvSmF/H6DuX54sBT2B6n8qwp+qyGW6cVlKdy9WTEiWfh/6cd
KbuE8VC6B297p0B1lDVWruXeyYlPdO0kIwUHA6zhwDjexlAOWH513z+vloLq0qRHX1K0dOUFpCGn
27Fe6RZWbJ1GyOzpvV3RnJNnEacr9NL1uwlCBGgZuerADLjQp5a9Qxnqz63v+01ZjK02udcu9k46
6hKfUSBCkliujFooDINn0uPyfTDfvCwkk51FW6ZgWGNOLRCSp+Cgg5MpeGOkBrdeH7BCxm98wstT
5Ts4zH9YjCoMhRQVBhSiiJJUsn3DUYy0UHx4v/rl/DrZpEp/byYlVJv1PePfo465m5i2UKv2y9nr
5db2mjj7+3rDR3xbqCue2klT10W6oMuHyqLeXdZCBMmSkInp0ZU2pNDiVht8w79Lj8Gn/wghLTkx
WeO6RhDd1jRcWP2TlIidsPXqXbRuAmLFh95IdrdIDfgdvge1l4OFDn2ElvjwUIV+Wszh6v0+rITa
aLgdBO2+l4KJp7tnFoY2CNJklJ0HUFGcc9oBSIPuBg3IXr+cyRU6Y7yGpJuo/WlMuLu7Kx3k8xiK
z2AT+6HMkE5Doj7xoqEyI2UyHlgfnwv1TuqXggqGw9JlEstKEGzEaOCqnuqMVPSPL0SbsAWNb23R
9syM3s2IKqkjSLRXvXTrSVadCgYuqE3k4gvPbPF7JTPOivuoZs3i9PMcheJjDmnpbiUceEP7ITPN
9TxniD1sG+UwzaHsE6JVIsSQENE9PT4xK7csW3Hfh4RWJcQy1T+keNxq4IKQudrUeb5HJKgoUBdo
o6iMC0VheUD1PEnmg3eyfK446hFFJKvDn57gq2cxSi6okKbP9xZ0NJXbS1EdYoLEfLbW0TPr2jNY
ADu/4W+UmxPUyhAMOHj3EANNc8tA48WpTNKNb3KDeJp308KSRTt8NkXk3sLFI6V8zvGmPyGRv9x1
gst3YRPvvcMXBRvxJgY5jw13/BQcERsScwclDbdVUZ1G29vqZCTfC72U243h7y1qwKsMpVPvbOW+
W6R57cW4hNys/3lLtzUfr2NqEb8Vb86aypxxuv6+c+oRY5/D9umhnPqovr507sbnw3U4twjmmItx
OLJC8slmvB15bd/ZHHs2etshbxsWvhv3hG3T3EHqdJUWv721yUHtnFSElJeHwLRlYuDRmV0vIk9h
CqPvQdWmOHVPlXX8elQpub2BTbCyFkZUY0wMH+CrHGlDCy4Aw3dLSLOlvuQWcRb3dkZD2c7j+5ni
JgqSNvSSE5k3SB+Bc1dUCBFmijwkAxkreY3QCHNCu1/iKnfZ3+IwDOgUOGvqz8n+lAEEcSUTuTEy
qBPsLj0vX9kEtAlgKFP0wcqS6sLOpaXpshGDYDHM2ErxxwvZCN8VzWr0bMAvbk469Nmzj4K+9uhj
j8E8SvZBlLivjEyTb6HBTp+2W45p0zQFBc1Bbkx61x1llawcz9yd0FUNmJcKgjZzsLM0r2nXLU4N
aW/97b0qOO6Ct9RyMD2zK+I2TLehOXCyXzhWMSBzB543g/YWbK8WAzC+FbKuLMOLwXh7MvBEr9kB
lKSGg52EBlfV4yKZD68cPR11vb8Zf7/rsm1PvJWheys/czVKffKKZW81/BP/1uREJKpp2YGGDkbm
qHhpIRsjTyhxBmp4DanCM5wND3l4zxEfRHMTWWyqILLQtAB1VI78XO6TGd234W+gcKEEbWysb0Md
lYwBHtGkuOn0AINjADzc2tEwyLGd5llXi9PyLdEGQ93+5ovw90Hp49PEyLB/EGlgkxOS6UwnZykO
jMiOqcR0U0Ji4Yho6x3HNzOL9IFpdL/IzilUEjWnreQeot9akm/INIWpoZY+9WSCoNtvmQXqJZpZ
dteEANgJrSdnm2U2KtcK5HDu8MTwJKTeqK9sBsB9/Ec9cW4KJu84uD7Ac2jRvO7hzzRlihM2ENKi
dy/QfCDFBtXbYC0q6KW/Ytu+P1I72WQpCEi+IYxr64yk1XawKMjhDUqrqviycu4c9RALImGehiFd
XinwHmBQWD0ocMPrs35hZmjyCqtOE4XQ/b8SUs9Be+3zB87/WD4FsBKMoLQpnS7Y+ZUPaCXxfEWS
B/jTWiZDDl67V8TSHpkH6KTF7eo9Zr2gGdMskA07to6GyYAgXNYdT7nIULYJ7rkEYWRDohIN0mEH
0CfXXjCgiutCq3HoAQ6Y8JuQrvQhmabbjChEyhSjBHxBJUFBVy8E7IGJ2vd30owLXmERLWtBStbk
uSaZUQur8eQkC/nntBmzF8zkD4jhPXVc9RXy2I4lRGsQOrquGXz6Ihm+HneYzw2QW0+Yx6TCJ+Nw
JPU3q8EHN6qAuNmy+m+H/Z4xz4s140V3CrEhpky4lV6VAYDF4hYZZ5SCjuYAfoteFRiRDDzIlfNU
4orUacpqU0fIFMma5tWflpB5XqCXIpt/xlSXCiUYr8RpYq7eHgdaXvX+lwMo2rHOHxrbQn6JQw7K
Bol4D2XfmrpCaI68po8dxVMZ5MYTEyIMa8I6HqOzoSThwpikJ7ZX5MvofdvshDtBRXd4tX8xhugn
oo9koT8Pdg8nmVYSDzFG3N1um47Ct2+KTlMmnhayA/GnjJNY83UKK+FdBkA10WmthYBXEBX4jusz
3u+2f6TZZ1f3jqq4D1V0p+j46JJWY2hYIwpLekmnfJ6To6pU4Ko/yYqP1jbcUkB9Be+6s9T2L4/x
26rdlB5qa9WCmA6NQ9H7RmTD3ri5ath7qGRquMrF5slHRrmYgkOk6gj+6HEQu4uUgbA65rgP2WZc
Tjm1eB+DuCqVzBK4/xx5bNi8zWsALhYMwudjbQuH0MgnhlpEjS2nECWAMx22ZuYBRfRLWdvheBjZ
ecG/s2tNsKs3FoAt6jwRIcaUanMSsZqiSHl9LHbW7fOf6IHCDuzfKra7qU6etCBis/48vTRejsN1
n4wCPAKPEFiKBR//lzlinfwaTXXIj9pgpdMGZjR2mXvcRTjJwk9odIKCMI6d0nlW+3MNb3HGBXdx
h2wDMqDm4wKZD47/OaDicpovMo69FIXOwYQFAj5t+qlg2ABMGr0Vp/dy3KVYKeyx1beX/zPVKgb0
3bKE3c+OQONQPQEbSBsxma5SWxRmhDDqxadF9nE1jKkqLTLre3lKnEy/xFGwo8ZsSTwhgN/UGQR7
yS7/ysugjnlc+q9qnbcS000MJLlrue/JyBjHhK1xW87/OGQoOvv7toNrr6/t7y19SudnfEMyYNXm
O1EUN57quODu8G00xnncDQeHxpvA9MGNHy8Qjbh8MzzgZQP9GtJaKSPY0eK5zKLO1XEZfOV+NNoV
xeCfpWJ4YcLvKVGqutD8fN1CVREtoCarYkSKVzUzkPCF7k0vOgxxjBz/98Kpaz4zeDrQ7hOY7FHP
qUoPt4y83dE0j4Li4otcxug1ySyeVnRbhTLNsFl0v1wEeeaTimiurJ5WH9boYWM+CKX1vOlSYMxm
D2opqVspfbInOl4U8655zlBSlFib0ZwlQ6erE+kTecaaFTwP8iEIIxQ4y08ANg3ojAc9npPscnRw
41es2mZrUD21/sYyq8pg31IxJqND9SL8duwB27wr6MGcJha6rBEbN4drwaxlkjc8PA2VS0XNbnZd
HSG5ZmM1LSK+yPxozoQWNHH0jviVjPxGN2MEt0onGRPF8kOU2OHCAs4u3yx18zm7sOXg7iRYqCfl
VLKnKbPQJw6VojvgK+0EYOWPUwcXblxDQKTq3ZcGG69D7SjI45W8SrvWUvrGu8x81Bx3j8cIC+mg
tN5GTyX0tsNX+lzaKMbgq8q0WYv4Zs4oxu/BWtUIuCPV+etK1zRFTJGmPkeWmra7gVfalN5lxprX
R8afEET0x2pnLdLttMItutEixTmUR9K1l61fuL3fPEpBjicUKD6sRjYew90pAOZgkOa0YBWbBxc5
xPvr2idy7RWZIL4TvXA7rueQWOioDaYTbBTN6W+ts5xZLcnxJP3t38QTwpjTpwoHeUuIN63hsynf
+ANaH4Yk0H+hamgRmGXFKsRRBkTCID3NyvyJOqmtGz82dcZGxFJBGhvHr3qbx1NFh2bgilyDRby9
3GsLjMLMnPaDGgxwqgWWK7LiRLKFpzMUe4cfCy3JvJnv/PEofQTdEfoeQNaLj+ZK+rXak6TVfGV1
qYYh4lequ8PB0d5CFYezi9gcIdbaNxb1qAGmlA+PFVjgtiO8sic/Y58GP2euN24Fzl0args7C0IW
/RlftlW/UzXSEKCOxTFiAErT/6bj2+g/9N7ro1oTgqLicsaa5PK+BGR/0qhQ2ZTXggF9lrUdcIGe
hsyLNu1c8pBYmmkKwROZJfHGBi7VknHkeTwxkXj1X31busRRHE0FYYvK8berjQGvxDpbyrQqGUV+
cSI6ROUKC84OFyQMv3fKtmTdKYwP4J6FOvCi18tgVYKx/FFmcYYdMXmme6CWltrux13rs445AyQK
Qnj7s0/llgKjgDiXgqwxZgaOM4Pilnw+7Hi534vA0+LlCHNyewuAQzeFsVPAbeTb6Ce6NnrydH0c
Luuo1wMv6aRCmefvimBTVtbj01D2RNIqVVqLroWHJpnXrE9iao6vYsZf4yk+qqK5Sgpi7ScuRj95
vYgAABcZWA/Si6LbjLrOic4ImhdG2rFySGvBPjVYb5fQeMGga9zVXDmItTj7jYOWY0fSw2dVn3WX
JPhp8bcBklFsBv19L8P408k+YG21AW5pnK3IWqUUhPyJCVkWFUHlmMJEfsV/j7PTzTMptp8G0WJk
qfee74tOkXtlaYd8MRWU4a7SCGkK+7v4oB4kdm4n6Df5uv1Grox8SO0813WN3NTi8TmQcmQlvJtt
QdVrXIbiCZxsoDAKvPQBKu7IqYBXOtVruO5WQgEeGjxKuxthRM7i7+ZBIcdeQCZWTm6/Y96IgeLV
rifwazLUEbpkYjebR9yXW+QpGqVgcGJh4LBr3DMQz3B94C5g7Bh/Rcp745FTEfQRihTP0AYwhS1r
ea4SjhKy6UxZJtVgrEadlJmdyEJCDrkWwnYdcsquLE71Hst+cULmwS2GNs2KToWL/EgY2xSBVAMG
ZawrGJUk2tutwVr+ewzbtYTeBYUTQH8TO67+KTDWhwisakVMzsE/bHJ2PsCEF9XBZqsXEhN51adC
w3H4cFK7Ov9Ex6jG72w89NijjMkC8ahAHRq2zjZed/BzmqcJ2AsQEml++9qpQRTIUFBabSJXZSql
pwEYAECwVpmEWYG8wFsxSk9YnadAZ2DgZL7bAcwstYeXzVuRoYd2XcNqZthTIlKkTvLKk1wCGeOv
7u2Wqr4A62lqDzNApMPQoGHZb1lylZo+vVeYHosR/N+uXPtfPaZV3lXFgITmRTUhpO1K6LrDJ/KZ
S9hsWLMmv0ArYSM1Q6Tj+Qto9mJCK/yOGMZKpLWvWXbhnGDPIjEUb9dYiWvMSmmOuR7a6JdyZ1uL
UcmOLNbOZdodkA2wAECmWXLIQ5c6t1DCxtUelDHCTXu//3FVqydVQosaj5slLIRYI3lw6POmdL2u
S8pb8J9+K+clxwlqqfhP1mf9FgykMo54HEq7TvYylL3vdVSbdbtiiSYm5E3l4bkHnmk4kBtePaKF
4X2kSjWu11iEBFJN+tOM6W4fm3rt/5Wsai3E59/wrpwRblH+HrUvXVBe134fG9BeYhS/Hsvc2ewU
h6UpeNb2remIXUGeMLQIqGymnauU4nXzAMqWqMXWj4XoEFOOSudMbvbUDQUXMzM8vRA5WxfxSgsN
sqRxlZAQ2s6QreDPU3nai6JoSs3v4qm0XDgmbmRLUY/s7lpesCf8ZdHrFtNqlQMcyNwzu302y43+
7LtXvERVCWnuhhoCvmDIwQ/YXMZ0+Zq+TMw99bL2rm7fotHu9OgPFXK31JgNfhigiehZ8A4PlEjP
tdpRVuDqI/cq6HZLKwIsDroPHM/ZOp8nGA9b2iVGtTLUJdcPHL1oJsujO7b7AngB9ite/KKeUfqq
erJBqQhghmGoJAbvIpTl8WD+dvKS+NTwP1kogmN4KxGw+Vcl75wlEKt2cWfM3aHwDVCZja3v1E3l
NwgnTNYU2xeO7xRwQr6xbUynDDQMLL7j4DneBV/cExB57+Jvgra1DCUoIu4G/65YLdersyMuwymn
YyMUbgsENT+Y7Kg8R9Ha53Lx5GvUhiWZGOTwH2V4ZUF/P1mZAsTQkEaDbYmBBNm+BrveOYuZ1Ars
DODagQ4TUT1cXHr0jmKz+ufvtbGRoaq6B6YPV3ufZacoZOvIKtMmeCK2RXsHpktdLsUT+2A6qB8F
p1cvFTaBIgIkx0ZvPUCkjZDZ5QHltJIehlMgB3FQmuLkwKg0Psmn2IZxq+1z1kOMjQGPzfoImvKd
9ZN9Rj/v9NFEvXsNSPmrJskPlHDraR6WS5K0c0XtQSzFC1AXFjKWluV8+DUJoN52fTfnp5ntKAcr
W6k7AiD6WEkVPQlXEsyJFF6nM8rOEsjqgAT8uLkcE1KXOzTEyFtfvrAPM1WhdBw7oOED5gNBksXt
McnD+cjdOdaMR625LEbywA88VRdNbMcaq3rmbJIGaGcGcD9GbKktcHjeBNVrRAMoiKawE/JIn2J6
4jFSda9Qxz3kFp4PVpV4pM28n/hyf2ihgVIzCdT5z4HG+cBXK0a3X4qPMGkdlKBdxbUwapVWHnL5
EVPFWY12DbUZX0Ig4O0PDqNAr8b9eSwyO3YY6p6O30FECnkfpoQaG6nNMfi2mvGq6Mkd+JSIvUI7
1ojp3E52u/uYeCoJKAHyql/Vi5vlV9k0IsDdEC+tUjMYulX5AM+y+A3AZbKybrA/8p3emBC2xqbS
Mgusz4RE5NzxEAgFu2fhfcq9pGzPYGbgRAHIpmg39TV0cgkTV1dkwKcPtMia7BkQxIRFVJSteIO3
Dpi0JWX2BYb3tLf8cODjcqfck6l7Nm2jKC3+89QdmB7riNbyD67lXkAYLLCAxsg88cR7BG1pryG/
6BXwFNrG3d42orl+L1z/5489lQXy4EYZRaLvG4hwhrfGVVSZ0JWQfYx92D69e+zmvCbhfNTJ51P1
+pZ84uKESMoT3drMF+OHpdLBKg3uPsJ4SqrO8jOk9d+r4L1IJehCB6uXAl5njFYh9bKP6NgzAjtX
CFkzb6NsaeGMrcPHRaroOLKlqPXU1ZNutkdC9Fq3uJpe/FQxzl4SmtMhQulXYH5ON6kTIRhFhRrO
A1QSdvPfu077GLzrD3DWd+jKDVh7NcBt4B17FVmH7XQTY2MtycnCmamqPnIcz2/jCQVlMnKkZFFp
kwtL56hi0+eVMUjaE1yEs3eopgUEPdpV/DmK8660h+g5cnOM0rQ0T43Pr6AabN9fdmE2lzEYdn5v
v88pOVWZh/qXSD4qI5vX3QM9jOGREvGFNAHoXEf2U3XrOBTmqkQlT6433eOi3UjynJfqkPhNNmKa
G4Je3q1mg4nc5rzXRsdNdkyIwhugDGG8rJEN0ejYUkhwVKBM5dgKUULfxzq+m7S35wEIwQNNaGK9
Z1An/T9VTmkAEWfRehq9JF+sZkCSato1gFipRfyf5L0oPtXVALxNZrUIfbhshVyc/rWub1hwoJqc
ti8IsdxmeRawBjsnsVuJciMrycw0BLvR2r+nK0kwuMm0tSHLsUqp+yVs6InXCFs/Yt4Epsw2gNDI
kIW7GuM3F6rktUiVKf1J9cW1uxWNG0rSuz3EX5WIqEHE+tJj+ivRu1RweGOhW4Qj+cXx+9mdv/tE
7r7EsJR/MC9rWlwVvAUIaVHcmUXYSY8SE4AznVVAPo9TwYY9+cxBdTHceFBaysl0ACmDOSa7DRC6
29EMlSRqYhk85UyxWc6N8LgdYyv8ev+HW4ILsrJQMpxOAspL+IcHJVkV7Gg5WITxcT418AsQ2DL+
+jtycrJnLtlp8l5Jbn5Mf29yfPkvs7kIKyCL4B94hjNl7hqAPPgMau2I14mKoW9Qy0BeYaCcGrcE
GmIVlRS1d+ImPOPq30eF3FpoR96QPAzm1WVt5KsZbJZuYhRgwKcdVttI6d9B/TJqgQ5XVWmms/Kg
Ul8UAu/SARyv+qc8velN7nmEdDfk9FO8zFZdAvaHwesyxa/qO8LukFznH7AFH0Tv1KIfA9a7248A
Sy8/u4JX+lWji6K04wQEx0RzX9YIHHyjcaMQLvO4LdPN7qCZhcDpYqYOLhKi3jDapwO295jsVGH1
dkxV5ew41Tf/7i+plBAeZ5ETsxqhk+rKUbTWpZpBQveExNbOQlhOrokoSgskX+Zas7O+CerZOFj2
iwLor/EFmi61w6ptPY7FRe/m7O39K7OTTRuWsH9wuoWukN0yyEZEXFnQeqQsNuy4+zMpoebpTRRn
ysFCdnFzRMzUifDBz39x1Fo7BKe53AEqr5qKUIB37GhdIO7wNAUsrrqpMiGnDNjJVzh/Atr9NJbL
Axas3gbWg1weJCfqF0OquEXs2FEaEc9sYLiLnpakiZTkcHziNptweYMXkpaykF7JqfHC7SJhuA/L
LPJh7VcDHHBDMsvkC0g8Qt75jaV/7/+AgOkZa9g0sLcqe0w1p3NQfVdeqqrlYeEiAQVkvKjuK5rJ
RYu0DA3eQYMYfFeRkfvifV6ujbkP6HH/risU0RZbZOizIdL+d/Dtf1Lt1J1z1E4Aqz4FAFH57rB8
kKySlCTUrWV03FRQvFOQXUuCVPdzObnf27WXRgZL1EmpUmf706S6A/EtSbfbVG17ebBRgWda17LX
YIm/EtjetHcR/MxUrMQ2X2+h37C6ndyD5WxACO4sHYn7CkKKbdYhPW8b0nOmsXaLuxTi3V+thKPF
msKYrq9/EtD1z49TyCRO5nQ08bXXv/0kX+bo20NA+tk/4d5fYCUcKNOlu+RQ6OMZ/xHklvqP5yeY
JJCIjh0tUI7edxjjeP+8yd6CqdeoFqt/csulQXO/YOVvWhOJ3tBZqspDDuLhellyLa4/UM6rSfEs
vnXJfpbwJmkYXYgqfd9XfIzE9pCK1A/9cKOmismqaIjeXQv0A81szCt1tl8zXAHhihsdZ6h7Lroe
5PLw+FhPZe3lUyOnz7/ENwrtlFP3LvTBvKV9JlqlzQWefN+JWd/h6H7lLSKGyyNoqx6KzqCrPGXL
dVVZ6Qyv8fBfRxXyO5lyNQa/3Gb4g7geyb726Voxwnc5MlQF9vB/0VtLRgZ6uXUF4xABm9L92sdB
VPJ99S2aQ/fkchd2KB1AAIrrS5nuO45cpvfUS/dUh+IhzGMvC+EXtEiWfKXUq+4ppXKoVr2KKBUz
Ocv25j3gKVDNWZdkCg3eJyBiSQuNeErxV84UWSAGu9wdtR9EKx76kPjZx7vxHI8A3Zoz9Ir+yVz4
9mNrz5h5mVkYL6md8xHJP60k1fwjeLQ1kNjr1FPmyIdysz8ll0bhtnejRq85SuiTKMIr/GueOxhv
ykZA4tAlafPd4Dxfq5JM+mjLLu51UNJqvB9Zef5CoqoEoxYOUrklf5MWsU2H1YET0jhqGxe/29RW
vdWetWwp7zhWjfoC+kEFsXlvWI2sMN7ZtSWu/kyDUKaF+iz3hLVBEfb5MAn2hfdOAh2XImC1h8aN
6bYcF22iGwIPj2nxU5eUm5b/Nr5feKrPfalisar8YWXYxi9uLC+ncjFoMi5ISIAAlR1C9X8ZMOXn
b8pUVZJzlil6iYI5YVqIzwIx/nAefkBoJAAZJjN/3cq4WwRfGl0awtR0MW4nge0rJJ1/HL9CMY05
ThFAAU0cBCj4l0B0NiILhNqtzgFw7NgzgtQ3xYkk6nQmrwK/0Wlg6KcDW9wgWz8/aHAGyZt8jt0E
v7N3Cxhy5LhGARN0JDgOMUEIzxOwJN3En4fZsh2JZ+8hPkBsRfCKdpfDzz20qSiL+bQ3TxFWpexa
e/vePvihBl6dhP6lsbGr0XzQ2ewmfKt871BzrNDKVbOyvSJ4yjK0bOdBh2cyriNLxSMb4wXQxIFW
4EsQUfOOlqcCuvFEB+ixd55Isd5xiKN4UAiBpAo1fcwPFBcuVfC81A16J4nTR0/cthzYKuqFQVoZ
2U3nBspoMlIjKtfrU+Zuos8kMcm4858O2NWSl7h2Vwg/bhtW5Yz98KzJtuqtC+RYB1GCFqIXlxqq
tDMeFhPZGcNLnuP44ZpRCD3BL8Oy05yfVyHLl4tpd8YJG+UZdZzLu/gTH1r/pJn/hbw/q/NAKuoI
xNsy5WnHu6NuDeC9/71MeOdiqPYLO1PW8pUXPaMSgVVbryhxtjADGOQb8RPuWSOmvqCzmkvP6aOu
RH0XZZfv728DBh4oCxji5X+AgtOIIPqauCjdmIQKvkuytgbsjvsIsHcggnTUvcrYYoc7pPp0VDmL
NPMKpt6ElUW8zzTpd6Dv0jn8mDLdGOIxRh+AQ+pb3dxnX1fO/AjNSkpAosszBhNOT7Gplm4+Z3X+
z4/Z9m5O1LiDpgh0Pi62qOO3eRVhYOu4YL5Kuly68kdsluxns0WpKDXuYg4TppFA/KKDPUvsT94z
mxeYdqtaRvtyRTjmr658+/8rJ3IeJHBcDTbG7XqBs1UckwhFvSxc3lj70ZAQA7bzGA7j8Mkso4ap
t8xewdywx2IohSocKs+1wuclH5Jmdy1JeuW13wM4sN4blNmlfLpdGyxUpVeuZGdMsW+BqcFVo3nh
10Ydkz2iCAQVMgOWnen0+wHKzuQttpCIxsGab2Sh2VGqLHKZvy4tBlhYDFOhMTEc3Z8sIp5IT5Lo
JNYzU8h+yN/o0TKCbzLdR3ByziQqKVcE3KZPzTsX4RURC88N8sBHM8q85hc+nLVpIqCj0LwL17yI
ctANhAhf+RmA336uMkUyJHLOz2bGw8LnjCbTZAlZv5tMzVat49GJuMmf4PV6q1orIwtP5dwk0DGb
gVrPcByQUY0NGvKj0qJlr1c+KwrIWNruc2ywfYulZYwQo5ND9u81pDcjl0Sav8RwXxIhDPReszyM
B2+Yl2vvwOmnxJusds1zn/p0gE7z27Ro7SxAyG1hfRM3jDynrqcIL+O490YcHeODHnx+lZfMXnNO
IvD+3+kl9W8o9ClZO+yluug9ju4HTbLHwW390OcRvN4kSlTkj/dNeWh5pbtbMfCRDyseh45xAiO8
QLxF8yILLXt85i186rixx00Pnyawl3xZH0ehcX9grbCL/+i9hMfcKsg31rLG3aV6/HVYfJ6hcO37
4DERtq9YEzuW+nx8c+m/v6fUI/DtWqQKY4e8SmqFn2/8ki3e9GVo87P5fzJM5QMBbMOyCGzulCc4
JgLXWOXuuk9CRTMWm6j5o9prSAhujiAXgna0n/ZzdWmCZo0aowxpbxzsXKiiKQSQpmGgr4yH/5rK
bjt+Vqz8xdrt9VJw68Vx0DTHAG9qebDpn2K/HeNGwOPhg8itvGcd2xA0uTq6Jaj2Klr0Qz/TNnrF
GsO81CILcUVHy8XtvYjtHXlkbXSPXlyYfdGzIg8BaeBI4VusVD4zW25V4pbYlvM4KsADHqudKPgu
pLbSbSslnF6ve/5dzf38qLbSnMqYsu6pZLe2Axt1Q71lVW96kyJy1o4/UHrJr/6dZuBfM34ZvdH2
iIr9tqfrAvrToX76/MYuzSomZodbPEQGebdtLVmjy9fZHiTNva+LhiL2tm02pcJZ+cJ3I2K9/sM9
G+dbPnWyW5Sex3P5SwTrBJFeq2m2AYVx1HNEVAkCMJNlMK2qNDdEO/9w2ez3PvW/seeoZfjLsVhC
oykvaqm9d8vcRCFZBGdG3xlWGI1gw/I0LFky+awCatNrGyyHED98RDmCafPYNkZfVrzg9EQkhN09
T4fGuVsGmy2Q5+NWYz/Znm3mUjmP8Qu1ir10jdrrowhY/YRokHRS/4/8uxs0DfUadiJ7BJ6eZj7t
3zvj/+TLnQw3tNXnAe0N8Fu7NNwouuGLMUQoN052Acp1qp0o44MdCQ/d46S2Jb/dB7K67KLZ2JBF
zpZmOYrkpDO4+b1o04+nS3gfg/682+s6Cm3wT+lEBTEaAR6ZZqOVVtgYbxVt41n+F1PUsb/icaOf
+V55Az3Aockq3Z7aI4biBQ9ck+GDZ02iUeO/GQSHWP1uCASprTLddstT+Exv8cFDQUw6jHhhx9mg
s3g3Fj8Zc6SZMrH3WJKomihmQdX4uOnIj4h+MrB9ijBMoKcJ+f7yae4RiFM+sC1sqzygQmI7Kwm3
qhh/uKKTBKN6phknqoeA/G6H4ANWtzzChiaNQVkfF03TGD8Wo8uQBOoO0mt1EGLZ/PnbupnPuyZ4
iRmNdBGAGafT/XZQv+xg0u9G0N8bu2qZMKqF3ncJMZww19Xelupk6DAvyRJyMdlRggJ02w4I9nye
6ilYyqtPcogsbXRKuJObK+754BYrDq78BHInVueWNC1TJl3a78+o3BvZLOia5Zu6nrAdp5CBRjAr
/JNJyojgDBqhYUa6snfYzlJHPJqgHQKqs2a/bg3Y+JNqo7o5vJVXhYv2XG6baG62xRnnSEaNOkY3
R5GjdrXiaZHGFdQain5Dw20Dayh951KvXCGtEcde+yS/XNmn37GgLWpksj6s8BmjQd9qBjMUe9B+
8LcSGy6P9lPSnjNUCxJAXECQX2OUu4loTwaqRfuVzwNSq/kOq1tCi0EyQTGxogj1XpOFVbFVZxlf
ibFro8SxCNDdaQGGigZ34tLk2WC9EoAaYJ1dyuf/oK5QOxB7upERsWZqDgmIDu1BVKymz5p1U6fd
few2w2x8oA9y+L6aW9fJMbtLBBkNaPCtiYnvR7PG/1Ftm3vWUeRPA63Bt2SqC6rGNOjOOkA3TI4x
XsQu24n0kebZNmjCHf9AsH60ZaOGbDL8dKccRT4xEopgL+7zVCg8VAzhtjVCTiQsg4GF56tmluJe
dhmhGHBjOCKdXoGqSzGV/7Bjdts5eozlyvUAbeDgbikH9sVNE7VLYsW3DaBYFn1MGD2ZdMsymr4B
LOJ2ZLwtk98w7RcY5XHJHW6ZX6Wy/OtovCcUgq9lu+ztcq4H3orEkXfoGoBSzLQn0gZ//61oYiNK
osKlwdrh4mP+y5CPAvlgdttUdtH8KM+j7QVz7w79Dw5nfcgYC7XCrhLoIUIQmU0du1ff6oOIhoo7
MKBtmFcgU+mHpm2GERC0PmbOJbqUdHPOBPvo3F1MQUtGuX+FxagogE210aop8mkspzU6dd4f/gY7
z1t9H7fO13Ayu7w59dfKR3vlcTiC0hKyVwQMdw8iq1hbvOx1liE/zibIEE6j+LibTmBgeXz3g0lR
8N9EgWnR+GGDlWxrFWmoVFiaig6B3UM0gX7j9IAYWqF1pP2PUWRGFQuPfSGZy+U2POItH8dXH+9N
5+xbwgUj5X1m3FSPPWtVLb4Sq5EUwKp8Vm5pVUwySIcSzNKJ+HUAEu44jD+lAXTLsuLz2b49YvqS
tj+N4lVX/nlPIgAIj6Y6eKqOcy/fKltzaERlauZXV0PPTwApFoCqyc16GbVyB1nlSTH4O6sA+Bdv
V29L2QWeQH2/2lBwmMIkOsujoZ14tkiAG+qKd96d6hqlMVXaukmM53XaPG1iVQZMZdGso3i5fwmu
yGvUliCClGsVsvRgE6+A4QYLyG/Y/so0m8GA8sofVNGegkB3DB4D7C7w8hvnC8vmZDBAXVHRwFE8
3VcengQ7qw2v8LJlZURLS8JAaeW3wEzg45kqDjKD+C74X2J6z5t9wW1X/YdHI9GNLPBAf0x3RWvZ
0alqauXD/n0rc4e/gzQnR2fVvTNjbQCsplzL2w8LA1g6Q4t2/1UbAwbV2PWJhZEU98IoVzhyjcQn
mSunIdW+tD+J2Wf99Jt9cXRGV7cc1bz9VHS0Fxe/zMeKJ+IgZZ8EJsuH7JWtzUXXHLq7v3AYxQXU
45LzyrpRZFFWyZDFN73pARqni3b0fX4UzqOZMna4KP9eJyJMSpk1hoUiNzfFf+dnZKyYVMnQzFXy
NbSu30EpkVKdAQD3UWu4ogRU3sCf0EDJSmnxn4ozn+8rucBEo3lCPbye9yLN4MUShupECkVDwBnf
1imJ1cCWjtbP2lOSGvhcEPG/hNgrXJQNqZig5EMwa3cZNLY2vH+JEn0xHhrlhx7i1WPmWx51XLBT
RzuJVOzRrkbeqNNTr+y19d8nYgp76ufBnU/RtiYWPzTNvqO0xzJq3sRfd5RG7T8+smdvzHji6dOT
QQ38a+WNPJN/KAl6xgvI1zbvZFN05Tb2/IOXYvCgnUolZrrODWNGvS5YnuH47/2zJQ63q39laLLs
KQq55KbI2O/lo+CCz9qIUhDsYg5z1hadeX2+Q8xJyzuGzLhcEhicEBxkvpIFdwjczIFlPprSR2TG
gejBohtUz82oH1M4+199Y2c3HIt/+s5nClN/oAqzTgQ6z3LB+2v0C8YYfohuF/ixrOEksOT41fyi
PcsYp3zi3xLXveuzkJiLNu5qGADwL+hHjHMvZw7ZH9Ewum0cWuANad97eqYv1bO3JMWwjBAoyC/I
7Xa7Ym0gqRuSBq7lcx7+J6rAXiWWt5+hY3s5HJh3NwrDW5u3j6J4WhO44ZXNSMsAzEi09SQ4lz8A
+fMgEUEBC8f7/iAWwW+hbOq0N/xA95XVFju/bcfrAqlKp9DFRGb1ppa4Klng4DrnlnTUxqsGI0Nf
sT4LxLAoMnHXqybMhXhpFno4Wxnu/l1HsasJvdiRxty5aYz95p++8QDSEyYNDVqxWRP/BC9m0zcn
QpiKy5ZanHFH+6wzZwMNGOz410gKJ9Wgpc1tjrVVZuTnDWqZ2bEfPprGeu/IY0A9QKbhUXn1Q8OC
iFbjIhVU6BC56JUyg1FRo2cJqSyyGdQsY5cOyKajP/3qGjf91EiN+pJvoJo1B34NtUVHROz/Xnpr
8VY8q+B+6Q8aSJ1wcMvQTyjNky4UNl6UD5MJ0AnogdqFMsw8UKCTfiehbkIoW+SK4XsrLauU338J
CHZ5SWREf0etbLG4Hg3Yw4gynrsWGWgE/H/61T5UHdKntW8PpdyAKQViE86A9j+MV1Ix+Wnr1g+r
IGPJ71RKewUCnJMAl2tZf57QtXkXDAvjqD0MYsu1ihL4d+2NBHUH+xWFqw0l1GewiU2bzsouotiQ
9J/pdvStI5QY7cNYuuaHXVKQP5dkeU11Oiyy+NaxaKP24JSeAqZM3hZrBUyWbvPG+outvIu3nOaH
L2lrxkaWJ8TB+aFWniiImhABc2JiduXs5sfwoIRdgGOSC0F19oQNpDAt94W8CQz1grAgQIefoto/
Lq0lBRsu98NqatxZGcCGTl9w5AIbi5Uv9zbwYoUUXKxP2EEl4ktwjIBv56IoVDIIsTy4BkjD2qir
x+Dh0W84OyvWS56fv8DOjLh3HJnY8GTq+ec04yAncZ4sieBEJaiE/4LoJRVa1egp5yfAW2u/BbsA
uhnnXRIwNjrRwISzPLC/toCgNCGNiT4d5+L6Ao78x3itwUK6369nKzcAXnMzWLUMH2LkC4TphiHb
uAjO6GhF+COCsrBGq8fFOjQRp29fo0K9HcxSlE9XxRVRmJRZKH0Ey4DJX6wCG3ENbMF+TCVTNlrg
b0INsklYtmH3GwTbq6ntorLSJ3CDugsZgPIzfD3IYLZZ70JjShPklCimuKs6Q0r1/vPeok61ry8G
7nITblBudIpCdsav/5ogsR5P9y2gVz0jsr8tCoioAZmf46a6QIdEOKn77mS6Mm3D8bwjGGwtn0ex
eWPi0uK3JthdfSjNu5s12b/jd9kt81mTQOt3RmhqZPPgvdk8CcWlZzpKKSFGF3ObZUvvuuAE/ec/
TBBiXcaEeHoQpuZriOWReU/6Syi+XtIcpyfx0Hsc9TiJj1D9xUeDC62uHcrJ+q8mm/6qGDjqvbeT
CIasxIvOtG+FnujmnU6JXVzyuahUAo2n7D9/xLcv+vMzO9tkbpEjt6H0SWgi1a2Y8aTv21FCxwYP
uqnKWiE+6BwMevjAZoqUsr3vIjBUjwMQXSc5k5dyIh1IRTdhw+PtgrhdO+FQS0op8oI53gU+36aJ
N+rCOXT96b7y/P5HfVf41VBJF0brH7I2AqUkJo/rYv0QWKm7sMNSbvqYywApp55cvu0lmZRz65Rz
hqntjR+6A2XPiiHD95mXj3Sc2zMxQorU/SMxr3OZ29vXXpIWNM4jlKDQL+3xEty9cMRuWCE9Er21
g9TnkpyfxbdfyuUpeLt/LOEMEtO+4yi+uc/0r5TlUQThTrMYhrlXT12de2bih81E6l13oWKYNazI
lq9TUZYNC8+13NNMP/t0Gfi2eORsqDCgj6PZMYx0zoVD18BUb4fxi0zBLkX6sshVkVKGxb9RzWAU
hmAf2FXqjGXtxGgKXQT1w3NCj6JxHb9N95PPgg7CP4XzidV440+yAKDvAvYYvvrQtnnvSQp5VW73
PD2rlhOENkQJkOoQ060DOIB1qYF4sh5EZhnNtQ4zLXvRKPMoAMktABwVN4Mgqckddv/7RzMGxWwr
FoajBwOvOa3KnNS9KrARR99pU3pq8WDpu5Kszrv8zHU/KPYv0Z+Ws6liDJdEZpgNz7q8rQDuym+A
39QIDeplnLFtmaRogj/dAUTZngXsQFXVlK9aXCzyGVaYm2KTjWsghKoi7ay/mptyp2DrEDi+9S9R
P4A/QHue5egLIYM9bS3p9tq37yb4z+bPEWUh6evZN6uA/HuLZakonGC4384K2fY2JVXCmJ/7nqUV
pzd3pS5zZyAb272e9AxOkaqn7zTLM4aU2nu6cOd0Iskgk5vdhJZ7/CtRAdC7N0verejSR/2PdRw4
S1yTs0eXS0zTyXZumzP/JSDVIT1hA4a5XRzQ9vfVukDqAQLStk2ybVZJyXKpynQzS31h4RyNPCob
8XskZp9Uovhx2PjzTpp49erPzpFYP/hx/M6RmjQE3TgBpcUkHuFFw/JTpewEfT/5gX2yuwPqNl9h
6VIzdAyj0V+abFM5wA8vGNMP1qg1noE7JvXYSaEnD917dKF7UgPgFvFDOlJot/tWb+i+4WJoIEjb
SOP6gmbkQUL9+Z0MZATWLakEbpA5BOdMhixuu6nHWdJIY4uq327J0gnJFGkJe9IjZQE8UkRGblVb
tBCIu030mFK0jfno2VTbGh4HtANDMN42dEU0E212b0NjSFboqVPVh5sOq5mYaYlC4NnAi+A6LBOQ
NxHUI5WuHHMP8wSXpkZypqKH/jPUAjLijTAuj+pakkGUraWOD3kLRZ5yh9ZCupH6rPHjcZS/MHTu
d5p5BXZojEspqQf2KHSQ/+BKkFpLC9coQSrniFT9HV7BhNH/1WEW98Bi/A1zx6xyps8ng6zmJiIf
IoNriUTIVmQ0OWPMGltHUXP6ztgBxgtyI6zf5X1034eoZu6cvzfX5TLlYBnPiTpWdY/Lxpr4brZY
PxJNOu4Dvl9ZtoSh+Vyr32eyd1vzTTila+jWInxAr9mgXvkDf7Uot9kuvpOFcoKQVHA8DWmjCVZq
Ze/cl1cLYt41D03zMTStVAEQmzGlDW8r0Cln5MqwHVeKD0TuXCKss3t+9XZQiTDYMGkNyNSpQP3V
K3laCxgfFFpMDpIcgiXKgPPZhUy0ehIJwK6v2LCGE1dsoyBCE9bziBYlHxeS/c2h2LrGOZWMuj5V
StJ6eaJeW+Cc9DaIhcKtTKJaE4rWsH0+hgJ8POlEAcaJYQQ7oOybcTZwwDptdHIRrq1R1tR8aRup
PjWk4O+AiyA7uaiUZoHmV0TYBKu41y9/YRUdlpyRm4XE2MBMLPvl2ropWpwWxq8CAC2T4SwkwMwp
JaiCCytSoJ5qV7SDVL7WdCmppR8+68XzNdiTiWsTNqlIcIupNjvLq8JCVDR1rGaQBYllDtwOOEr2
nx2ZdPZF6l0gTIOhxeZDAYtddI8YFG5nYnxDeudtBW5b9bXtkMp4OBTCeH6yzeBDnhiL3IwJpt6D
+uz2eGslEsGPZAhYDRCe8NOfgAC8PgHjQHrflGVb1WJzCgy7mLdWb1iVsa6iSWaxkA8LanZ6GAc6
Z7oCQolQvXUVXzot6VrFEoKMsyTcMb1HmwMWYb/NO5Pzram0wjjIjd3RJHk6nfy47gGRyQ149RBo
cVTPB/pYavNFH+nWWkHtgWoCVcBKM26BwBst7Wd5PEACNHqmts9pxKJw+GNvAnHd7NcLSQG3kSwS
EnXlOHl0z9DIXtGIhCn6/MBeT8mgM/0zYaGa2riegTfJWxUpPNow/LopH65gUarTLVcP7i9T9rzE
YMoY3D+up52nhzFg7LXy3InyzjkW8BdBOzXBcOTFN1j4fBVf4NGTK4vJxXRyaGEVhkdmE7vgN5+K
2qL6vrG6qEIEt7u5A8gv3aPQvJ+NqgJJClQGIEaM40Rrwwq6WUpuxw3kboFy/UEiXqp+nNIpPrK6
6nXCvsUpXwneOxLFQPtGbxvca86sctZeb4S3fqrkXRgkNc331bZyVLRG9xSkicqe4jqhXgNxE8MC
4CjD/a5h4S5RdMTIEBWGyf7/UgjOVt/OLPlCFxpy7foK6wak0xi+vBteU26vj+sf+mBlmTA0zE0h
wLeXFgADpnaXOaA9hl9iXG5IsIlO6IVF5OBGtGn9JORDgj+YN83aeW4ox6qQQEhhKCBWgFMh7cKs
PhGzBScuwEc9KPbH+bnqqQCfkUq9OVz5uX6mbghI+GlBk7Elod9Ao3Ojx5c2+hGCvietqOqJzrhe
wZxhkBiDFgEVDUiBqZuney23IaEpffBkQldHq7d2HQJZZ2AZO88wq8rGH/YWHNWtOjMrPKKC7n13
z3Z8RDpkZhhgUAgg2Ajk2Ns2g5wtqtFQyLozi+yxT3srcbSo98aVnEMBRmbmojPnfQqZKV8vMlnJ
MQDp/MAv5AXHQsAhDB0jUa39MM766zMipkXMCP8vsViT/TJLcI3EyWaXoD18jgA/p7fbAM38kpT4
YNQkzg3rK1yeazx/6236P0ptZ6ZKxSsaJ7ZnaciKqytef/Fl95quOhCj5eB3MBBeOhAwXQ7vVhao
e+POqEfGxINu5VXcsWK/KOfnluit7D0MefnhnkZRnABXqJw4/n68oGzD3fzvc3Dl2fXaHnS5jzEr
d6c0f9WQ0VZq0ZEUEqr9fx6YaBgyLrWg6ng5Xi9lk/pPGsYG9WUrZD1YSZUkaovWIV6SSQg1I5IX
m64LnqS2fVuDla5bxvTb5gGpDBzV9lOlHzRcU05E7TlfvfSo9urgigPcZoZzGVxnBC5NW54/d6id
Jt1vrrCzap+3VBXksj3AK2rHvPC1VyhLcx+e1tUZjoW4/u+hjOjDbfnB3wLNIhAUmBfO3UnjGMVU
wJgRYqPrAmK0E1HcFpFzCkFlNBQVOToEz2OKVwWhnHF5ZIUhzy809d47YXjat1Ul6varGIhr74+b
KBWaCwlOagaaUpXGY0mYmw5IUJfZZ344aPBOThGxNAMsRr3AoRmFyP4ImXO4morGRCRuBYNlvA8S
T+QWY2EteSeJc3Sf6WZd+ruA9VV/4Ta0WFnG7OjPc772RPR0zOQZphxuScYNE/3giMnkHwcnyqLV
PzZeILqGsIr0TuOG4JRDnugV05zwqWV5iCKUVfI//dgF1kgDWGT5JpqniIPYBwbAjNgu+SoPnNG9
zJ+bvXzyN8TIy85GPD0CxH9Q961asB8gUPduP11WWOiUcecRkCyJCNz/H4o5eLjpe++8BzOFG8Ba
0v4Pm1hj7LFcYG68UalX0d8fUIOcijbUdnh2U4youFJBXwWoh8bJcIEpccoVhw42VPjAs06xHLR3
sswwpDrRWyoIvmaPWt1TJkhLncxeIoAcQUgdx2/eC1ApDc5KCvN/4p4h9JT87cBvkHhlJeuTxOh2
JgA6YrQCvUxL3+K21b+DObuzZkybCeG+QLkLwwyQ00m98ZyR/tbe7fz41ax62HEz8tiIker3NuCL
JlP+qpDayaRQm0JgUmfhvc63j2IHtlH0JAHE2YZ4todsgaeFzojWJ1gVzCEaHJuV6qzzrZ3cgkpe
XBMaBpXms5xk1oXsG64tHM5+fhjWImgg3aVzoNhQfRUYRm06/+iSKQeTu7ahP+2K3WtFXEAM9zvC
9Dj+qIjop6rPQLonODzmK3owRUKGWNqx4y6fyzUBcbP+ttHiDZjU3CVqZmJodWJSVHcMGYXXcauD
7MOr32u1OcmzKj2sRzgyvGu5eTKMEw784G7wqmFS9KY32Y5IE8WzVj6mL+AX4PQYISg08/C8FarU
FlCYKSjLw6Hec/BYaIHv2jrHdpIiqYVUBY+3uNFFK62KJCAWfq6KE5QuwZ3xCfyXKaXYC5MJ48lL
PlBka4ouz2fHkCqlSTWtgaA0xT+d1UMQag9prAGxXKaEHLDW7+0FX51hzAHX3rKzgJ1DjBIYoBtx
X/E7owdByFNpYj2Wh4oK+D/ic40W3tdZpqm6meDlb28g26nNi6bsYskmaOp8seMR04UHiIWnCJv2
dfC8CzCiBNn6sHCxatvSRp55xkuF51VicLBneI98Sue/vjVjwwRLPhpdRaOWWQ9mmckGL8oPS13s
2zWDX2Uf7uLVu1SfShtDugvcbPZOL2FMI5ntrNrNzziesExt3YrZ+M2eWcvf9PbdSWRdJJW/cpU3
4uOvSatWUGMx2K7cKg4uD5Xjz5QQd5OmnkLG3boOIurwFbZyPV26hrs8+94DBYGZYljUxQeg3H9z
j0+vXh0/PYHXOV22RMYNrUyyT4JsOHQ8g00fcYYr8PWyUtJjXwRmKQ52I99I1CgltOzrOXOpQ7Lm
ksVDB62tViKbl/5qrVCmd/NXu/VKcD3J6y26+Sg1xYTvomh6xStXQt5vFECjUj5k2/raHGiK9Mp2
eA6YXkeRDhQxQAyKDcpeU0+GR0qM7VVSm9YM6o9Ij8jKOiwE6ACy9/1NAkTUPXPqr3Lm3024PIsk
DYJoUXGWWFDQ0Jv8CxQUOVxmIvOhZLCRYD4brQnvlzyBKmFmS/IKTSxd6tjrUNnE1gI9gLwBibXU
NVRrmXT0NGzZBkSAtHZgHkXii2MvZURJMDSSa0iVYMiqdnrHVTWR98yEw2a6HMOq9+5+Y+HcNeb8
Oy5qS3HFmSpaP87+EBqb9CR1BUvti+Fn6RJr6xr88tYMbaIhJXoAhyHwpQyME1twxblSsLSS/Dr5
Etybko22mLDaOJGbwW6BZlvW1n4ApH/xUuf+Zqf7OgUjEW7/wCQjFNAeSa/mbY4k+BMADDM9p843
wVMMpk0O6qmhNXyYzCO/uBQKp9ZGiBtkAxdJwUunY1vy68+WY42Y3q0Uai5ahwOieuSD+FC9iq8i
LMQx2SREKjO1XqJH6LUwdXy01qhIeKatmhy+QXFRDCvx1iRKY2sRV5CtZAUt4/SSXrXg9S+vTtgW
de/wmWNoNVE8eA3v0IJxHhTnjGGm8W+QP3hIufULfGakca/Rdu4AU4EDJ1ffQwTJo2B3OhGarWtP
+gye/lQkiCA1stcksexn8mgRjTXumHO373k9KvTzMIIZFiRbO2kqZYyr73jbp84osZ08aLfyABlU
ktCQQbhAedBKtNLJzO2BsxytMbYaBLcNeJAYa9sbhWkHPQrP7b102aBsdv2zuuXlyNleW2gwtowO
71hHCE3YDXZ3jPYQntiFa0pGpkEAycnP3uOIinw2Rg6uoGCF8RAOeD/Sb1ol87YqEXWs9D1ivSj/
u7luQB5qd/YADeN0Y7/CVz+EInO+Ns8V66Vg2yZVPBmt2yu3QtVqU6jAhh+BU/vn40n9vFJrwpjW
an7LrHZ2a/tC9AXtiSfJCbjeqHRM2KBO2XI4B2ZU9lq/TLIOoU+rapYaeUdUvDxN2x2mv0BJYm93
TJbqKLkrc1YHzR4uE7Hqq6UN4FRLkHQlofeb9IaBbii+xPx1pkkT9b0Byln0vfBK+E5RGAVk96Pi
dmvrp4CEJOEscygedJeZ1ktokgK+I8WvsVwv3Yapu3dgGytWNnZsYlcfMKQe3l6El+YlBGHvGZuz
MOHe99EYCPs/Ao4hHuEFmOuv7KhpEkqTzDkO9WbLid6WTK+Bt6lU8bTjecSE9Z6ckjl3Lz41XkMR
7t1126CgjCuKhWeHnFPs1cMUmOTVfQYeGQEvAbwf6e6QAk+cqpLuha4E4eYey2LE8nzo8dpML+oM
2PYYYE1t0rgGZs/zmqyfai/aorrwY8nDTbajZin/xlADbsLKII3cRevJao9mRw4PnXLiRKUSKu2n
0Mem+5hsgWYPFB32pggL1VfzIk4M9qBFKnJ9w8jzYA5HJ/JX7p+oQZpbMJILhvMrdfyyYhdYgZv6
+LgcjSA6T22/ykLUkGy6Lgc1s0Y1XzbE7EJfBMxDVtfQMhNH8BsM+KYEYCG3AY39sGuYo+mFpzk6
0ajfix64l0WbEkWPHqJ+n0LnruUvR9vG27glGN9RYNgd1aFcq2Ua9fT3SvLARiNOoPmrpY5W1gA2
2TYMcLCdpX2GkPqDEo0F2rDIy4Z9K/Xz5xFERCRdFXIWtX7h6OwisTxWOMlZzIa/VwNJcdH4hfMl
RbWAOXl+A/OhL9abozG4MQq/AQVo+jxCObzP6FrMSdCyOBOWCCn29ibtZLaamk+NLOEpTGtgJ58z
BFUsMiwXk7Olpo35baOtwdQoZo3bb4JBbH8FyMYOGOkosdvA5jv4jRPQsWz7orSpxE+JHit6bq3b
AeD2AwA0ET3sjlk99yR4AGKumlqEdMqTew+jnJztYJ0g9G7wlgm52Y7pAb2yY+70BopxVZ5dRZD9
X0c5HTzuXra3bPnrGoTU/FYolaqXocpdu4KuCKO7JO6ZcbY4bsRdHa9KiSeQpNmKFnluwQfGlgT7
1Bb7hZwPBP84857xmbB7B1SQSsoKbBaDGKHJQMRRdHJ9ZPVHwJz+dlXPrKhZtK5+bxoBZc/InKfv
Z5Xu3QeBKXf9IJFTJgkSSBZMBTXv8/OYhindQUsY4AxRJTUpRx8Nodxh6dK6iLaOPdthDGsI/Kg4
lTPh72o9iYJC/rV7Hj/Cs4jHIxabngxfqRpJIPxFhZY6t8rcc6j+tIiWvYk6kgxS0q1Tx2CXEN+u
c1x6bQ5Kfo1sqmws4bsEKHWcD+JQ3PUar8bo14yEOMGo5C6jsOGbTmkS1vYrYfWK2qxO8IJ+mrpl
LfHVEd940MN31c7m7LQSn2e0NFCpPlYo8L39moTV5hvn8baVVoM9pJk4rBAfqAD4bW3dFUmnC1Yi
G9XCPoA+BzssMo9cM2pPhNAqb33lUZoUjKrb/0TTdh9yy5fIbqecSCABE1KOjljNL5SKgspjUs/f
WSfa/FHfjoDAXiexKeua1luka3BH4fUf8xRMWkLQmeVnHlZh1AtairYbIkfDb/oS2n7GIfBxYERv
+HZ/AvasNzdoxm+HuO74IMvUAg7BHNFlpKHdGXA6v+J1uUA4czQjc1E+7/FSMUAz9gl7bES7K4zo
IGIuJ/4TsMiXOQrHkuAD3oh9YUIz0v7dIYT4TRPmHObQ1C3RiJNKCDb0/F+xO5IkOLU/IXIhTgKu
REL41+sDFfCGp4AMwhNevWmENjsL86CCzbD92HiavzlPQxm1MaRbDA6NZ5ulYKiN/wVj6UeB3Dns
05wlCXiL/rZSSTK01+gHG4uZQSpiAJBIPrioUww7MvhBV/Yi0BnyCxfzVwyT9GV7l7R3upY9IhH0
VwiPKUu4h6X7tIW7KAYgHCdBLtjobAkha2Vn1ctsqXJSaGGFm+4ysoruhPGGRiLS05fNgG32SjHK
9UzCsXYQS6els3IidwB+Wb7hv6HBw1Cih2NZRRJvov848YT1VpXIDPlywG5U0OK7r4T0UPM89fVA
wp3MMAeAc8OIcB86LeFKd0radoMe72bzS4iLwRmzi198kfusPz5WiGtVfa3fwH0jcNR28QaEzoDF
9bSiBe4jxB90KBGEQD63wj2O1tv5nPEYaT1l/oMDOF6cBIDwpOJb7LGFzyB42+/hljJMDNF+pMxZ
xKyepJWUUNGFgN8bwEWbCydXz8G0JRN8M1fwmskbzTEpq1btqy7J+Yi1ji8P9gtzmTknzKXJMkNM
Ob4/ZFEELINKSH3uRHWB6yzGWzWD5Q1d3IBmyl94YBRXSH5cCmjiWJJE3jPYDIl2l9fEzEYRpBSq
HHEsqOOUAk/1y017iGrY7JPlot1gIaYgS6DHKBQYd9LvsDc8SmbzqG+et58MH8loizVd1t5oOqAg
Qiu/kl/Z0ohxzGFNV/f3ToMlc3UaHgLX0qnLAzJaTbOCPrW8xhbTPa1xH52LKomGbhfSomciurEO
QmSGaEuAsz6NBpIp7ysIWshVluFvAMKHbkRJkxUlzq8LZ8kjRCBQ7yCt0YV73/Q5Ir6wqcI8pJxg
dW35cnwyJgaGE+IfDiZoBNRQenmo8HcRS/1FOzOZHGFIGWWXcigDZSpcZ1MITh5ouRMLBmbwJP9K
Xqc1nRjlL62mBsnzn1caSjqKetezIxzdUSiXjy7O8slOWR9bwwJt97uXUKLiBChaUCTEtFTJnfhW
VvqONxfV+/Mq7ehrWcv746+LuMzrTSmLtREQ2Psnortif8Je5TSlb6I5HKMVbYfXQ8sFp9axJZ9x
BJwTqo2zqlOW5tBKLLBVOY5Z5KDpF3MmjRkmWM8a6kH/Fg1XjGSNacjWUFhXfBO76a4QIxTeio3R
amTZ1sjEpFp6ah6tFcxVo8qyDCAIQOBb1XiANCr3DKI4s3ZEvsGnWW557lIpKMxXJ+2iXEeS7KUD
qWn3om5KxmDPxRNW6V41f60cNM2zHc8i0jkDTtRAgBoVgc4eai0zL88ZlBQkz1l2v6G8bn+0Htis
h3+BlXelRLoDi+ykHHveo5rZrjlrOGM1e0ZYknlgNDUQF4aSpPABb+PFSnEt2g4jqxokfgBgYeU7
2ZWXz5DuFosRNM7DrnUPsDtkHQ3A3piVrJE2QRsHtyqa3DHYnUbGfaqeYA0+LyR2pITx80vSd90U
hdRK6qtCOlVxaM3ee/d8Irn73i8lFA1wSsdzuBXtvuH3iYS5DIGuIOfgbIxZOGo5zRPMmk/UyikM
JRYNrcveTXXvOLAsnhoIM8XmfKvKQ/+xvl00E5W4aBKu1/OdDU6gMyxZNg+Ox+MHBWTv9EeCJxti
2tUGh6AyfIxPc4syQ7Fpsfgh6EKMQTGLtOPBRsdx28DZZOVaG0q0D7K7NJq0E5owDaCJSiGft23q
jtjXa8InCtIxOB2Vv3fqM7QT5QjhgioUGgL7ntok5ch6547np8k+k7sa0iXDCajuMEcJt0v1meXC
eXgC84vhC0goALDeWkj5a1z7lR8ymp8KasfW9IWA17ajn7pfLchcnQ+A6sHcIjoWCfScI+MmhAj0
isyP86BLqxhsNPcvKi93VbZM+uJkudQKRtTmYIRr4iN4hU/6DtlA+wTl5nglBVOFxpsJ6N8CEXW+
/q0vKmoXOCTJXCPkk5t0GZ7MUxXO82SU3B1ROn49WEcGApl6RYY2vH61exHe3NgDa4ce5+a8PPgG
MzgdOWKwJyTkdlkcjzLiMpps0V0PWUxVsIfLMOMYlDutfKZUdL4thr8twOLZuMFzXKYoz9F1G0vh
EYt0gbxpQgwjulD1Jtv7A1ebjdqMj+IqYkrWqD7jfQyE+rluJwOShCERR1b33fKXn95kRIAX2g73
BF2IfjKzsX5IlQ/cm0XaNd4uX3mixtTnRP0ZEe6VKX+WJoVFe6zw4kVLMEKZakZwrwXrNV7YBJJn
SgUxtom/q7GRUEmDJyz6dPPzvPvOz2mnSTaCgnyacOKpcOEoeqUl0mgyiBuGA1yp8XnQooUEbqeQ
iguJaKx++XnRmjtdOR2gyvlONghf/mYwMKtDNhHwdy5aUjtc+BLU1aopbl/Y0wqRmRimLfw9/bAw
CXPUik5e23jNdpMtYhFHvh35kcYXwyurIkK8jI7SOZMhh3jQhE4DqPv951/eyKEv1s5d6n+6kvU+
TVxo9OGXGySCVmjLqXx/FGu7GBf29QpRpu0zXsqKyPUaoTdUzGoT/Gaeq94Z8u7+D3GhFva+9HNh
ArF1rEF5G5vLeNMYMh0OMs+pbzNOH4tmM2It9p/sWLwdJQAv88hP+yI+nWryDBX+XOLOwmP+F1eB
DSrmnlKYuO37z9SQvg3P3XP8CvBig45yXwmmNKwYvMIV3NkSajDJ/YzotnqnRHpmkl8+Xuhv8UnE
KoQFeMIkXTtKaaro17amxfGoSE4xDQNb5gSoDA4jRpAxdu2Hr4iz/oJ+hwmGgQgy+MZS8DhO7XIM
khNR7kf10BhcWf9JqcQfCGzVl+nS+8E95nIeoIiKOp2MPtBOZ5K3CnhoBdiYNACez44j25KxkhZ9
5g6xkTCIhsKBV0q+3aXSXpXOtOApCGI+qxq1TqVpRVXF/qjY7W6uiJFc7+afUsEAKIrHKi1ebDeG
oyeXbFkhFemjvAJ9hDZmcy/ZNyw3T7BxeG/57UtrMu5/FyT/NOUiipbwT1gU/NMoaYzPmt2U4w18
6EnvhxII01UIGoNjgjBJuL3TUtiy/GI9CY5/JDSSG6YFwhj8umsDURcJW+KLrL5Wbcrz33Fj5Qrq
WN3wlLr00DuUy1FMwn70OSqzoVtCSoXRZbDGiuAU9+1qRBm6Lbnrun2EFtWuxMsAkQB5tSwgUKFe
xXf2JJ/yWT8naa21s5d6OJwzLRevy+oZp1eRuASK29v1hQuHT3alzIaJHOqas+iovjUDQtYjfy6O
RDZd/twahEfnuXu/cNgZPy4+2wPAsQIeYZ6Gl0d1dn3f6KTtDFLWRy9VFj5QbVTWjBOvy7Q3YUGz
PV0bfDz6oM62kdiCftRTUjnVid2OyKj0XlZcAQEdb3VJsEyS1d+ul/kXH0YcsWjjICv8p1v9Ds5m
0z0UZdjX385oV+88TbLmQ+m2rDOf83IE9A/oMkfRehUDdOr6gksBQkYyk0MnatqqONsov8yjeuRK
5TkySqs5LxD9aU67fz514WMmWCObzGwiL5/m5sXHBK6VjvX0mEbjdXn6nsWE+9zHXvZ9uGP0mqAl
5X5SXswdpkZ20OT+uv3uIj1NFJ69vr2s0K46GXUbJ0QyqhNQB4vzWOoBINpt6mjeVyPXqP+L9kj5
Y0eXHtDuzjFFbwTLRHXHlUz17pxJ7u7gmaT+/RSxLDH4yfCnbfabOtXzQatcyLQs+hI6QSYKAQPz
ijNWe3aG5cmYiJJX7FtLHm2BUKZm+VCaoNUGM+59biGowIPbBNhfc2ru2tVlEReKEqinpY+uXNPW
RUWudmWLOuWgma8uzRxUVmPQEcIkay39CvfuOBcwIhvJ01+XRg4qIjL/CsHlKxeFc98N/s6WjDqK
sqMPgQ+iJtReYVC1Rpv6iLqkQ8C2eWwNRgSdM00v7szfddLq/CxNMrYhYGbktkh79Xs09F0g30Ft
60Khc8ThAwj/lNYDw//dZodtttqLF/Z5kG6OYpwBArUJ7q2sG9HDxiL8OPaH0PyyaBwHr7eov1br
aTnuL2ar0pqI4uQUYMMScGdBp1sCvUYitgsr1zO0/HstRfchMnWsIZhjILQHIM361C1hYLE29m+9
vfUh9EhpQZxjw4pXHQx1nRjBL5cHe2jiJhGEExQTyG4HPk6mVBxZjctNYwLzwVaNWNCf2qPGMK6Q
JsLQfY5PXzMEVfOn0UaIpjdWmyV5kGModlDQD11BVnlAiWvKVLSU+2vYDtFcBUoA3OOw8vS9kgMt
fq2V44UI5JuVjkQ1W834HHLMIwbuUHVvSC31g6Fl/qYAgUhV8ZjnSYhP1o4pCQqBvNM0kTmOy+wC
mpeSZmwmviexcHOADI0KYGlR4GHseufFo+KQ7wX1jkp+4NXmRWyjQp9qLiSVNDh+7U2Z+H1tNwIt
Yyvb8DZHYgqnNuHXys5rz/MUTtXuhdOCBnVpvkDXrwl7k2kb+fUC0Ia5rJrXRxG8qByZTHmHMVcC
6vfInmOp+y+TOudJT6GG05/D+/9yWgjbiIqH3ustYOD+dH0rOkqsRjab8qQ5sl63l0sHNZWwB6ud
f5oUQ7dCGqmx6TWXkR8WNnq3INGPlmDSJgxIWUdZX2kRGxDOgJsTRR7uiPY3xa7opTRssUk1ynxv
shWkxttPkHERXGznvmbGMw0pf4aSadaPraoVhBmtrBxRuhSfcrkXrgwKruuYCx1qSTE8VOPNtC4E
Xjv88+SQotmzpdkfdGJq3VroUQ3kuDeLnXqHZHiDlDYnstGLcKY4DFCu9PAHFz8YZQQwBP81A3sF
28wr4aOHG+Qv7uSGGIENFet6yzNnqOL0UU5WNHNagcd2rSxHO+vnxOnKTH6G9eMH3B++KjGghshy
JBjnGYdqJw2dQDEs1jcv38IIE349JvRWl0N2Uw+jsOpojq6GYAbwLJTyHty5irk0mdnhMLhv5cwg
PcFV8rt4Us0Q60YWI++TfRAVjkZ+GdgVa0Rshfxy2J/FbTzRACyAMnTeRXBpH8mxXiMjiAYvik5l
qIzEJ+OCNS5HdFAw0hA4ZkmRsNEn2YELwg5i4mJCcuqRkZ4CMa6aVcayB8xK3H3w6SmL0wCyft0y
XTJwPCjhApq2yXx5yrQ/F789CHu/0fzDFmPAgEOvqdjFdDsz8+RvkmDfKKXHXIWLd15HIO6J+wEp
04Sg9E4TdeGrfxgy907rriR9+wBc8h4fWNSEP39bvSVgSADOqIAuOnRKV74ivlwOZ2lRmU6+Lkpl
DjGdJWKXlVCH/5Rt7CVt+ZEOdewoSMFq7lHYM5NAo0WTWzZP7S+7cbhGvN8W5f7Ak0lrZc/UxnvM
0jYFBHzXyZMyBwBI066Xnlzv0JQpbm0CCfb3ERnu3Fe1APcdknd95fFra1m6+JF0Wjmub1EUjLa0
RCJuUkcrObSq6ltUdeeVJEAALhfF01VABsBDuW4pjuRdcInvJekL1oZTk/FbB9uh6ZmUc1/L6KjK
ESm0lF/XXhE7OewA4lySf/7730C+ks2PlI/m9x+OJD43XCXxOrTieJNvDRe5BJOtG7hUAmPBpfM3
P8DjweoPUM08vDMuA4F/Ig+FxIsYBYo20sFNtAihamROV/c/U60kzpoSNa8HdHqgK7PxMR6i+wEd
DETR3SvrJoJmslNmjKHOGEOhThVFjPs4OCTYRJ21TWjwE127d97N3GnIG9c6ckmtROkUbwm6sIX+
5i90ZN0H0zZv7iJkG0IZRqzzOBbttpmcfc7TBqvV2TM07/X7lpnkGU57+Kgkrzz6wRGeBs9OmjYO
jxCnHmsVuM6aTLdBwcM0nCjQaCDqz413qurlekzPrDScWvRqGOyFp8RxgCUCOPwg6UT73qFpM6O6
50cFYPhIVPH/3rEYkoOQnAbUJSRbvTCODPK2gbwLwZa6JnAegIkDWTnNFWjMzUvESWICr3InbKB6
7WkyoRC3+9LhECpzobnT3O0pAcpbkLw0339yyrjCGCPwuG51yVosaXW1ZZsOU1ADFZ9aLVVu6oN3
1HXXwtc+JsLtzBVzAv+pqfbVncGxfN+vSOIMtjSO9DMVnAojwihWshPRsm1wj8KtwTc6XsRtjvx2
Fc+0mII80pE60gfWmqRT/GANxKeY4uy5j5obYzK/plegnIJjh/CQzGmkh2/0s4utZjT0LTnACxon
pqW2J18YFhC2dYUsvyyr8aRWhmyGxvEy2LEBoOC2GZosPCbXuS27czNmypM3WCH13jSWHE8kO75s
AfgsfBclsr+yHcD/Dxihrai+DVKfCN5rIolcndZmQytbDSM6ljDSR9cHdlakzz5q4tDrk+SRUAyM
vJO6ntw0Zud89vaGXO/1y1A1wEYWQxedZadbtHSDd6yfyWfCS3WgUnRO0bGUzxu0D0bZjKQos4Y3
1LVWyD1YJpXOuvcAmmLqkLq0gBQF91hVe8Lz1xYfGXgFhYjcYVsrrioDrF2LKqdj8/SxFbbfK+uj
OYuM6B5I8OkYAxcXxfgfvtS40iCjYpyqKZDth4c/epkmLp6hoXDLRz5z/xrxu0g1DPpiLr7HHczF
NmksSrcDBZOSxRMT/dq8meisQk7eWJ9yF4EcoEz166g5rjhyc3ENMsufUGrr/FjO/1v2Vz31Jx2+
0cDFyD8CflWEbGvgcxbY9+oXL0zPoAuNiuKa+nDPaLSoE7XtKu0m9E9rKXfJDkz+6PaGo5Uzeshu
+znUy0U48oJ1CuRNJ2scNuDGlvtVLSWemttWSpmi2HyGuOjcBqBnnbj35iLeyVe8UKm6VXiF7MXE
6ivYVTtXGJEOJ9pePZc5CuiFKDKSrDqhdRTGAT7yx6faxdPTXabSWr3vqjeff5GRzwqV7OtZW2I8
zINhXnZeGSLlo0fzaBXBVKvBOMQ7uwqoa3FSZaJfa96RXGP+N9Vd1R78lCxCfZhfH0yF2j+HjRdw
Ocrinrv+mQhvLgII07CvGLii9dahB2/QvYCxrXeYfqNRdffNP0Czp2nGxW75DKirqnue7aDk/fRU
JlwDcz5TZWYfCZAaKbW+eL5JWSu2yE0OWsDy/c/t4sIqDsTyNYLuMxfzFms9FaxhBOfURU0J/45/
zNFL3V3zmusKXwScZhpEMAnggh9cRheXwWRBCzDgJy5y2hdlsUwa8NmT+Y6ryvnsSsRm8/fnJ540
jmMO2JRfDFfNa6L/VUwU2R4psOgH0YOnzYA00+UAqSa3f6J74f7KbkJKrc9axjU1JptBvznKgqLF
qbIhUOAXFhXwNxRry+iPlvYcn+XHuRf8BCywfcrzzJS1zmCpjbP1rof8j5Qzd2BqzNh2gfeP6Ig/
7BY2FJNWLAirgnWo25qWT2HNaOidMzrOAVCsB5TH3EHK/Cz1/pJgd3RVXQp0fbdaZlvUZdCq7c7b
QnXbro/0IEyT13H8SF4PbBjXr7bbKwyGjV7jHpQYyH/qiOQDYxJL+fwE0oMFmrIystWc0a5Fx0YL
H2VIv4M/8q9lRZ1A4lNxGrkGvd549b8FIasSw9wFy18CeidvuzWes+rBvYQbOuw9IV0MTY1b15d1
JP3xSPWZQn3NlTYzN2BI9wYgBevLe7MW/jn5zzJnPEGo2fFnXEDNj9nCrIF7ycyLuAVgE0tUoFgj
LfsexfsUWEdTI95gwUmnpLao+aHQ+jOlWNgQRiaqsuVwzcntpuxRV3R8nNO0c01Hs8aU+R6tYVDg
HRh6T0MGSAZwEm7HR0CoLjHoTBXTTYTKhKZgCV9jQMokI3F7rgBrIGnG1oj0cJFIQQ/wK+fc0pAG
AamYYDpgetm8TeF0alnF/FOboAKprRmjjt+yglPsgQu25cF3kUQesh5WHVFY/Cv4lKxHe35q8L4j
Yq+0fUI6JWTKx4vAx8woFYJDo/uKfGW7K3r03dnu6p4hwcRGlxpHAQgxriTCKM1Q/XRvC9cK9w7N
SV71ABPySUG9CmdD48REM2I5LZAc3r6hPP/m7EQT5ZY4vmlK7M00VhfOYkihnajpI9ifIug6pYog
i/knnFUto11ZF48raotvzyRqnFLcjIm1syiYrLkH0N0YGHvg+kHg40Unk3+fmrFhxqK+IqQqNsFO
zuXPU+zmDeGqCvw+7xaYCO+yxpouXZ0Sh91bhx0FgKs8VxYQPl8/yS8ZIMgt9XWSPxTXwZwO+H+D
Gq0OZ8Vaf1SQmxpH4hapFtjSSzIDv3rh0BRk9TN1mRXmSbNG5TdieIOVtABvCPU0H4ITdW/xOqKk
Grus8jfxr3OPb3EDMrLaI0DLgLxYfkT7cpqIjSHRwpLXCBeLbHdX60Tr4d9HBpGi5rqqI0vv0tNP
LNMj9ToepPBA1dwdcrklqMvclHdFiLcPMSLUn831UHuY29wDLdVOnfdpuqYVaSXlLeAFii9Tn0iW
ZDnS8uJ0ggwYGs4NneDYoNSTXzfQJbkEqAuzqaD4o9I8suCbNwjXHKkSbKgYiiMBiLmDfryF1PHn
bakMVFypehK/bOqo35wFFHkGv2pUVHPsJ08GY0+zC3v/8IgHANUtI2B2S+pFXRJYSAS+ikgnx/WD
q+UajDabli5qbCaM3CqJIvQzTAHMFzO1n7pNDq45X250Ip7ABDrNajnt6yE7WsDeOiR6KZ5+GXS+
6Qwq2H7Rt4rmgpgwr+rwSDH+O8NbVJO8nrkYFS70JR+GyysPdZsZxd7kLRmc3qNKnL0GgrMl7R7j
GGXUrqFbHEFEgi48n6qe4HeDWfb2o+GAtqcLVGbMpnTptg2j2oQlPc/TBUtbB6L/+r2qNcIFZOpI
fCAZ1Nbxg6+wAb6qd7fTpe7fuWpIOXD+UPkX3vQGxnW5cmrGrBQfCGfwQxR6SDqt0MYVl1py39Zw
DwrojSssxkt0YhBqLFMkWPIhG/yrKiVPD/DeNzSpDLmSzpuzGB4NvRcZAkXt6jUu/IADc2zw7KEp
Y144021LTZt1aErqlYulKLc1jnrUYvGKekxrRq/VK1cdQj6L94KTAT7p7lYaWoa+l+qDPrI3Q/7L
JUm4ce1vhaQP0YzzHTPWLoCwBcco/VGCHAp+EVztW8SRW6NiFTTIotWPU+JgoHBuzx/aTDNz/J0o
Y9dPsxI/R4ApnASK5C+RotRUJwcBLNnwX8Utay/PzisVPIqN7VbTW4t1AxquY/czyis7UH9/ggTx
FbDB7I+3X53QDSfaymgT40cRVjrTSX+MoA9ygrxeLWkIbtZ4p8YJiL74txltXVpBt8LR7GGbzutx
AFygkWlorVvBzYotTJ2zdpXTF+3an9V+aL6lua9e4N17IKmo/eNKorBUuHTHeEnwpe33ahI7F3EG
NskmSu3sOqT4bOw1VOLY/vZw8KQUsvLjWM19hRjaIneVtdzZoZRCRmfR0XshN1Y6yL1cqMXmEmIk
h9OSUSUl7+FPLbZ49XDglnWKvbDeiNYD1rx4f7dukzzlikc/0DUiADw5xxZRlAb3TMTEuy/V7TtK
Due7Zk0OId74kepCWKWSs0L404SSU71MaPp4Ncf/tmKDlCZvqVtzy512rNtoY5HlNEch6J6bs6eX
XLwJ/TRLXDGrsUKyH01TumwhF+GAo0WFvkzBubMuxFYW0QD7tbI+RU8pgch8FnG2FGa1qiOEPrkD
o+1nJd+0btrPRic30gF3y+99b6FUq2RTCG68X7Xdo2cRL5qwICnZLchjWCzXu5LQouR8mL4V0drf
yUA1rydMohcquu1xmGMuxnxFfF5IxwMOZ+9VCYsN3lfvbweaYoQjJZx78hOan26/7LV2Sh4O6jVn
2qqVQbT+ceZKjqKftGBMGTeu5/yXmQ11Jn0PrX0P5H3r6XgN33F2UjmJxdxGAcbA00uGuyWQYt70
anS7GnBbFh8PDZoCNSrmr4v2Aa89uY5t5CFo4F5o7/D6G3UcYnk3GwzvRiaT1So3ONIdhOYWFQ3p
4+jKyeuXEP9QlJGuL+IZ9D40d45mSiWnEsJPnqFcOWZAQFcUd4Y6xQ/e2nDYHJugTJXp6gdfEda5
SvfmqMD3csknFxOX8R19DZbjE4GmgN66tH4uBMyKJADKrX3DkT4kbzlfxnd3mDwtHgOJz0YkRnu4
PAa9Oy5vsL0+8tV3BIaSEUNUnFtOnPnCGjZPm/C31aKPYYJUpgpzf3n91yZQSWXv1pGhPa7q50v8
/TeOBveIWLt3YXyOnkanFpY0AuqiHRdR3D68DnJe9HFWZRvuGCqvyMgT3yTZFmS9JQE1lyBckG1E
l/LaVOKJSEAhB0aXIMPo39nExa981SLfPFbxF5Z+22WsLrZhbIUPiayg17EHFRWmfq0PZBUZLEkC
lkExwtTwPEE49fYBLkyqavbbYxc0IqjgfFcBWuQuDsu4jqoB+ndUtWXRYFJ3yUr9VbjVsMY8SqOh
CBOBfusl/PEwfO6eKMkgi967rjMy9v8LF9BbSfKGczA+au4KTwRH9fb0AsBaXVUApb4GYBAW2ZGV
m6E0J0o+McXcrdIm1Xhl+vStYwtAKYtkAu0UzjKNwiuyD8A9xNTmbPJBZpdRlzOSBqBa4O7s+wPq
YxsDyT8rZBYTqLNhyP5i2LWcRDkPJgJJKH9YbcWL37rVLYYQZ2HSufu8rp7B+QLmVesXOs8WMFWX
hHvHiUEN14h666lnCFoOAECyGOwSFgce6D58lPZPV72ci+swL7r9cZwhh58wGwxUWkvvGMgQPBEj
W1GijqTGUv3lkllT2yJ/hpunr1BMU/2uebnMdu63VnX5md3Z8tZMph+BdAHC24UATliyOlO0XNTU
1AaBaF3k3mW9oQq7ilczeZdbNNhRo0mLZQaHrjxJzDEJ7wR64ilRd2VrtpBBu0r1VDQuubGoye/l
RuJ0jIQq7zFJ7TLY0kkPOhsISmtPa7h8bSH+3HDZBKdUKwxphY6w23jA9zXrRqOM/a0mfcsSsGep
pKljGSjDzqL6Pq6V06mEP4HxzpFEEPwoxBli3njVwGwyTtERYmlgkwpgZsgoEjtiUQdmNDX+yb5U
93q6ElTbvEGWCndmC4XUFqNMMBzX59TTD5KF+av8ZDgNYdb6j0DaQOTptRi1+PuymGiG63yuzHKk
nhqUVNUlqkRZy9W2vYXWsx+NMqDce8GpOtW0101uUVBnq52zhD/arFMeexVU0KwXLU1abfsGyu3c
Ty1dJ6Pn3kMebgo/BWTka7dS+QLu92n9y+3212+pCGJ7ngXCd+bXnRtkaUj3DA+9bLC29ElmF1c3
YPxiZfJuF2XvVLyi3/HawYi4XW8InDvF9lC8S2xHdCBb65JkyvrpdoYPvqub1yWi906q8L6XNfAe
Gf378HKOPVurS2Kl+3Qyim5APWQh9rsUEnu0XAnJ2wDTh3TlHHLRnILmQOyD/MlCf9rN76svz0MV
h6XZJjwc19sYMjxrsb7Bx1DvYR2qwFgeSSjm6S5MlfVN8nnoVKewHnrJynoUm6JgfLrQfUUPEkhH
QYWAfLw8hoc7NQFDui4XGTtHGZKf++vzp39sYRe2xvgt/aHDTjtSdKNnG4qb6S5Dq2u4rJZxA6yp
zSP1OUuaQMU1sSY+gFVjHy0sF8gkq8mXWs9mOMJrmEmIw6fCKQ/mkwQC5XjdJi/FJpJ6ZO0rueAN
4Bcu8+pzOtTzBHxSC55Iz0zLIcujSnKsGhbeKeyC0qji4ohrJnGFxfhvF+hxJO0kDeGUHL0U6Vx9
6peFV9rMpO9QchgII+Jsyzk9Z+tKfU5ihfDowYJmnk/t4ZGe98PtlQbbS6B92ZBZHxTDlwYN4uhs
lX5E2fyfW+lxvyKlCDHHFEdj4ta1VX9vElerIFZ2/VIkSJyFVmsojnU32jpzSEyMeR8gtyXjdZKb
VkIq6a8nVIMHm+DGQ1+/ULDTuK7TVJXNFvsPtMjhXeW3AG2Hwxdx5mBx00zlbR5iZzlIL49vTfHC
eTBwDE9kQq0MUw1JRlSXDjI/ro7BIoCt621uziNgZRqetXeH3SBoJsahRuCRm5MHSXBdeWmudQHm
Z4gCeKmDxqTbB0uazpIad0okB786LlW7CHOp2T+dmhw6M7QkCFStS06JhYKuSdDdXiwAjBtq3EjX
u5z0m8K5DwasOqxpIpyrrvaTPxAf3SzpEBexs2vg8xA4fxIQXyuskwhM43JkuSz9asLMhSZzGgoq
xeXESlsRpZML0ZdXtYBcZC9U4WAnStsETPdOsZTd9qtzp7FCauwwHScOZo3XHgQZjoNcFiiXB3zR
WvOCQVxuwRE9TgYXyI+wp/TEgeJ/ENecUFE4TRDii8VIoqePHwY3o6+7FLxL8tJsSoCpEYBu4pW9
Hp2056ixFJGsVQqV+AMVJTX2VWdq6gybzZZBzTslsuLMj0+OqqZgQTPFd6apzUBFLJo4EdjhBl/B
eT8GZxuX54Dk2aRrajGWIB9xBD7RcReUnDdxNkMa4Eb3R7qh1SgMvRdhb/cM+9QXEH239PK5dufq
CE2xZe5u/gzIiopL2QW0DvZeat9cOFczKRkdYtapcA85wErC69fswhIJQW8C6y0OnGoisdnMPmhd
pSz6vKgbPV+VQfIx+6dZ5Glswter1/SSocDuhnxBZ+zS7S747GMsGbWnadAU0iV1yMhRdM/M/vtz
7FuSALJ0DOdyQSc+MAENPny5Jsj1bg8waUqouCyaO2kBfKfWiVw6tSG3blp91EQLndoM8rvll4yi
uQZBblPqyJ6PwVow5NaEEbv7ocnJ52Xowwod1yS3NMvBOhAGd4IRHnn8XTDTGd3ZxgdFMO/gIpkB
5sy2DVjp39/lsK+36qnDnW7Ysh4MSRsLemHHACtgjHOvTlJIs8X4KUc4HPnHUeYonmk6vPqq4Gxr
JIZLoMVoFkJFYjf0dDKyrSrLc0ccLq+/vIoDK2ePY6Vm64cj1skiKXlh4NvipomzAfz7BaNGZVFh
tBvLvGmDDbLMyjQT4t5iqa7LnaFMll6GGnYthPHS1gNL0nzzE9sMzF+XJGUGmCt43tRAdMBBuZkH
kfuUvWMuxdV48C5E2hPgfIGGL0DO9Php5sIgYYgKQPjTQKQl6erxV/0eemuQIZ0tJUWPeDacejYe
zHDJNbqg7PO3VuRnBS9zN6nj81YXNb+HLVv9XXv6VRI8w0/EHCaT5rnQma/LA/qlaYtpT6AKRpld
oAwX/65vUNtH+ZctUK/uk4N/2z+96+0qJJoKrRqJEWOSp6brGr666pW+zgsHzyZlVNhtKAVNWqyQ
+g10CSa2K61zdcYnzoJ7aqxtY8uDUfupOr6UcTMHfnV5SwEHu/PTQYmq40cwyyAeJQf45mAPS4Py
eMlh7OaR361aYAdPCjc7I/hxCuVhczVy3dRC8T7aBhh0IKDcCxl6WaW0WhT6d6PzIP1lmOp+d7wy
BuOJ/ukw4gL9+y2ekL9EPsRBSoOQsugzeMxJfGDXKSI2xosWZisHvaGLZl4lHG0Lg0kJJ7rwfO3V
XWhdTY59nH3XZR2d3m2FYATfgG6uQ7LIMde7g+cfeNYFj+MBkwFaspjyp6iSN5uLB/uNK/bMS/OQ
PWrLGJE5tHSU+nLwSx/+V0bwyET7WIXk+UVrtiIjUaninyQnFv+b/ZBRXqLYmVI29PMXyOudATfS
mumnxpuiBOQPcOdVLj8zKNczKlZ4ykZBN+BRv2iOhqelfw5Jll9XJgqABfgWqT/nGuQsgvduGM53
IWpBO9MPLjBUGtIUzIM3w5pssbMGzqH83tAPzTGDIiXI1rBeTK9qM2w7olhTZSutHVoT3wx+42F9
xEs/ZsfGf3SlcfAQu6l+fEuJhzsOGSOJryJUyL6mve0BAnb3rgnkEpsd8MyFUobqMMZ3HL4bn6SF
ufWHMlvZrADSk1zRoGSRDK2XG9p0V+FuHJayddGFZKrk+7G8dcslJhtBGol+1xXopxDjaC8S1k36
bil0qx8bsp2Tm5gGmO2VEkVrKd4z2sPykjjYeNzYXrbKEuwhr+vvE8VhY1qfsbkZC+y6je5nKdvq
TnOLc31kwOV2URwnDmFIK6oB7Mz4hv6jr1Gtq9Uyu9Jsd61rovbDd3LuoKJJLZz0Bhq0b8d2yCLl
sG8HOiWF6/b75RZXlC+69viP6WXzC8UaEZXDggWtOCXr70kUQMVk1qXWYF62qQ6fU1Dn9dpntJoG
uqq/mwe/6Q5sACY1nnhn3XJRSjnm7kQ0x6VC40TtfPVkxs0eNaj4lLmyAiDf3QaHIssiwo5SvI5Z
ER5hSNvu2kIXEMnhQNpl3vGt3qsPX/CWfKSsGSp5uilZ5uQg3UI3pQ7eTmlzHGFy9lhCnLBVDrmj
/kVhd/qftQGEg1VkkLdWbbBqdQLMRR3NuvKYxm9hV0YJaQ7WHCtlBoDIoaXdmLPefJyw3sdmI3bU
z66xrQQen/hwEbyyDPgu/FtGxsVzonybcyGq15OuS0AWfxqboZPfjTGYZWeHft/ZJ3qvOA6baDmT
5BRQMcoYk80p+a/xn1yR1jYfBtaY5L1dMhYn+QGN6Z/k31xXTkaxAnN0mdYmMFsm3EZkqJQF6+NH
htDVIVagKvAg3xrB+4cWZECc6xmHhT9bG6wFTSlJWAea+yAORltJDXo+dcOVncYoOQBOxOiixKLz
K5zkR1KglPh4jI8gyCb/PRmA3lOTdhONKHhrpsjn6W+YvKtQ6BI23gAIQj6+lyJpwKQ5Uh/hJILh
6NqnahPmwyNLin+VofH1jXGHCL7gFIBPPFoO887mF1WB8cJIzHWiLMe9p8pbIWRBtjhASRqLDTJ9
akFz5qRQ7tCZpWZogodI5hXotuaWyX2QKVfzRH/JNnfTtUo70A/dhOYzHbO7RL2cg85T+UayoBse
jg2OiPpoMLnDSCVUFnDaaaJy6lOdSiu62pgqjbB/8OvdDjXFOkbF/7OKNAF5T8V3K0cZzO05PIMd
P4AaYRDeSpMNBtRoGTQPqb9GSopz+u4XlOMRlnL/19A5GAzMggRdRg8a0CsB1U8shsPoFXihiI4T
GJrVUgduW4avcqInxyr/EC7Ty6aj/qK6Xk1WUQkeUPUMhwoSVG5gu5cDilr9P3QGz13WPvSVbWhc
iw6mybDdg/qswAtNmi+lOAUynqdvK9GNyHqUbb6yRIBo+BZqMZAXCvT5sPfSUb1FSgo8rjMoQ7t5
TUWyoAKJQSXAvzweDajycYCdITwK7gUBOj3WelGGVPXmFS7ftoKJ1qIwskavf+SXityx7/fy+hPA
PFb/iTss+bUPxsvrjMlmvxVsty5/mp+0OrdFAnrGHFpZted+YVWT2f3xFZVfa5UqPV/W7NcJBtzO
b9jUT0PtM/0e6J5z5TYqQ46nOmx7sqTY5v39Zu+pAjkPw0W2IkQjFouApycOMb40Wuy6wN0Q4eGR
Q6muCTHwLSCGx8j0+PbzqmTj+Di3KOH/K3lJq4zd5ye0GKJZK3vG3qbxpZT2cbfRAt2iEPh5kIgH
dCTmm0cjeGPo91qkDuzFtWJ1NIBhWkbvtWIRaflVthXNr26hvn3dDZwKls6rmjH9UvksSYhsMmKx
l69LOlYWTEXTnp/VRKSpiXWYvKgxUwVlkCOKQPHe8GFpFEUXnX8MrlJrHhrRYVt7ydsT2i0d2jfR
Im4ovghyhh5P87+v15knkB1kwAMZIrLVrzpAkDYY54iUIauoMrfEnyv8Cy5nGKVr6zbE3Uv/637+
kbd5RDPdEa79GLSRA4kZaq4MgENyuEWQCj2uyHO0Lf8cVIEKrBdn7wF6VoNtsezOn+mv57YEabCW
mF8XC9yJB59x1czMYQPKDGDCVJGy3wj06SDmrfMx7FVcjwmUni52AFEIZESOZ8bppZQl9X2fmLS0
Sckoa9JkGu7BFf29b/wROVdmHAQILboEzaFHynbK7Jg9Fim8/Cbe7XBRet3yGipfcsCnt3wLh5RS
bh0ivkx0qO3dYqsLyYy0gBeclN+c8Um7t0JraI0ZzsDUrzRk/+YAwhbR7APhwugIGZw2iJH8DNmD
Sxb6skn0LJ1lLMK1ZlsfaJ2ZxyOqL6htJ5UfdC6dT1AwmujFUFksAUXZakCfwO2pqdChLLuoEUyP
AOETuZ8IONTRJX921xD49rxgVAwNGH57certDiC565f9JLsxWILi+s+04hxOr+XI6GcedVDvmqKv
ZDgqF5TZaGsf54XTUgIBBJ4tvBjdchLXZUsq/lRapRGPoPVQC12P7XOUC93ijix1kqgwCzhOSFLX
m34v1Tiwjmv+vHKfWbLT6Qbe23jADRlC2imBA/Emp2EvCwGcT8m5onuC3+57ogwLM+uRJN1QOWzP
Gi6ltJVnt4OpxMp0+7rb1lyIHzCkM5/B4BgyNjUoJx5fqaMiQiZ+wSJBAMxcAwtz2Uc+UA/nPCt5
97M3Zk4QI3tBImDPV0enAERcU9UrrZSagIPvoQPub6irsCtT6ErHAu42tb5HUptYET1Vf0WcoMr2
/2wTtWhP4vEW5ZI95Cjoj8JEw6ielrYtaE5knbnIfTgN8XqcT5Kl8MLKMl+zh9yIsquuQKrmx6GH
TUrLzxLvhFsnVDE2lon7CIUDgXxpu5/BehHuXLwKfsgWqgeRcYdztEFjiDt+UKlVeMaDKsPQ3yAa
9/dd2hNg6Rqx+LAQNEej5Fbe2Iz4q+T/crZ4I5mi3v6h7nNWmclnBHBFzZhcH9lrAMnD97TkTsty
l1AervkjasG50ZAgU7mMN2QCbelDVH4m0Fd77qzMIrROB32SeYvxZEvlYZhQTVquVUhpfjxSg2Xa
TFlp21PD9D6RdHQlWxIZOKLHV5RiFb13ATehnFYw2We7iUhH4BS778+ZSXdQ6haX6uJ0z8GpNYwf
hF1l/3yaTf6PRT9hMhJm+hPS24EcZZW7o+OA7E/F/IKkKh+ILLOzRpnHPLWyRWomyEQJecVSTXAu
O9zSIb9u4n1EodgmfVjK9SlNTxpejEl6j6y5qgjdNnVfomD+YIYr4S7Lj+bsE/blxitOdv/la65L
6bL9ZYxF49AwChdwzWtJvo6bzjkHE36oLu+oVyVac6gFI0+FKHlQz+YNUYOWqpGqzeB7xn5bthh3
W5k/2kM/F+By8aXlcJRrP1rI0FlkgYXJah8WR0qNwwgnMVsMFijfY2OHMwoJtaV6kjI18AZaYwRN
k+1vrlBFS10fETYRQQPrONooIxUkgTTLHP7KgvhR/yic1QnX0luGuP+NqzsK3tTx0MFpcyVlaU8r
FOkx0scHBYB4PeoED50CK97fkh+7dgyf0muBUH3I7KrKygqqekR+btqFGw2sLK/PWTKsXGinn6Ja
4qLiW8ZPU1rWVwQYwFlMKvW10C46TEhkXjj63Kccrn6t/u6hdmfXt0MSDov33ilpKdxEQmujMpnY
moeAxd2lZdWQu4aNfAgyDTOe4WHdSIjhFbayfza4GvgrA9//nVYPGr9SMopdTrtwkWRgT6NHlO1S
CtR9SdnPwe1ffk3qKk9r6rkGsPiy3Vza6g1oK0pnCZpQxdy6Eb65SoYCvvTFYDFIlbMX9TVQ/aQS
wTiWd0ZeEfYeNzRPmPyn7XLG65LBO93Hkqt3kZ/kkNmlfNPZEoPtwhZNL9s22Pd4HfAHtnKccW5k
r4I4uZ26zwef0JObIPPflitsCaaPWxHa9IMa49Q08l/1lj4Kl0w7YY/WPWS4WYchN+QM1ew+O31L
PhVqo0TMjRF8VyQOuyD6fyYamY9c8aPQjc+0A7+3EvOvipBi16K4fc5FYXU26wE/uorcFbqo04kf
Ek9Eo/MsTkxqxlW3u5XhDyHpuhr01C/IeAY50IHlTnd4iMa3nL9p4ba7OFUQoE2IGtwG/bkq9t2k
Gq85x30VHRmJ09W7EgA1haR2zFBRF58euf48zR1770ZYdIcBVdZ6fL3cUeg0wsbvLY8L0Vg1Py54
RJhL6HlJPiUhMP8yJt5Syg7ez8BJX6RcwrkvHfGdYX9N0EWQij0LYvFNBfnJzJKmj3X3W1Jf9UZa
fYMM0jNF8oKZgNsa6vJomfzVhKN6bSlyxmguPo1mcc83klVzUBKVZDkEXhzuO83zs0hszM03jDfh
FHuVl9jV2kV+93mdggPMn5jTmxs2nFF8XwvOda/9U6OiKMx4KGbr+2d+unpzh9YlMETqLX1iDiOS
tX5KqFNfN612MaA6HV71BDYKbCv0rMPXrCbdjFcc3LpNLceWBFyG5+F6/v45rj9bqKmNNuWrGES6
DF1qWD/hBPKhfXzbqXjD7S54p+/jddWjsjqhko8Q905xUNdYYv8DF88rav/UV/ORDgj6mkiUIFmM
z5YdRUjaxsnes2s7g4G0CNEAFHNWheqY7vrmY6fJLGrWIKtyTSfvxxuV2NpZMDfRbu6XMYMl0TDP
+hsQUaC8SfH0cd8eID+LLGdk5ELfLQ5sZ0NNDXXDL8xJumoiokxSObZRCmvWHchh+C3ebbzy6YDd
XxLKTynbdaF+GEW49At73vjv7wPHKpN3kupHnvC7zduJhEQNDtma/dKMsA0COq48XtSy2wAPG100
TTsyhrLIifLoekSwZ1poWSMFcJ4sphrP0bCbjCn+xzX30AQPc8XamVjcVoAe82Gva6nH8d/L2/Wn
iwEo6CpMBDcSaTRVIiVl8J+8F0DzjB5SNRv7wtBxkznUP0m3jkeX1HshHxKINyqvj83cXMyRH/bz
zFeccVpB7N20Oc6OhoJBHG3JDAEWLaK7hLGSBCMNpdXDUlRG1YN/7PFGj4SnTijpdhSCjeG6lXIK
kHQ3WJ2hvrVuqz2ju/jMLvQqrXd8NjWICgMdTxGAXcxgvm/+1/QVLWnumYrrl/g0Xb73qJAUR6oQ
7Z89iWIpPZLUmoBC8l4x6Swrs0zd+WBQwzhhmD7Pf69Bf+t4LI6rwh0zii9lTjuNHAEaW0oyxM7S
zH8Lg+CqAUJkwwgWgSQnFpFocr8sB2679lH999l5p9yb+KT/S8yST1B2DfSPTaW90uGArviVe9UF
O+8lEJapDNiDlf3fqx0XzGbvnomlFTThfUXsfpi0mQVVMLLUkeUmaS+hJmF0exU8LKe46f5sqRCH
IVmlcf6IuFciQUgpNacJQmjwBqvbrnB/7EfRIz7T0OhnFmLsrkGME7XAIhHy1qbNWHGdBSnv96s1
PoN/WE5ds2/lr9LNwJc2/GJ/YLJdqXhWGrMbpU8bhUI+2zx6GrzXqlE9nQk5qUasVoc0Kid6mupV
aDX92WsF27YyKz8KRswsH+mQYVVqk9ZuobZ2N26rXzDQHq4jExccULDLRianqn85raH0XnZRzoz1
MRwmsPKz3PDCnT6pJj4WoTv12LOaFW3CzHtoJIWRYi5FfEe3a49MGq2KSFHh1cV4KJNsEqEGFqPb
bNY8kEtqRDR7FvO8bwGodE6Vw+fnIKkaw3JEWNrPzSLeZXavHQ+txYu6z/dt1jYo1CtJVwGxNz3Y
MHR/erIT+9TF2N4u1oVVbBW4PvDaqim1fqePpbVZ1xhpP9ikDc5Z5kQHPMEW2d+GG1Gg5QYV1wQv
Nlo3a3LItmQTic8KNgbeYQrdIbCd42eiRutamKKN5dUjeBispfWVFh7Si8nfpeU9m6orMcPJ+Qnj
KNuwAGvlhCbxlsO8J5DFwhF0Y7i8zpal57mJnpd1w7HVKXAYLBdX3pE04TcuEiL76UH5K0ohSQCy
fMIgFxYDQpmcUY48ADSI4UKBjlQbHsyqKORANqY9aUjq45YRT1FKX9ejA73qgELg8qvsjoK9QASM
zhE00jQj+lsKlU3X+U3wuDerL2s1cmeXyShDkE/u+2yi4BNHIYmQJMYjlAU4iVT1jX5oX/1iltfM
VosOmk7V/YC3BEuocHgcxhP0+sE6GqgSbvvvsS3PqozlDCKs46Oh65JntfJ0Nn+6vHQN/YOMVeWI
G/bzbx4HuYc78DAxFTyo1vnuon9QyClheVs5LIaf0n3u9PGDGYBgC2ZsvJ75g4K8Qp3iCWcZncc8
GCKGeJ+y9lxek3cJ94BqSpOog6Fg76OLqVh7b9MVRk+XzT+1g6sfIs9P3zHz2Pu/DxxEEPh7vo0y
vk+ts6FFhIlO9hSIn45GcWErQICEhGR/jy66LTBYu89876bO7CxRIEkprVat81QnSH8IcXVTiOZ1
pKqk3Dd9XaPNLNYxgxiyviFC7IJBiQrv0Q4F6y8/cFtNBH3y2t3SPuvActsswnEk9l5P53iN7hvC
9srXQT3U8OdpJAeWtMENZixpRGN/lY7WR1WEzGaaVNHTqgWpK+STBQfSgIVp92xhN6wGjQ+CRfLH
F3aINzv4JAiYlCBo6K4CO2qiJlPq7kbqeu2/P3NJb2NsHOpOZeMokUV8cN2sf7cc+XGAHCoj9lqr
7bKGJTvq7ju/aTbFnjGq/RqbpHvSD+tdqfVVtbXLAteY7IcotDiVRDDUoOzEPiDYKAiUplsxD9Mq
xaoe53CF5Wi1i2TkzCrwEFu34uS0h8Jbngg8n3EtiaV50T6jbVW5NFkRm2saCRMSbCaUOesMkRzF
IFAeAWWVptSXjS10MeLuQgiAFzrC3i85nLiKWyEz8vY6P6Dvbz5U6kb+vU4fxwkbTizPHpdRfIpM
fTpIlZOHyPty544c6J07tzknbeOSuYqto2IxguCndK0wpe5Gjqb2n4P4vOem8N4fdiNnRb5oVlo0
tyJUZJSfN8C0rwxg8ZdwhYpm9d7Adn3iXbjuqmL/AyIxz5cWxZBCuvRJSvW7Ews5juIHxJSD3fnD
+IVrgqBOhNL8jIUHTHDV+ehAorfQkfS2kF7km3KVf+5DkZMg4UMgKnYYjRgsuzNZpmg5FIbdEYAC
RaaqSXFhkyPvunYk2WPAJlJOBuhaiC/lGUyoEXVmL1gOmd6uqJUMBNqLW2fvTXsrFafmcLXhYPjP
eZ7Rll+KoDVqPv7Zhsq8jUKj5pMoyJnl1oD3eNq3EgD/vl7angmgiuCsPoKq6jTFyyNyQFqUhJT0
eCiCC7acPVcSfAwog40foiDovfaBxyxOCqYoHa5kmtLW5g2uRPwweDxf1Mq6NUteE+QH/vTVAY/E
hdbiFp0xksdFx96ttdu0ZxxmjclDg4Yowjk/el0Z2TdiSw8eAvsr4/kXhqPtZkTDH8a2XseJitN7
iCHfZsUeg48zsFJBQzEiqGMQHTzJg7uzrEbh13K6gANL6+smLG/bSXiUmeb619yrqQ4QzWH2jsX7
/+nEV7BIZbP7Fo6pjwo4yxPATbPwwHy5VQcfzyrfsilHhgFf0NU1HaAQ6svfa36F4hNozOZcWSXk
D8OvsWDk6qqETDVmKlJbTH1hr3VjE1KN/TNMofAMcEVA+tP5DhfWxG86iGHB8tmyOARcgX9U3gtL
yuLszXpC5hqs19MSdeHYIlAe4edjpldEGLXpEfEZpQH6CgaDp3E3gbuJyG44GyHwYl5AbHX808Wj
NY5YOrOXWiJbP5jkPkc//3CGAPV8OyktGr6fW4Q4pS8g/M16MfFyLlVa+I5/rJhJ385NhyUfYZkx
uHs9mmY51O4iCSlyfYO378Bv4AhVJm41lDCrLVWzI2ShWy8uzltsdq15bScY/zkA2q3VQYktvwmq
wE09T30ChWk3kHA/RBr84LwnYSj1HRYrBzqV556J/ScDwDklfdaISS84sM1iekFipSfJKE7nPqBr
2j1kw1x1cDawi7zRF9wVg253AwQxeo64uR9B3MU0AvtJYwPx4+r+qD73jVZJ0XQt8nCbY7fkk6tL
YkrgugPg6MEHsCDDOGQZlYxxnvFhc8OGcm/H6Iuuj1x9lomJJhSsW3wwPaJrKCXH49crYn/BQ1U2
EUJS6k38GT1rt3fOKuBGUfYhbvFd7UAIQJJmHuJn3AOkGDM5dWaIWFtXBe9GlnKJOXcKBIopBJCk
LfEFm4UAfS3mJjremBgGjdjSHqYf4IUfgrkYGmrr5IoAOQ/VakE6/Ev2dDS+g0qFC8rcwRmMXsFB
whsKqzV61kZQWQVi28FpTUkwv32yw8co2AET44SNBGFAaywRz0rRpHUkNDSV8oVDr/gKFkGI6X3N
WAXRB7S+0y1SPMyRteYgVaVtOIaIzc4v+BRHGZGhv1oqqSfGRXcmv/gmyxsFYSMPyt3fixaXDGqB
hO4nNWUnbx7wyhbZ0v8CI6KeYv0UPNnerWb0Iu9OqC5YwIZ49J3UTIPjINt9Ok3Tmul4vjeZ3pdr
qbVO5OjY7hbkFupzkQRfEqEMdZoH2xyAF0GYqpmQ7+GlqXJ4t3ClvfMTnyx4oN7r/ZI9nd6tureW
2BSxQwKfoWkicoRjNeY1AhJ+Y4jEBAjOJaLuPeYMqWzUtrjn4AP9ekvhnpaJ9+f3pT6gg0Oq24j5
Tfnz1f3s4yFNrHqefqIK9EgAzl9f8Qwy6xFxdfR8DdEpCQewnDYuwb3mGrEHi5tPiOBSHuc3RO6H
R0eorasrsHoeUS5nVMVhAOR3/j7IUCCvFuXpNTTNx90XpUQiJh3+8UVI6yy8mVUWHl38IihUaz94
X/o+S8Rmxc0SyEKj6St6qZKF2v9w0ozdcpyyPXZM36+6uxC8gUiN3cLDgV4r+Kb4vBCceLBxvrmv
i9xTiYJcJMiqMXOzMBs8KE7n8ffPv17d6MFwBH7auiZgAwZydD3xPoAOZPrxUcrd3SXNmg5DzFi6
GmWLHdGdrYvzW36Z8EjEooaY0SGSPFHV5gCaKbP6mlqpXdkqd13Scen7LAOBixVyV0bGBXAwqdHQ
NwgdYmpiL3bQGOQBcAa7xa1KqSjZg0TPpLlgwhwFOSBDuCtSN8Vw8KI/01BhWrXKDBDtHMzHWJqJ
uVGFSdebO4kiEAg+K0tYhJ0pJPelx6HUaznYA9q2gt9M1QZk5Gea822W1WkoiJCbtaRYuurOhfJj
icK7sfPWk5JMguIqCOCrlc0XPjouWUBooWop8P+z72rjwanI6jQ1FPparER2wcp81HCpP3/1XmlZ
blmIash3lkJiCvmquzj450xiZ8T6h67Pq2g0n+U3XeCZ39b/eohZkYhnWDR2tHosuuTB+VDfJNM+
CpohC8oUM/54AVzRMo+8l1qH6uh3txIQUvKU66V47IneOwbiedDFTulBAkEqNrXIymIXLrHfbq+t
n/KwsssRC5v0pdL0cTqjiWGO72hmWyKrPZU8mW4lJPSITlpGBW1I+0/z8n7n/mUHobU6pSHgf67S
kW2X8jnJwxlPrvhobioQPgn+IF266MCGulVUIQXCq3jVekkeUvYslaH0AE+xfFmZ82Ge3J/KCBet
SapeinEGX2HAlNUBcCs6bMyZHnhYeQ6ZiYdMhZeHXCflJW3hgV7Yxw+piQCUeuVoK/01scAxN0jl
U5u+aVHEN2lIjrOGD0jB8IzsEn944H0vjkqE2i+PaBSnC0T9VeSxtpxaNpbGNK/w7bF54zYm/EwJ
oqe5Q9XReN4Du52zDkLngak/A6rxoHsV45V7flDZsci5rL38NAuxR8bbPA0fOibCGGoBCceFU3bw
YIlPaZa3DPYjub2owIZ4IjQSqbvrCkoYaTVtYMeTUtV2SfVDVS23PI/UC/7sdd9DbopDOBeSzmLC
3WPJCZaoLgEyW/ziQaaa6Er5AHUqu31aPu7+OUNGElTWVxWvtj0zLzBHrZ63fhHctr67Cs3p7B4D
z6XuUVOvoW6hUEGshKwlLN4TasNeOzCQFnMB1BPf6eZnRYqkT1eYyoTosu7fx/qXu+0i/WolNV9h
X9BmpeoBh3FnZOLs2+APuICQuudhNYWe/bxMJomoxpdO1Ynsgh1ApLsNVSbG5sndDtEJOtkopFTN
VCx+zIpPT9VA8oSE44nB1qkIUT6OS2BjhNJZnps48W5NsrJw2Emf81uMl+V7cKMUqwqXamsdexpu
ptw+3UxjuBV6B0oXPw2ypUSg7l1h/uGmGr9OtCq3pWi1QUFP9ICEC1GQxFy0WphSuCggpUiZXbD4
dVUqHBvQaIUB9XtxbWW2g6nkTXJc2NgIEzkmmIYEJW3cnL91M3G999c5gUD79HIMGl2RmanornYD
EJjiWBc+woDs6CHZ16mL3NqFyJwHMJ5KE/YmPD96tgWAftP0ZIlEcRcfWdRgedzdEojfM9DVQN43
NW6TlwAwRUAhR4UHp3hsHgnkw8gpzBWs8Yd9YT3LrbTYFGSwD1BzbN5ipYKUDnD4eComBuNXbYhj
vGh5g++v/hFTcMgrPuAKFEtEHJirASbA24y12Mqt3uFXvAA1BbQ2Hg4Qq9rpxrxdPeEhVARmJwSl
FiyWiSyDmJlxXzY/7byTDrF5yHaQHoz4pbn943Ww+UlTkWR+s2JzpQ351SZvHUFliDJZ7VsdfRg7
7TOFsWIStxYlArJ+a7ro6QfmJ7a9R5YyVWOb0TMZsgDUzN2hgdkUWdysIlbsYq2vMNXxHZ33yVT8
6MfuhDVRAxfQOojdVBNcLJHUU4qDba8u4m1RNvEzfSmi0PgCW4IcU0JD5ene5+14rQNglVm+3oE2
DaRH/541sMSskgIzg6zyRG3sqk7QjQpfKczqYoQTvjDh3Rsb0uOLzSwkmEc9UtP5sQA/dLpzQWDR
jnAD3FXwGB/GlnsbKgZgj2Qtw5F4O3ZDuKu5EbkhOR3AO+hlZAL+7cctUwru6OlCdfZ3rk97XpPg
zkYC0VrLs6+Ul1pZCJl4cKL9vS6JCtQ0K3RXbkKBVFyibMJROyT0Ob9/ZUMOEYFbGrCzNPotfJrb
pzkQUllXuBxN2FDZ1IOuMz1PRjCjTk3YYX4Xn7345sXdNnFK9+84PdZ/BL8HES1YQ2am40TvsEfC
j5Rk0MV/iUnSxGT8MM9ywf5GPg0lbq3yFkW6FwYvdUlxwFjuaLvtv+i2+/O36GXPBqiAPXmtv6p0
NvEbc8CUyZsYdNkMowv9cG5GITf8gF/ajiHun0ThSHZYwp0mEur0/vMaUjXUFvnRCR02+vYCni18
DFr+3u+4sip9s56KNcXssPv+bsHpMVV2VoqdAZ55AZcHjhgX888V+0U9DDE+YbiF2QXkpPRof4zh
ZtX/RAxV4EnX8r5IrLZSSuwFbkLBYJGyOJ0Gi3RB+0JeCBCokQsHsbI5G8mvXgMZDUaUmgRzRm6+
m9iU9bLaeixG7UcuAYiZWBJpuN0B1K1CeNTQBzLjKuhkv5WUCa5srM7PHQCI7dZXfmho+0WtQtfk
CZxw3VOX2exv8R3c0n2am8yBCJfKbl/6htDp0hQMuOTxc0s9tKmKL5QNS2MKAPVGa23yhcJS9IBX
r7XQAh+I87/agMGqYMT7Wp2C7hTp/rPEC61I1/xnuuF/WDSptjPK/rJZWyQJTW4GmIk+YCMG3Zt3
Qm1jMcUdyQkjgugFZpWByXYOOjGoTaD2a9ZB1RhT9cot3lhpx2fvoc/Xnq68lqD2w1o6GWpmWNWw
en57XtL1vIwXKlNxUcqRXRku9IlxB90unKj7p4caciRD7gw8aIRXw98SCnLZR5skAHc15GeARV5s
k2W5rjXlVptawq90AY++iYeNvGGGxcfhTxayTL5BJM+hA4H8bEKCw2Qpjo1PMT1H9IJh6O8/yylV
CCTUpXOeRfvFsMHjt74tIDgm4Wodc2xqzHzDxwD516oZOpGgqQg1w/zSmblGWMXWrPcmUxMB/oAs
XxM60Yy1GWZ6G5/SiKftphUxjDb/raf+qfGxP86rqfGgVl6YSuU2Fta4RsCwEXAa1MK1TU+HIibI
3nt+9KKUO2bitebO6z59AO6mY3ACqv+HJOmdc7ih6dncSLkOySYrZcWbR5+fRXk2VpuwptqXykib
1l4wfAqM1l47F9SsBj97VZPJEBsaUyYxK3Rt5hAqVhb5c66Nu8pf8pS04qRVVFjgY0QETDFPNs59
+biOJ0au0cyK5+bpesvi00zJG8QpmpRPli7RPOVn9F+I/EZ2fHRYdoWmZevsvKwIfhb2sYB6iuha
2P4yeC/Y5gHfljj8qjtS5zy8ZEw+wPcWOxs7jLKzh7GZEYIEJXzDLSpoilblVGenMlCJ3ciX79QH
/hq2R1ZQ6nR2Ftav+jWPVn11S8rMoUbhrouH7puk2Sf1My9sZ4aDsMyxsPlx/etIcBb5hLs2TDzH
pLo29vWSdYj31O0d+BKugLoHg+Bo2+fG0Lco0IeaxeUYHhAettPGF0KN8eEnmWw+OrNQG94EVA8w
NKQkI0KwQlJMAUEM0Fdt6+dKrfIZgGsGMUaumXIoHAYJCde1kD6PYX4OQEq0ox28U/sX5sKY2hoj
gSufQjk/ec1/SWtM1FFNFY+dcMfgQ/9J5bJ1P3IZoajwTpKkiIlKEsxWUyE2kN57eEl7OPY1p48f
UDo9M7A5EjBqW3t7g5unijqh8dLc/0wr1LtbWl1BDD2dIJhwwnWguus2ByBlDDJodgUAtesEx7Pp
wbEeTzShVwmsgdXFu9lDVtD68N6umA2XMFpF16mtj19FDEr50FuPG5Ck5YpQewcdXcLi8xJTI/4f
Iv5PUTryVx5gIBzxVivyB86J0KEkO2GPC9SBTOAb/77YNlAtl0vWxCgwje3ZbM7I2AB1tFz0Zqmg
fIAOh5OaxETqhOwTRJKwZY+zwAa4JRepzWbPjCEcXM3BKaE7xeID+RPJWO+yTNxJjfCYgXiZIK4n
6lMP11NzlFGbCOlN09GrnYfLCv4pjU8SyGKJedpy5qNoMXGT4XGnRKzecGeMIFhHrlJkWbBm8QZN
w4q8AGr+RL26zVlgXtG6wtScSc/tU/PCkSu94PmHWJIzkndsZqHcKv2n1y3xXsy4hf1lEOL2ezNQ
5GqYb6phNb5qzCZJURg/M35Mv5TiPBOCSmqc7O1PqFVwxrNxhu1Ii81U2Zz9lyowZv+u5r6W09sJ
J1WKDLd0NrpAbmB62jU+beD3M/QaWD+Km4ir9Z9AGdPYf5PRV+MSW+uZxoFIVowevYqnDOHcWxmV
VO4f7J96k1T0GVM4TK4hkGEStIvUaI7mHoTxLjUIvYWdxlujBYPOGAJG49P5idHahdKKplLFz4ui
ESFwTNEwMLSjQyxMcK4nu63h5hxCPBkUcwISf2pQ2BweB1FUHghMlcq+cFdU3wl9AX0ZU3gT6fjJ
xo73rSIe0/8YnPNmdzp0dUuJUtAw5lX3ScvrwcaAqtivQoNv++cMCtyWKa1qbi640VLKRM0koU9C
kIYBLaILUCFevjMXsvqg9ZvizBLGoovoC/wRigbhPGsrC+OpSEZFIp/eXeGpTk1kaiiZZkna2MBn
Yhnw8Avvz6E+X7fu6nMTOq4ZaEjlthg+Rp7LfKSWi4T1ZBtPahCcAPV564x4siwnRiNhK5LB/hO+
0YS17gEG917T2VSvqxXZEuti49r57Sy+x3ZARQmECIn15Vhb/WgHiwej/vQUh3nODAZE0AnAHPLJ
9h2uCSXTpXss8+l+IqqMC5LOcWFecSF6S2c9Kg8Bj5/K1F4C1o+y0e3veWflw6R9zPrbyJGou3L3
HhS6IB5upD+C2J0Ph2YmJziUX+gP4bzbH+to3hZlBvDPN4l65JWscAb5PIDNaaPs4UaF/e6yrm1B
lFaiyB0W76BnRm1CSZuXaW139tcVzrsZ7pJK0rfuI310kw1o+lEMSRS+m32ggpTvU4NAKZVE5D+m
cf9md8gogCsJY+23Qxgz9J4RjutJ8U6VRviFYPQ0u+g21chBHUWrXp5+QTnbzJst/kOpDY5lXfZ3
kEqNifsrt/vW2bYmIwWKl6+sz6rYLk80JWSzIbE3VNSwDQokejWDLbYhlnxMJi6Q9RcWeByjEn4a
vrhulCv+UqVxfYa402lVr6bIxrYe3gABFn9S1I+KVhtdXSTCVBVrWhT+P0OrZniO7W/hqHc0+8nk
7vznJF8wzq3vQDekyxyeuNL82hbeM8Ah84NTWhy91AUtahuYAJO72lTVuqY+SWBjmUe4vL8zj89c
epDoRMa1XelJ8xbWrqcKfFLMA7roDrWYfI9abZNDcqZCDOPdiDJwIQcS3Y1dcb7vb6qwS7qLgW4E
db5oMoEKIjG7aAuvVXCIx53OF+DBQwws4cLWeUueidH+6RqTuw8iqorGnpc1tooFaD24cVM6fL5M
5BvUnkEGdv9GlCkguLbgtSXzHeKpuWtsCUOwnuo5ARW+NicYDsmgC+v99e1HwPcnfaDDT0i0KM5a
TxuR47hc3Eh6C24Kpk23sCfZZCOquaCuERI2Ot0BR8nZoUplIllLdPl7yPqziKo6F36l8oqas01j
A8RP7N5rh6Y+FB+zGmQFIJmJ9US82CizbQygd4fLi7h9Uue9Op2Z+2pcwkvOPxs4WMT6OuDcgClA
ogfgMGDTYu4f0f0NU1fFYyacz4k4Lgrxo0dIINW9rXcS4n1u6GRhouN/T5ubYR/Cj8olOA3WBLDr
XyKgqqiNYNZMKP6ng5Bc8TeCCyz4S54NCebSuaouAW6+YTd0lxmrVtNafhi+bcOzuzSvFzSrV2+o
6MsoIsj7eC7FFdNu9emiFQ1W6XpeRCtDvpWcKATQEGJ0VfjZ7QJTQRaPtyWjj+IGYjzPJId4cIpc
OHpD15OiyXWwPCpuud8TGc2M5vxk7+sfi8SNgXxe9saHu/hC9/jIM8Q/Tspvw3trsJbv1fEvypi3
+lhdVNkRv/TPXmKCeYCkjpXcRXClc4wEqGPf+MPBPgIvfqXDqMv1pJhh7vytP7h5RZFngSLsAc6Z
lJPHgGSbiWERuG1U+Co4sJwk9x4tc39RjMHiilNnngORff2RGgmrtecNpUrO+I3CCi75F9jEZ5K1
OfzAH3zYlyjhflfkrbIso5Hyt+KmUAv8kTQXf8w+J8yP+8cEuItu8Ap+YI6wlkR1uiPb4NSA/C4D
HYdm+lcWD+OP7n7tB1Qp7XZ17qt5L5UnEygCfXMfkN2Y9mi6l1zovuL5NLCXRdrprnPx3FIJoT8o
NSLfhXW+wxnZyjcrCKysj5uSBvb9I1h95ME7e2At4n/kUsCD0wp+jZFFEobERsfD/XcHLFpLylsn
5FeqT9SdkXYZxTsM4jK0WRoAifjS6AkQR0RiVEiEdNSK+TsDMMYo92Jd6bI0eyp6umVkZmhQk67b
Zc8e8Ly5xzc4kKsStSozo5zMzitOPiCLBvxhzwvhpoAP3qXbThHAx76izenC1xeFORcrxLAQfRIr
vg22/SOeFYuvTXKSI1bfiyIQymGj3biQVZvmDI3DvLZzKocbB9ouZ77OXd7Hekn91/4VfY6Vjbj7
7guhCNWOMp9ENqSDb0W8aG+DGylXt9C9ZIAxlG16RhbImoFJ9VEJe1lbV4YGKKJiDo3DcJ5XKqjq
XHyWbcU1meVctSktjRmyAdUBASnsXO4EKlNRKgTflplZ9AA+5S5QsKzDZYFWHe3sC/im27mnQTHl
ZIp1NmK+LkqKOoPCv1v5HjmlrJt79EeL2idrB8vhtEyx/rqq2qQn5Fn6Arr5ozUKZo/DDpkItlvx
nO2mXlhrO/x0YxvOLK3pVtfM3S/HKUAmtdaZfDiBVkrfSK45mY5mONDgYFSpgCCVChSZj/mcu9xR
W+yOW13wrLwnsj7Pf8K3ICVl5PlfpABywXIcXVpk/hGwjO7zuAkzGNCaFZlKUVMn54+QjWSRx4mc
10pgouwybNM/lHsTBrWvZ5EZ4fwC1mtPAvjGJqkxnzE2MI8XL76ULQnDfn1kj12PHnLvOObzwTQd
bm8X1IOf8LzSDp+3Au5wzXrwo1n+XSKD7+quEDKLk1pqp0xtzBKCrs2tFTME7VgTwQtNMjfuDZZT
FzijtQa4Qt67wtO5X/x5m3AqciDQNdcKY6mp9dwfL1oSoXVW+Fy2Y46cKcrKNANZEHfmxjdwO/y8
0zJz0kRZHJ3CEft3KkmFJJZRjh7tKwoIFHXpyKfVCdXWshxYWky2zetxs0s7HM4tNZfDU+SyusaI
+G/NmXC4MFk5LmWwuW1eSAftbwX74UbAdHqBcPYRq0bOu08ac8/hlKd+g0i6OkhmcgLkrLwDI6E6
ZOOhoe/VCvM4dcsJs5ZUMiZe6QydSywKwGPvUjDEAu9YUOmucO0/5mm/Fsa3y/ld1ocszY3OeTzq
wT/MbtWjmZp/QjHYrLaC9GoU/BdXvfIXv3Q8pC6YKMum9Dlq0n4I5Lhg/yWsgZtpMBHnwulaynyx
K/zSqkD/YCFh1iEdFvAyIpyHXX6swMN/GtY0hx2beM2nY81RDa3BaRJAs5pqPA/PT6Wx3DngvtMH
/ETGBAn9zbI7mt5/FZGUE9vtqnB50G2jv0MNuas1taZ8w4RPWqNrGcECzYun6XdHZrhxkvErGrRV
Hm/PuVpEZgyc6589b/kHveM0uTtjlAByIxQo2BV0fwCSp23gvb4v+0WC3cx6iWhvbc/EJxM9cPnG
D6v1tp8Kr85kZgUugcz+xhss4nAM4qmpyOzEF/HOx8JmW0uCCknnbqKHnto7762l7hiUN/5JFpck
d+EBbdlsAgO577nPmDvE6qTdqq7R1rZMp5eaLs4jm2lQB8Hwok2JrlxMIB2wcl0rJGpvoHHZgMBz
ics0hw+EgMzRZ0uJFrLzULCYcmNo628S7URb5TsIxfYfxaEjsA8laS2zeYx5ncEN3f/zvkB6+L4Q
t1Mm+0oZAzTvQvKW8tvMwCAvBH8rfiBf1+w2t/+2l5qYIqWmUx/VilRUKQUUY9Uwp/GEQ1FP7ZPl
4XOhhl56CUT25bnAyXPZHM7oEwI3Yd1EqRZWGCX2cNOrGjzvtwhsvMmPjJUcwY9tGOHyptq5bs+G
lTLbsVzTX/l09liat83Yt/t26YzMblLZjTlDEmoxcigbbRCWG8YFgZj66J4WAjoxiBqou4h1XK9u
4x5pnHji2vDKVsQ7kxKCmaF9LtIrHLD8r7d8L5Ju3uVTx3NSCD5BCE7j4C6yaNa3ziAZnTvkfKnR
jfKEYjXnBAt7p7MGKFfcTsZeKtSLx+Gx+XnT3oz+N7SmSWY9hDoc133GwtdPRE2FCn12DRJc+Tpq
ipzVgi1zIxqTB5x7yW+Pu+xj5vlSbGj86fHfnFyLStEzaPphB95P/4bdR+d9EhhfCZ3XOpKzkZgj
wLW3AvG5bPN6t46gJL0foSkqQB5ulqNmW0XDAO532RwL1vaVdZPPVm2s6HLsIb6Eak5Ealr9KRcC
VP06GqqelINIt73pQGNN4bNtJdEX9YuDSyFxv/3xgFeVuP14GUfE7kpJtDpmG3sJT0EspltdfGwN
4lZ4Sb96Je7nX4AurqMVIO+/DVnQSdYL2PXaG+t1jNf15a0QixOyPuLIblLaZ2BPPspMHaF8mXZI
XR0Gz1j7UpX4nwbOUbK4qMuj+EqVDqBI6KlZBVE3upUduhqwuUy/WgYoi5txwMtrHKYqyQc0+CY3
ybG8cG2/rZP2yrCYnKZ0ru8d/vG2KIHyHANXA5GNOywYiWm8Y5/1gDaWJIMnIEIIcp+HACfdnXvG
evY7jns95gbgVgfHoNlTBlgHI4OQdR83pmOZWBiYKAAzL/vMNjtcn+cbI8FOmEuPuD0zsQaBhhQ6
5x73Yaq6D6jsaxOeG9lzDrN8RCrWN3N3lOhQKZdvZN+dvCWb+5sRz+hqMKzA0r598I43WqPS6xg8
uk8yJ+T2t8ViXa3ltUOH8M2TSJ7n9IkG4f2lLsTbIUtn+mJ+tbmVpz/4YGAq5MzM6XE+exauiPnG
ImMr5kmt0FPM+dXJ42l9m2AcUhsaRlQdzKBtBv2zv9UAZsVVP1vKV8c/83CZ2Z//SVR10mYbgB2l
7owPEugRU+ghVogM7U1XcUn0cJscdLZ5OSV3cxzAe280F7PVNL90HRat1JaWqFxcTHTGeA6t+dvP
CrnaudADO5GV0orbbV1f5gzUBLxJfFvumoR2muR5i78VqAvWOerde4TSydJYRaYFS+T/hzqOka/9
t17IWzjFAu1AsJItKDuKZQA5evVj80StUyAYQP9XmUwJkCY6eFahmB6mmbdmwSkTBMuICOQxSoov
Arb89SvC/wOkpPBUDVH5tLShCnXnrJDf5UR0jgYVbzUKK+aH5lxKr5z1ZP5mc/GGmwKZbrntUOhd
NDMovz9jDMhQ13mYToEnt8Jh5fXId6EN7gFGWPvwjDuGwTtZhDFmziuv8rQnbTNy8Kx8n1JR/vLr
UNioSFefsjmNQloChTGSHVW26A+JoE4d2DWl/lL6oDCTBUaMc6fK0sGDKsjzhb/1H25991NsN1Rh
L+2qwOBcKDeMmchca9YvsNMbpprJU6iXydh3q+n4/jQKP0ubaPwejo7OH0BwlujEQfJlWS0TIrDu
Vb5wRtyDpOSUMA3HTOQTf7QiRozvylLXFYvJjYYlglINvSSgWFkJd48pU0QEDjJP8xGykaDV8Yvs
XEgWSEHWVFNZNAoXATZpC+gmkFGmrWzVGADSjdrv4RuoPZuHo+uORkMbo3hfmKZ89z16k8jqgrLo
XG+t82AKrl+OppJUCljBI7dPvH160HGgKsbPdAT3RVtAkmzeGxnCsyoICrUCBXaC+dqiSJCQu/2P
7bCpIyYNVJd8EW4TGBOh7KgZ+FtUXUpbVkgb4EH5iO4LOj0C/pQt6dSwLOXoVaXAe4KVwegGIqa+
DTBKRfXw8yTUOelkl6lz/O0kr3jQHuFZmgBGfhf/duFWSfxstLRxw4/g8wIh6Ie2zkDvFyjFYGGR
n4M+mNWtmBEJqvDhnw0f7vvYG0fpvMbDT0On9VsQNnvt9+GYSkZxlOv92Par5yEbQ113MogWsn/D
j2JPMfMB/IrxBLhGCbkMkgAxkngJCekqM17KWTndTwD2iro1R/mqlJvWHGG9PWL7wxasdVgDEVGA
egb2x+fQChv9ETC/beufwWU5pCP2iInkPwuVS4G6rBhiXbZR30qhPei6U9587lTwC3QVsN4vr/bF
xbYEsNF+xlaQtkSPpGJblgXr5fS7QSOefWUOu/ZoK/D+rpzyRD04BuQfKHjRms0s9H++XbHOfyX9
aKHU5z8nBotlw69Ol3ya7f+aUtMO2rSHlEeuyKvsjxSZQAZ1x6FPoXYj0RSZBUvRj2n2guiIremm
mkQGaqOSMZQAXWAbctt9DZmzb9q9iRpcuc3yO2Bg7R4VUf1hXD2/Xk5ykRb8XPoRKQFP0uSs6GIr
CMjgnt/n/7K28vzKWgYyCdbfnMaSL5Sm3vE2VyoPQKMebkVdv3r6l3/7CymVp22G35f3Ph+O/rA2
rlyB/onwvZDc3g3O2Sv0EEP3Xm9i6gyc2NeqcTT4xL2FhYfxFUd4Dwu4L5o1UCNnXSZNe/NgAA0w
Uu3QlGZvc3fty/vAPf8dJ9O/sQAGW8acl9a65YYVYDS5c3EQdUm1I+1lGrVYlh7y/+y6OXHk9mSk
znYkDV0pj829/DCcNVBwvIktsfJYlnwaYghTydc/8un0dH8Zy/i5tqFbiLFr5zebmcgqQdy/gYtm
RhEWg/ZJ8nXkT3cdNBs+p1J5i/2MQd7/kQ6VAcIs7FuR+ligz3bWIQ56/u69arir4kcqWux9hxdz
PqfK2xkI/74DAgyYqu0XRE89a4UNDzmvBl3EOxydtYzjyY/RD1ZVka9aaWZbE17sLKZeyzVoILQP
o5V+svsuJzBt2JcezXRcTovM5L6JESaWObVdjVnAidL1gmVtokhyxM/TvwMRQIL97MMgsA9m/+wL
P4VPJW2De10rLsGpvSBpaUcG+tVwT1u1659O1ZHsyJXXtsKWa+L4BxRSUIdwRU/Vk8Ri5ynxvXz6
zap6kLUZpzNV5MwTrkyW2kFqNEFKyHjsbSQi8nTDhpchJ0nbV1YVVmz3fuhNLAWujqLirwd6lbr9
JA6KqqF5byekCcOwtOb0c5pgGbVB+4Ee/xVlwMLA9rXet6Q3TutEmkzK4unASgxm0TXeD7ZcOAqy
PPIHs/nrLpDLjQT5fnrkzD5FkZoMvepK9GNH+zIOYWhabfmpMcFuNYuiTIm3VmoOnM71IDO1IcEm
8dIT5Zsf9tdTbs/jMcKKyIg6cpPF5qfOHePcFruyG0TtxJeka3VUiI4CMVMP1r3BpP2aRfyJBp7P
v5AqWX7wHOfKtZk/2NfNpgNoC7zoo+SLfoOEdr2lpUjcn90m83tLG4B4fFfCL9Uxfrn3WAS10EnK
yA+lwj6DB40+7XXwoaigbHbXu321RDyKLGp7udWYdhoZmwvYg7avOBHdt6zKDaLeQXVluZ6tB3Cn
L3YWhm4GvQciHGHSX4a6+Xj96q/4wR7Grau8GMK10XrkuQr6N6VzP3AkrIbG5Ia+mFUZFC0tTXw8
1gXqUOuNxgbnP/LnU77b80wOdJCQbKtAc87tanPJFkauMXFbF2PwVeOC2NBJkaqTtS4AJXuluAMs
0e72TTwiIoiBqgsXOLpyB9541/NHmLkcuUhMdLRAFyR3GpbgVPkZhrYFcHVfMj1vnQNyweZ6itSr
gKdb4pzSuMIprn22UXKk015oBKfz1WH8/0wkdFKaD3/DPLFBbbD9O0grpk5G0TfGd8sj+1SMa4+z
3YMMbuct29oZp+OgrcY6h0WtwdTrtViUxFNrXsHWZFL63Kq3GTS0vfELSnLAlEEPSpKvMAKP3zyg
xGSwif+7kaTA44h6U6HYyxEWrEMl16vsMAYMthHQBWXGrvTQOqf7Pqm889pN6V/XpUo0ZBlndD7W
5vN3I5PWcZeAG4dh2Pi7aU4DjWTYDZvt3DJ3YMCOGEJ9erScML9GPbmq8AUFRjZTGAyZ/o6hkBWT
J8KIqTrU1llLc5hsCIi6XXqXQvCn7c4NTH7Lsup68aQnVnJjig8lqVsIKcxvWLztB4xMA3Eh1R1y
gGakqHMWiTzQTkayBX3F8SqcC3HFERL9kKbb4OsmtREibYao4V3Wc3+LYpbIwQVzEaae6nxx2D7G
T4teK94LpYWedPr+AVAnORQN8tmVBRn8fR0toRq62ac50X1IPvfUW+52uiCO1GfVLMugRHRPMuMh
Y13gBsuNUEmtzCUQm6jTWNFtKY8p16hr6n67GB1DItlxYFA6/qx5AsU1ydTbvmWgt789Hb4G7lfy
76QaRNYUbB4Jol/rUQ+jOpUdys+d/pBUCwbekWZU9QJvvj86hmuG2ao1UbMdJpsPwX05Pfavq8H+
dPmUuH4YbElpD9nbva95HWdvx1m3jk7/lkc6HtZeVHgCC/dDjufNsPB1lbG8UBHNKx2XA5ErX+Vh
Rvm7LKtLcqF+wMdt25tucq1YgfP/jUgVJ/GvB6Ewz/rPZXDkhACVhHHGHbxCwnvD93M6iJus8hpC
D2oX/7UZcCmLRbB3lqPgZeH2xXMl/++LPsURdO2XduTaU3FFR5AImF3fdXGnwGsY3cQi/5x5bLgR
k6oXSIn6kSqEltA2DDn1a4I7fmkukt9pi2pBcicrMeEuPXOcf+dhZg5xR4inKGHwmImRRYLDY6BA
Q5Dey40F99gxxBEUDQKckL+yoZ6+aejRyO+QZlSim9chWbf3m82OW42Y0KLxvBpC9Lg/Vcev3+JZ
oYqW56M9qKa3nhbEJwOHivgbZSdh0PosVW2bcANqnYEbTpO5B/pVWgHUGmPf40i/iUdolUU5JIio
QgUuxrkI5ZV2NSK9jS0Z0wkUQlIsRHi3X8U2NyJS28UVzvgNzYWfrKBnJfuBSJHLajx9q79WxTE9
VbPU/RWeQRejPG3XwVozWM+mxl8mbuu5AICyJJD8toAE8gW0BKX+vbkohUc8fG5ExFCmVVL8AOeR
H0fayUzADmrm4NUbIY3zx+6lEVVJE1aumSvvlwIPpV0RK/w9ZzaZDVeMrKUu4R8koLB8v8n4NVev
mprMrtK32Tr6EBMcsLDToINgDh/Yn8KV8lLcs0mAhLoQrZ4IHvRIPlHVhewhp43AjF+NhiLAhgKQ
5ZxoR3kxME5rbyA2AeVvM3KHhzdb2GMYPd6hQvepkgssACdNalDUXUNzduzUgxXA24IxhDXeyMH2
+rN0OiZF1R8k8Jkx4r7vkgVIUCfnj+PFZvT9V8GKHmFOuQIcKZpJhnn8nXWljy9w6iFBavUFyKVI
TkymsQsqXmcchMT0/ZoQYxlvn+QWyuWjeMe//5G7SJjZTXz7j2l+c2r6YoEY+K4C3I7uXmX3Pj4P
I5t820UzFRRToJHurc0Z4kIhocsXCpXUF21etRn+TkGbabDQZ6Hyr/sGgF00O8PQIsbzjMKxmSu9
LYU2y4XqYxrnlK8m3HlcJhylCY7qX2rVhUxkPj4MdHSRLKMPDLwSmzuL4ImdCr7K9CVBxCkQQxs2
Sf5h7Vx+GiMQ04f8ZjnDuvy690DtbI/HbDR2MsRuoRdruyzT5ga13ZQs8kITGwdaUA6t/2RRqfY5
4usm4sJ3PnY8wHbN444qdD7T/5EZkGtCWFSGaXlWRxctw3miH6ELJP3aP0fAIUYEcVuyVaxJbq8M
aw2xeMBNElI/KSm69+PtbBEgRWit8tgDtCsD/wmc1exZX3WWmsv+UfBs5putvb3cSz2q35etCHPq
xTl0hwn3m9BrOI2yVJfVEhtIZLKH7ri29Yoyv7OaqohOCInGOIeaY8TzRCm4m2Q4DtqQlKB24yd4
NEVv6NDhRvZoGfxNSN86hNtWnNsXn2/7rSGArTOJeqevq3O85E4kKazi17cRqAQYR5+g4j0P85Xc
6sPibsMGUPIBbtexDGPXz99b2V4ra4hPvU6ldPGW1G3uZy0swQxkHhG3P8rkgqVQCM694vNS9Ai7
TvP0KidU8k3JwI3Tr/C6zvJiwVTZYJ6szeGdpfC4dmxKN7I35iQgzp1ptmpobpQVXqMN7otieZmN
ps2Ujc1jsdxBQv3JQLo7v4bIiB5G7gk8i9V6C0qCkhg6rosiCa0OJeA4ejaTzC60VYeGcZreVKQd
h5vZBwkFqH3Q0z2aCQeAfC0U9JN4tK+hCoOB3Erqg2b5MvqyHBBOn/uTdd0Ewm8FBEdaRWOpY3UW
/leFD3HNszxPtU5/BgZ4XKX0JaQ99ZWksO6JCjxhksXlc2eHKH1krVhi3kXG1m3m/wE/dxC+qIuz
0hJgqrBuIwCh4Q19gEF0d8Zuh0zNB/WNOMCJqyA9XcEgawumG+AtfK5e/6q1GKY08+M5BlBIlY/x
Xo7jz01xlyA/hq2q/ZqHyl2EF62BB0UdQo5CDB3rN0sUmVbrARJEt9/k4aLgmzwX8PiUghyLpqql
ARtRDboRScIgIIx1wMIVzGPMLMzGrCABNehEHW7AilTYEAogDhtPYQlgfiCBt5usuoFIBPwwHVL3
cjtuKLhkjXB/4+c+GALPj1R8qjlkruskDVzGbOXDpcm096UsiM66UniPXrxGIqMTss6eE2PL/oRX
NEiUnM/jzyXk6TL9xZ9o272hhzXTWBIQsCBJD1wq+cyFcXj4qjbevKLM2efn1OJAOnClJBI/tlnG
/qhfOHbJF2QbeeqiGZX6qqvQ/xEqyOHEPg/SB7su1HrUtI2aAhFhWIqmfSnlc352P5VAJO5PrKGX
5GV8OPCaH6VCY9o5k4eyDBrBjQL1NkTUlruiehfldA6MtvnKepgLGQzlITaswtT9yN82CgCsDF7A
Dkg3zQM+Ql5PRCXz5b5Wbv9AAxwKk/n3CR3IZtspxwyGoA0WA9E596s03V2II2m0YQ3GRz2vNUD/
/ToBmvlxblCu/uQVJjTsYwDkAqrT0pi3WI5ULH8E7S2T24O/exKYOrn/Vkg3gRjowpjD1JnOVEID
XgpguwX1l/Hk0BUrvZRwGa6BMhc3cda0l2bOtzZ8832ZUSmcMXjKqaZCYa5mVZ1A5kupDV88rXTb
KHNSmQv93A1AEBNHGTFzJjE1Ge+VJyFZoKBRXi9wve22BXEQ7HS4N9x23m1GAXpZuP02hXg/p4KB
/AD8J4cVoHUd8NvSH38yemOCMCBVlzoxxn6tJG/mu56k0sWHMF7QsvGRRGNTiqIAshC/J9/aD3iB
bKQ3cRuCFlvxOI8q1bGWBETPmA5UejKmP6SYbYjE3I471boXIuFivPMTBKzoo++Hv0kHqTrZ8BUy
epXxdSQzMnqNJ05BjP3oXmct3cWScmvG3ujEX/bsZ5OXx+31QlAvQd4smunFcOct4ahTNOXSuDKE
k/ELPK61syidigl3H2LqT+BwGTG0a5OpqgfOWI3ww15BwFTwbWosvduNZhQEbgqZDfoDxyuL6a1m
hH9M6px9+hLlW7WvhGX4cxdIu2Iwdb9qxWZZ+YViyXUXAsuxa2p9ld9wIhtQp8bxjlU2KfFWU1dK
z808kQKNq/hKzdFSr+yjXRQfNiYd9KLGFM++rxk71e/r3zWmuIKyGPLmjGQmOuIZDSmcNLL9oNvA
sUm3HLpfgLUvHiox3FZhihZQgAuXgd42BxUJuc2CiESSlHK9zj4Z9CM2yu6PlZzaleQkmMudBsYA
FrR1w69hXOG7h1yV+hUCVBwbqPAjsCC4ZaG7334+QqlFnal3Pd4WCz2CThVtu3ZClNRVLeLygVHh
qgMFIcWjtNKooU/l7miaJeB6k2bsgMXhHLhyD00QHNbcF3bI/ffTFzFiXU/R2Kl2tbmECPtX5+3b
hysatB2GAGEToXh6789HusFy9+NCW1lhFz+dIquaalEmFihRaxVsTMXKLR+puw89pOdkff5IRkkU
nt+5hIuliUYu5NZL8jXqNErpWNaVjtDmhea1rnUKt1iAnnvZAJZL+BTb6jW0sw9fyg8BX5fbwHDa
q+gIPZlYjkcySVF4eSr2UhKyhVfNJ3UrbUdWqFcCL6hoRl6klLduremNeRiASZV8uChFTm52pmBh
id76CcVTJS1n9U/Pt3etm3fandUUy35D6UJQETmG/SRWkqLWAGWcQbkGr3HbQHtrAUj5Mv+n0+ep
DSUJ5oDhE1t2FJ8kdAyl96ZPTY6a/0HmIB1I6gZcLj+4Cnhn/oJcaiPQ7sGe0SF8b7rTDDTlno5W
64Pg6m1BHJGwid0i//+095qm0O2zZeZAONfq7Sa4Vn+0G251rIFyvOx/IuCdu9Br8a7ebRJrwZnR
i2XYYJ+vehz0EWBAmymOczmC62EIqLJ1Dc8Q0dhvinRVQ+3fWAiZqGD+u5m7mNuaiRWCEdm20Mb/
RlXfPW3hgbDGPvwbRaVPc7svYspTCzF7kFbB+zu3CjwEdZXPfCO19Hglh8J/ESITT4s3wHeJG3/m
SPlrjKnx8hLuP7WEUzwowI+oUSK7QHdiQ5/lZsupPqN4U8Wt4FqBt/o+vGzVStJGqas4qpf2VkU3
r5G0EcVhfrxMhH38oc18GPwIvovwyNFDhWpe8MLwEcuX3fO8bTVcIKXKscuAvKAV8Beu/27ZoTX+
HWRS/jVBew338v8FYDRy49YYC4xYJ/H0YLw8cKHXSZ+CkHQNnlrt3ES3GNB9GvVM6GKUZMBmense
oe2DFWw38AXLXhLjZYgthhPenWEPtlhPI/phdY1edxOHYizbzj0yYKDViXB/7ET8DrSunJegqnnp
ZgvU4/IDbINE1TkE1ihCNCIlkfq2BHuXjsUBbyq2RTGAjvb+hvWimjywV6ap1GMgRPuUS7wDlv6/
J+5K+3psn/XQe5jcGXWVQuHeMB9r6X1yBG+lU3J02Y5NHlXgEqNxVk2KP7LQg5aTMLal+RCI9YBZ
gNii8/cQpxClIs+eUpyiYe6JH8vS/ArTToB0Awsg+SUctKTMHGOirdJPQwwkNaVrrv+p8AZaLyWI
ItDSF0wFYDyoXrlf6J1FwfJ1f9pDyQNPgM+r2ZaHT3FsVrX+qAcMv+wyWmgntFlKQO0z3rpG48AF
wSgZOpDT6Xlk3SeBW+KifPjB3r5Ttx1BkInDpXPLCQBavpisNIErKkIT+D7XbdI8xor4nft4DrVW
xhcYpWnnX2wCWs12XpRq9v+fR0bePv4wiRzWHNF6wCVwOn1poGQhHwot95uM6ukWuRe1gnjt9EzS
r8zf1Lv03q9nJodmbmN0cX2cfQekFkg0Q5/j/XTGpTOIt/CBZTDeaMe8lVFgTRKTcC6O4/Uo5AiD
pP2Q9rkBAmOvRqCboag0Z5o8IVKCTyBWz6tNT2YsydZiquq0w+bC2K8DC4vWJYjzXZl21JND1Zfv
D01o3JjFoMFsDY/jk1R6XrSSRwj/lZic0Ql8qG9QGbGObVrBh4uWIvS1IWXz+/ZGxP8L4Z/v9nlX
BSH+ORB9jk9mBadyru1PeTZftdOFiGXXcwNglEbqH22a+2dQeqIUK56gsIPXgSLvBUsAU8aQfxeR
RaOBoSqbtQa5Sx+yx7s6tnuLG8lwzU2MVkkcOgH+lkEd41zVuy1/AcxtXNxSze0Y/FXNuTe5bp6E
KykQrvJAUFMJKYYrzighFDNRypkCdpvr8SvTe/8BDWpjWBhWVjXIOjiHaQyM4YAQe5UAcpj4QfRz
rNnSeN46dUxqyn6UGc3OWOHGwHnNZB7/hs/joxoY4pX8+wMueGaagdpIhJGPu+m+G0f47Tv6tZ0D
huUEjNiIKKWNZ3hIStpecaA/sOmwzeLrEb3qffUEXbdXSMvqdu6rXSxe1sg9O0x61s5O0s7+30fQ
suDzvsKlfLyyANUMStnWAXPzGPWKkKkAEIgy8pXLAT1+LmjmjIs9TFVGBJYretvuh/bGuuM5KOJl
x84eVK4kI8H7j3TTNFgSaRvbB6vwadtqf7tRQFQi06HRorjYBCCLLJCeL+A6MuYXArdhXDsJBkqn
TacWhY5CCilwE17Fxkd45WPo0cS5+vjCGMTqP1pfzAtATAiiGVQdTMbtFOBnFY1S9cw5n5H0VYSk
bKHZmCQkMpQLUFtNoeBFf8OYrbLIqwvRBgiFycjIlROU6dQep5A4GDIUcoxXJkQfL9f6G8URCJdK
5ZkQpSCWZdYA/fiie6A23nqDUXrH2wZlQqcHUWTEdtarDjxJ8P+zuM+BLLyPIEqzzBUtlC/AiKkt
SPk5br3Xau7RsXkRKg1L3WRuvU/NAiNid/Iongm4COGQRrQVIbo93qDgtP7pNPElMvS0//Bztntf
O034cK/TJHGqwS1UAa9THTj63MflZyCRQqEXNfdozEP5tyKWIOvjOGuqo93Vd7WaXol2t69vdtM6
gIh2JtFjUZd7erjJfcV7RNCa5jB+35Yc19vv3UPHMSMUSsN1ff2H7vtJeuSffn9frpl2s0Rq1S7e
wMb2Yt04e+8CICdEvJoZ03VBSjWu3dIbI+UAsta8KwgcRWlZMdAivvNdX1U0vTEW7SPliRF6W5bL
OO/LKA2Gs9xQMLFg+xUXx4Tycpw7iczZfWJtatxpvVqpkVWe0OfJuvUhGJ/O+4SJCOJlpotyhtXt
BO7qIyVn48CDA7JBX1X/hE2pjSKjV5Q8OgkuEAljNMtqWpjS6GLugYksnTMluPN1sH8eU/a/OoHJ
pE5jttnUr7V4bJ3i804mmHM7nzMOafT0/GtEO7T3vSS/TjZ/H9wyJi8Y2a1zJxpkF9XSktl8MHC7
LlVOHlS0MfxbNKPwaOkIS5ahNPiRbx4l3bIcCT0s8oo1gackeFdPq8LfhEAHQu8jo3WL2eVeFna5
tZ//ftKeRJjiMgy9hJ29TgbgJNsl7c62qN68m16NrLtsuB+bGiz/lyiwgwJ+HbjHdNz7ZjhdOaEj
opp1B0Jr0km9wlap05kP6I918Ge8QrdkOI05pyXFFPb3ZkFlmZSE1Z7j8GHh9KorkmeMnz9KqJKw
KGwAwzrVN0efDUGOqOMk+Kr+nORGGK8KingPTkj8DgjsWVD48vtpzc18wZsxqwgurcc/ccKmFFnu
nGUquz4BqbQIuXH3UUX/jJhks450aMgeC2A7F3/HZsh46Nk6mmW/apwO0wZojkz7wZ2BImjDW7hd
rkZW6+J92QM9fRYs1y8LB2/aSh33n5FfeMkn+phm81WqQexj+u/79Vo+uEt9ONIk29gwtUlGv+eU
HVJCGsoZdYup7zkEz7SKg2+2TZ8WNTq6kAXNG+BJRAtCH9Xa7jixAXCEu1rOyWp9VcERgBkYNeVg
u8lIzd2RbCa4ZlHbJTWFfFZ92tg7bjxZcepaUnxrgUElAqL37S1h5QM5Ush4hE9/p4q/7yaf7Ljo
Ctfvm5GPgOBSaN7JRfJIelS0XY7/zIM7jCNheUoYgfsMFDW46rReOVFw2t2dk+Y7r9ZLr2YxUHqU
b0CkUg1pKfflwLfb1y5uMUgn4hJ35xPsRC9KLEtmJ+XCG3GjXvollf59PYPHOMYTgbmAYRvbu1pv
+dDETvg9dwnPCmCgYKKp10Bkjl0ECDUkpSU7oCYHcm7fvcf4hAaBNbthMsrZcI76Kp9uabkhajjp
2BXudE6D5aUHivFSSoS8RhyQoqpcIKq+apTrg7tzpCPLXzwKZNLwiUgqMnN+XtXJi239C7q4HIZs
weqb2/qxysvtyK2VeCPh+9LXN0IjM4J4N7BfDYiVunu6xtO1VClfNwJYiX/O16m56p1Wm9PXT3wo
AlH96E8ERqdGF1sgVuVaO4KU0Km3iHxNg2LbEW3RNjZkjpg+VaNJVqdX5M7uUFEJDVlNocIZqdH4
L42PV53BgeYdTAV6Bd5MD8ZdiB9m27LQz6czTsm6TtDVLDd8VwwZou2JccPtaKfIXS4fZcR8cFNd
QLxiL2t/7O4EMfjUhW19Uhg7FlX6AMTrlrhzBDJPub/t6U/QMFOyhOEfLdgNsL969LE6TkQfb5qz
BkTjwl6LQoppC8Pbt+uE6v/6zMv9P3sxWvUe/94Z10cVtny1NF0CJeq7IzuCIj9x+JW9yeK1t/iD
6ZrJkeIJunbyNtp3xpwcf2jLDOefgmLzzvWlJOGKfjXwAU01pg3Y1oprfY+V31JsvQxNZHDyIhx3
MEJYPWtPcXtU9jpaMsLOb4WanFWHG0Zsg3al9j1l+WIm9qHPaM2gX0LPhFS1iP2Uaok8I5eKibPX
N2kWDGje23j33TDJ3bsXrSS3qOlIHAhU1/edZzMugDmRu2bN3fV0vygjR4ZGdeo6GzNO+Hm+rozM
3p2f7nVQJsf3wq554cXk/SKbIlmlCt9DDYbouWLct+k788AAS10AAAIgS3VWydYonwc0wtSk2RP0
eoyl8/cS+rADivRL9mjlLwzc6XEiFHtvUBqehxDA5Eexe3uLSXK2Kjs32IwMrjuZAPVeKY8V/Gas
KREp3KlHY8QkNcNGNKRmV/us1gygh+3OyzcnRB83C12tSrNZwQRyt66nNibQRXar89+82J1Uy5u2
Rh6Zd1g9xB16+E+GpfLok8U11otRrdcq4pVkCscYBPaQ3g2qVg0rywzJfdh7RfnDVv7qYJDCb62k
0KPMQj5QR3MItwkNqY7BDJwROKe6H8aMfrSuTbY8Rvl12Z8Z/FqQXC1SUN3VoNHNXci6i2FUDqcT
+/P+Jm8XFnE0JL8S98jPjAOS8mU1M+lQqIBWZ9Z49p7BGA1vdUGSnblA+0UglOe0GA8ZrAiTe0WL
1eSU9MT2WtxFZMRdm/XeCgfKseFUytbSj+VWwcyeEXGftpcArPkAknRHEBe2D3YQ+g17gwE5CKUS
6nn7pXZDHvT3ef+W4bmK64Jow/w4N/9iba6jADyGSKQ9lhqOlplw4zaoJjyL67AgoX2cJGuh+OC9
9pxUGtQbnhuUb0GjwwT7EJegdJBt1bbII8YzmyQUdZEsyNOdjc3wt6F+/oSQ+0ifx/u9RgY2FHvt
83rmmUlKicKS6+BbzLcC/fXxEW8b8r9Oj9e9WQyxBZzdpYH5hBAfjdYW4xno+PZKhtq0lvT2KSKN
hnwsjW4I34uV0HbiLePF65EPv4nf3wG1Xe8jJ6uDAhoP36f8ZWigMczLgYKIPE9jkP2/INTrq95u
IF9DgWGox5Dl2nCe/l1ALvPitY+wFw8Qtd+Ync93gp/xhr6vobAvrU8ozlIG8x77mWh2jzgdQ864
LyIzGD28Qe3xt7oIuu+DG101u1zlNxbOmlyrs/+nzVIqaZL13syB0oKOQspKhkQI0nPjD50XT8KA
j7lOdJ+RzGPr6bUG1k/7cqCyF5QDYTU+VhnsQWSt9+ay0eRClkFgPdR8wu58XXTBYrtymdKID1Kj
ChOZHZFPMi9v69n5tesoyWXS//1XHtL1PQJnl83OEGuRXdW92/LGNVwpilPVldb5kFLKfm6XV2AP
vZlDHcAcq/whQ4vMEuxk7kOioB02r4JTF08yqDg9pq0rAvVgOMuaWVXB8pQsDAW6qTIZtkh8NlRm
HT1VUQCEVtUIWobkKiH3AIcv8Guu+v8M4tOgw0oNtdzDH7WFCJUkUHPtU05Wm1QcoB7r7wo2/0DH
YZKSFw2KiCUJrh0jvBOHcwpKGI69uaz6Cc0MfLwYVLvIdbDniDyVDYdE72PTEBu4S2fAic/W1pdy
YfQVIkEHD5bsNePZjW8zSdzBv6vjf7Wef+fsm3XmjC1DM6FueQsVYAs93UhLGCLIfzJzLufKg53V
H9/qB29eefP1JZupxCgUFw5ZZnk22tGD1F9ls9bjUs8DSIiEkFZeUO1r681EDbH0F3xlJK89NEWc
k0AxqYnkMAD1R0EKSL9dX+udpdenDIxWqpjCN5HwZaDHNhJc+N4eIrDOL8Efq9rgk8HlZjW1ReY9
8/VKxwegTIxrgGfEq/ZPA39hZ/pl+HhE6oxXGShUyn7o5eZpoDOeYFq8jV3ksa2ec/bh+25/RG0j
FRpDrlPWw+YTUUErLnQxTrfWG17gehmUwJv+j8rcy10vIG/21M5LVmeE/4usxRco3TgC+VQsuS61
/TRzuH6xauEGKsh9zrajOKauCYKxikrGF/7GNXM7ATqrOnEJPqxDxEEpm1sTStGFk4BfVXtVV2V4
tYY5Dn8GSIB5XJLzXvfikWAQDRdU4DyVFV+zvLe6SUZNYq0jE2p8LwwPFxtysgfmtRQnJZY2f+Dc
dfTTTCbuTBW3KxdQNKAiswIRiX1G6lTzAhGgzefZEG4ZxD85pIz0/YKzxKTA1l69ycg5KHG5gH3q
dHzdm3rq/inG7yHSMokZNk8MhApqUAtEHd9moghoVGQz9dHSovBMKJLlH9PxYFcJvDkeH8gVgQQi
ezMhackqIvxMKJI1lRwGwhDcAJYLnZ63scgAwJPY1k4c+NOq74OcdKHOfSR4A8U4s7VIO7LrocZH
VhzHkRVZTNcYj6Wyd/GDitFkwjTIGgssC7YZ+OsH22ps00NbC/xk6gsXbOjPApD7N4nMQ9u09NA2
Crkz8v8xeoKPCSGGO0HnYHSTSP1wTSvW3vZJDxyVRP/TeDGliD88ampXgzYK5R7TumCie1tc+9G3
DmUi2RorS81BvS0MwqiIkhLHckprOQO+rUnuATVYH8dwT3h4mqNl3WirakToBg4KZUzCdU9LFLdN
n2altZEJ5BxjTVtkg9tSfvoKyjM3hN6v/Z9awitQZCg8I6CSkqaTfaKJyijQuUZIiFeM6229qchH
jZQoiEDw8bZ1L6nqO4QvB3PAidH8yzRJHxYkggTEEJ8DJzpJbvtVgH2xCjBHtVzlwR2lUmsmsQFM
GrTt+9E3++ynzxOILylW7JRfpLNhts5tFer3rPm4vkyDE4DbA6MS6RbigbZEzkAJS1V8dOf1T9RD
4QqH8JUwB0LQgQkF3Gnidir3fcdmq5hFAdfdyecYs6qSuywM3viz68LRxLhx3yXU8fok24eQE7s1
4GUexIw+W/EOnrW9BKQ/BjDWTAG00lDbgGyjMu731V8ItdSsK1vdoAYxw6RNd4Hzdt5iY6ktzGDE
tw4CBWcHTtfgBieV5FRhOdYNAi/YrWp67PN3Tg6SX/ix0STKa793lW3zChqWNqzV8OLg7RSBMOJm
8ar4b2j3Nw+pepSZlljDKuI3n0mYYLvpnbVXy7MTqyhl+xUAmum//+bu4YRQ5IjBdq6m5JSJCkfc
UIdOB98I7tp6aLHAwxJCHUQw91n7sv3K2KwG5JgsozdEd3fNLCVrTi9HKa29wsyjJ6cJVDF3Hcy9
HHME97htIrvGNZzMak1bon0z7/zUGIFSkk4GdT7jMmOLGVuNXrAW5D/HProBFuyVYQdy2ciW4fdn
hrKqZ87G7nE+27fxnbQMV65g568Q+Blw1oO6mTVPPUgHHhC5pOKQDQDC3/ggmRHKBpZnilrYCqG+
fp7GTVj0Hw6sGQnu5wkamJOBkdcN1m2YhVyfmmg2Vae7uSD7CG6NrDyW3qSxgXxPtlXUoNTOfouk
Z3CleJfyWQ+AFCdBxRTj01TvSI2wpQJD/Y3ECKqsvi9wI4AGgejTsn/PpX17JK4Sbn1w5Lq1352J
egICBLbviN0biHHL9h+w2UqOMC490LlK6vnZah/a2onzPYjIkAvgcBOWyET6c0O+bmKN14A2/i7e
bdA9Alg8dT3bDKYDfZ0tBdWOLQZlZMo3HKOBV3uCBJjba/AJro/g71kkUQ1byWThet9gChWsO+53
hUY3yaOn/4fUL62XpdroentEh+W16bLbflTtxUrWXXLHZEcbUhv7kv20sZkPhjxovY2CqMbez7G9
/Wy7JaIlGEmzYPD0dHuDXSdL6q4bezU+m8VyxRzQPWSY9CfCdZQxDhRj0iB8rrU0odjLkORMzUA/
eIcF7Xll0sfcpIcKvQhJmxU4ara85E3spwh3kcnYAa8loxUIAtY1G4DezpAj20uSjSot07aqlSPG
kk7A3v3oRvps9pZDjSRBIbdX0xqcvt1si7w00fMCkvA73ihq8PTDDoPxLcRk5udRuyRScIMR7/x0
R2BXGRqIy/pLuWIY6gW7xsRsW8Bc7a+GkTpYPNkEb33sK0W0KYPind1lNzucLPQU8gWks+dtF0Vt
jn6lSdYm9E4n/+kj0yt04oE22yrnV1GIj9cV1XqLzhJEhSW3NB8e4aTAEx68yI8RA2FgJEJ4CzFb
rcIhY6kvHDTFi+dnIFt6TvNX3JplJw0oX3rd5sAN6XtgcDw6+Hldrul/F6fmbAe+S55AUa97XpTj
UnlwF0cnN8Zb/1KNBX/fou2Z2Dv3kR7cs0yCYu1hlw/clU/QsG5VewNTXPAeb63Qqmqo0+0bopqU
d0n0DVvaW0QvwokqpENT0Om4pEdIHadfqtvwFctemTx6ygGgjhFZwryTyAJU86cG+YmXNahc0ae7
7O2zAoK/3719TTbDwz30SgCtmujxPWBUdYxgzMj+tcll/4SND9aPie/VhCNiXZfPXADkX5y33n0S
17oShPKheJyT+yfEzcCywaAkfWIBXr77ULQDIJLjACOHVkCtEFRUAz6KQPXabdpwKQZzUKhv0XYi
AiVTVjXnTbQ00asNMztdnO+nAIPSztgk1VfiHpmQGFPauZwytoHy0wJRp0uYU5y7kkcTnf3S48PQ
Qo+8tFG6Qg0+5worvxWFVf8xNPCAjEIRx5QR7yd9tzY5FKEHirwrBWi/b5gj7cS+MVjAI12sDQnU
hUpDEfGZMLZtla+9ojPR9dkj4kyTe4XYjxyQQdx3zzZPun/rmKJierFtu7Q4MJTQYCwXYZ3fGrMH
P7xvxUO5boxZMrxyWMzg0sEQI5eeNWf8o6e7J9u3WLvkx5+cbD/eRTHaWcUkRizZhZpWVSOwW8ns
YvbUtSOCnwvhlCxK/DkZrDSg5eeAFePrTzMmMDQbb5gg8mqSzFR0IiIldvjz31PMWbnKVweobs3x
0kI6IaqfC7HOEox4FTaaFwy78B6aJNH7IRPEhMPtFkwEl6wCz2jjgJFbCxEmoXbF2KwLzlmGDJy6
ZkxhF4skpo0q+FphoFE9KPntKZysJkjuXfrmfo8442MxJSGie1yuocDlLGM3nHHfGCxQ/iHEE1xC
QU/CffHfF+peR8YDJ3GbQW5Q25M5j4pKZgot/meDXV+haNqITCpGGUtCVbdU4mLuUBhyrB8EybO7
XlARrjnTVsYeaw8RWHqrP43CQpTxlQiuWKx/XgShjIUafvikKmU8u03Fo+ZRWUjj7eBy37rvRTko
6f4UrwO2HsLA1Xxt0bWKn+WNRRIgpC74clYF1veUVEhtbWpVprZXKahI6g+wrgWFIhI6fn5e4jgV
bV9gao8iFVFav+1lzF62rMXud2W6WwHBAfaBoODOvm+0tq49JsCbvINmO280fMtv4vOxHCYswmhA
lyo9pFBEV8DizE65LswkUu6ut5rfT+6fw7O1MmakTtM+cV2jnek1Qm585r9ePL09sNo/3UUWI1vC
jQOiiSslwvieX/9Bk/W40U3W/XZXH2D1/R1/GyT2sJhDeGvpCO5Z87+ZibH8eCPTID8GuJdjnIUm
JYBFQZesPJEgCIG7ibSJkllzp6AsfGrWatjxNpt1pAgbNKCmCvq0XCkXHzkHUlGujGFiX1pNpVN3
dnIOhiR72cc1X0cDXPdvJ6l+Ctpw44mgY0uoCf5FdHEqExO2KEoYv5j59CxujrT4gcpHX7HW/t7V
YcERRZQFWP+ch1SevlJyP1PqBQpK6URsCipQ+WIncHI8lU+SFEdF/b27xVTqYTc7WxYIO6LDFxer
TA7k9+k3Mv5SxSXrE4USBWfb0Nx/ko2EgS2cPNrR+8IR5Oqt3YL80+LQ3tjYjTIbc7nBwO73aw6V
hSk8ELudW6x2clzN7SAyXBvFj2hqrdzaf5mpjuQku7jeMIK6vN9e620dt2nSlxQimchK01gqpR8r
NHAu8BnSNJjNK82tymSPMIjEsmKgEV0pj//voOy4r8zYV7jyLAa26blV/BgmiGP/5mOrOuAxJTnD
SgR/vczjj7vJg2Qj+ODz/ss3V6gFiruR5OZCiDp9259bPFHrj7I+OKt2PsBYXQQtXlhUzB3M+K7X
4YkU4801fhZ8jIFyZOyGSgHsuo/ptnMfoKkx4jxCDtmg7XGavKjtYyIIKa5BwpWxTh70v79A2WVC
9aKvxd6f2cp8TQxQRI8KVhdWj93eVyj+5SourGQFpCOp+RUhxoXvqxeAl5EAo3alamw8ygA6Y35D
i6TjjgzCdsUi8iTDM3uHB1iEyll/nkc9BrKJnc+pkPepzbGwBw09fJmpkPM65TRPgpKmt7C7gxnL
CytBHEmzhqUqq0KxaIOw85oEbX9DdR9hCd837q5VE5/agcdfOc7KFNdhUal5fp9Rvzen/QKdKW+F
lRZfw2BtUW1VeAjepYr1ledf3OGcz55N1lR2NLsVAnP9yd7tFyjG3oZ1othvGQcCZAJ7JqyYxROu
IScbhqzkhvcSRjbJBGcAGSDuQwHCgrfduvrrBj8lzr6ju7W8E4D2KbJPJLm6s9UxCHSrwQ70+SE5
cTdBhVpnj5+XHbS5e+YCx045L9OtlAeToFshzP20acrhyaC1ZEAid7u9MgZcnBFzlQbKVBbMXwop
VRYrd9WC80lJBbUn3AOEpuB2dI9vXLDSyvVbdajZZnI+vyzdtCGwEP7EqdY4PMZuziOmTee/AmYl
osw4z53dXBvuhQAfPDS5DUHewFH5hzhXtL+nCAAdRnobSp3Rulknlse49Nf1ZCsUZNSrKKoAqnPL
b+FvlAgmW9++FgZZ8TvBhAHUrboK0e7U/htniWvS54VHWHN6CxJcWKeJxMvlGYO5xy691YVey5Zi
gxPpko4oqdPrTjJW3gZSeLek/3ytZgo/cBrQtr6+gP7ugAasCuecWd0MUcGGOwCWrAt8lHFNvuPX
zzfIWucJsNK5IFqC9kIBUwYl285GoEC4wux8NDP15JRF06PJX4ziZyiEXTpX9ggYL1H0Hw2ruHoj
LEriE6ddS1XVOPG2wE8PsUK059ZqsIiRmoWmk5xwEFvlte7S0T+Fg7QC2aPrOwHgrhSDtpZkch9E
NbqcD1joa02+dMJjjKfQI+HCsHGqRCvQ2VfIQNix4dXuPCdzkuUTB4Lf/Os2I0zGZoPTotnV2K4j
B7Y0z/0sH4gcKFLLiZSSTTRQjmuJGF9vuK27j+o9VqETKx95lcz0BpvC7uKIzMjZrTUy0WrJnfLH
qjiEDi8OH7ol8f8+3xjDS+QZ95eOdx/kRBdAZOnEUJucv5LDUJyoC0Tz7/5PywU6q2EuO77bjV/a
5gyOKHiYwifTtsZvYQm08nBA/5rBxsSGRHPCjCnU75WLPrOFAg33met+Vvy/ZuxfBs8q8cvTaDzZ
spKTxCVIbbV9wuH1HGXnEHpMP7UTNvbZS2C+mEQ6NvcO2uiy+jFNJeXVEwdOnw/xnwaNovWIP7Cb
TVro2iuYjvBXbGhBAfAODPHtAKowna+fM7gQfB4Nnx6p21+pvdXIPIR0kVqr/us3inLejbBOhfiK
S+cBOd913Iyl90O3FTrfRONQ2GxaRPP5B7IUd1LMeb7UVv2vc6RrUHVgV830+x0CnIkE/6TNav9U
igKg5ZKoZIffX1JZX+znH1K6dB1TVgSfoFMpFYnsZbL2sBQ+g9mMedwxws331dyfZnabC4u8zsj1
//Kh1UgfXIJqE8ulrAtL20pvM57BI4YVeE8UaNT9cb56aqdGBAfw7L4+/5hTC9KReo83wKHLOjeE
C558nU/bYvh2lCr2ReeXhS5fmWC8UInCMzjZKga+ai39tOOwVDykOBI5XkAWonetJpLhbKek20Zh
tJkTfAPmsjhhPQYvZiBiR55NqJEOSrZnSBKHqwcmVPdYPkcm+RhwtwyfA+Sdr6aK+TCsNN/V5KjW
BaDhX1aLHaB9AUm4cRhXVa3fd0pJlqQ7uwZRVxmQ+cPQsnF43IgaoJUisNO6N0+Bra5GA1w1aG6v
Rt1J3oTrrHTX0Cdb9AKHtF2kIho1xj5CFgpUJJClWsxR51zQtE3VTQyNDgSsTzrz1LyowZvrY6jn
FhKxSCNb/Rfx1ZTTelsPBl2ftB1ORNWrwCWWlMOGEkCkVUYtbW3NrPmKvWD+mmySDooVSBgYhXrd
lEAh+d/OqYMLGZ4OWf8/02xlqQsD2U1CxuOBoOD66Y9Ub1vQ3JZmx+5a3gl87zza/KRe820l5dIu
pe8KV5MarlVpHlSWCw/u/OJ1SQbb+9IsDazVkiU8pv3lzQsumc5oRz5wOMgExXBD9EiGf9H3Op4o
o2o3QlX13qIBsrRBVbZzsFO5FkagCala28RznLAinD2YvJMgEVRzrh+6EN3P4LWNBL6On+RQJD4Z
GF3ubfFiYsSIIt60jEJWIAp63FSfWB+D/Poq3+4svl4b5Lj231+bQfKswjF/GPfa1xBuyRUqHcLK
+FrmZdc+m1PlQ3iRLimEDatFT6GoMzOHLEm9+DHdwbQsqDxB4UUAML1fhbkNvlq0Nsq5cwE7kLi7
Wm9UH29HAhlMBWADcVud8xR31CoFW3vBKXFVpzibrx98dug6gvibqWodxBQri1vcnoCm2oEavqcn
Wzjia685JrAFABvA2EXRjzsZbL7Px02DCqdyu9B8amyM7TeQ/T8YBSk3CK+b7+nokbmKfqeVuD82
lxEW7NWxhcdHcSBaBU+ysCJgzTAQipckD6LpWiG24npelZ3OiNYWRYFOAxbVXUDJIWYPj5bi4qbf
O4SndL5k7o2JvVdVR/S46q8FS7xs6QGA5YTEaqx7wVWvodxkqMMMVtRqpHfHhYgDi2KADse39Rqj
G1noso1Ht+qAAdr9relgJyftM5PzdJtnjwScnlZvop7CyiDlLpiRLtBHZEos9L5xxCdPz8sKqVFA
y5cKm3Y8P9XlznJQcHE8wTINf6n6WYI1i6s1GIFjkkouUCVhH/UYTrwvzPuiDVjk8D/YHV8v2fHw
DHo8cpEU6kGKNx2QhhKGAvMdYoCb7pOtGsK6hbCKqu1b3b0QVAcmSD2DMFUvrAmRNq2MnwdASo94
1deTlQkvzvEL3B8uACIrsghvKueToqYKuaycVcd/xrbXUkI86C9ZnW50KHFhfrjzcb9I6fCIkQ7K
1+N9MHWDEjW7GyjsphcAp7ySMYFFMJJsxNGl6UlkeiN7KkauWc/yKU7ObcuwyhizERlbOFkKnD9x
rokq9NSYY3KbQLPiLQdY6sS/X3rGHYRzFxSsuqe45XecH8HoDAQarh5bJ1ORhUQxqDqIlbBWrCeI
aFa4ZEhL8wG2rAUZ0MJJycBbnnvrSXYzIjcx9OuyGnl69TcHxbqBCNIgjMyWrSrFegs+NbrTsjSw
NeHWkMUKUPRycZZQsfC8KQdC17Ail+sYV+ilb1k/iXAz7Xd+6ze38S1ZrNFeRNxs45nTwm+xULNS
nnTu8g2RUQKjaIO3UK51fwzInTHtUmvWaJNHeEVfV3Mgd8M5yB4ihuOoiwYaAqCw+VVGp64TIuyo
vldkOO3viC/tbRaS3b2E9VB+3ceM1B1y78z5bm3cPhHGtPHlOTCwYJLThWb7eA2uYux3sLADJXUX
1nxxftBJSA2nZVA1cOmuAuT+X9o1jQs0F5s/phAnZqjNTMkXOPSRypOnk5z7EMcBAYbxQTpWbCCP
aY2ct1idXNL931xyC+DObLZZ4hJn8BCOkZsxKmJrkesVrFltrqVsHr5Rmxw4Dted6JNi9OJIt1FB
yJecSMb59Ruq41KC+jFSYmrMtSB0hVHdUY7s1itSLktNF7/MvNJ4GB++fu825S4pkSutDfW396RZ
y4nQUJQgf+zwwjM76+7z1MRe6k6xNPH7rxsZMW6o+l3y2UCKP7mZX6EFzhBLa7HLSp8aWWbSSGi7
ZTgTpOah07Ju4gFJG0cTvuYHphSGnVQYv97Kif0kuY8QwOvk4eTm31XxIDPIE+ouI79yjTeY6Khu
JbZDOFX8bNmbQqRPRNLn5hsv78ikJAOYhMEGxWVhMSz7xgyZztc7tiPFkiht0j/XREzMAxSoWDJw
b0e6mCxL4Rn7FVVzcAgKkPoCGnM0I7SUVUX1JGrcdSQ63ejiX/Shn+uA831/hT0wwZwuQV0QvMu/
J1SH5emLuCseLxeP5nwEGCTqQxoV9VIWs/100yBlu2S4PYk787zVhLXeX4nOP0N7nVxipbQGzxDR
I+eL38s4tWuc8Al0wrYhIFw0Lnunos+dnPg2CJbGY4RRM34o8rCsptleD0MJ9njh9e/Eq9vR5xVk
4WB9zk7hoGltLRpbjWYQeB6LduIn3+guhI2WRnHyMLfVJdky+lQ2W4Nxg9icnSrZqlOoMXe9WPhq
b5VLaSwHI+9KCetWT/FG3sP5smcNhaKIce413RSx3DDUleSRwS0zOlBfnsPa88Kgs8Giu/NC8Vh1
D9GWi8p6MgsdVD3ZBg5pK0xxZBf75L3vifBjHEkGRxL2/0xqR1OIPUEMiffBgrFJBfjyWVX3XU25
MK3aqC1Oek4Um6a+26xA4KOX7oYfsyENrl0ptDtxEgseehD5lSQUwYgHQa6m+gE3zOEpAQr9sXkH
eZePBZAvVgB3KwMdbb6i/G4Q2/XLk7MpiXAvwBMxZwPVfStp6TgGYs4ySqUu92ddl7goTS+grQZg
REPXX1tBL7hypRtyRluTPyyIqqXY1ecGGGOBFNHi9i5l6bQ3+AqDZbhjm4VLVpSTzbcfXPPbYFod
M3P1q6aMcAeDi2B0vln5Ac/e6wAuIp/s52lPJ9h0UNhfmQTCj0/UjU2nmsMKc8HN7vmxfuvbqgZv
fYgReFxJwIyL85AsmoMOI55ktn2/j4ZLAFq+A2yOWo8PhwVy0LcPCUegbYeXQO95QkFngyIivuo3
Qv9aK9gJwrZL8J3D/pksq0PgsImVA93TO+zbHa2LjgShjgGYLPB3p4TI1LprwbxB37OTbQwnxxyN
h6CcQWcFvz7iFQBUbUXK0zXPR6unaPgudaOVJBMxu08UyV2izRIN2hfzJW/SaFGyyTUWmSArbIgR
8i1oWSduyfu0fJ99BT1+zGliuFM6j2vxNhiNYNV74xYoWU/kNxVKM6Hd17NVRV1eorfdPlmt6Zvr
opbEzRbpBvTBPWFUwod0YmryYfaV8rJ6Zkd+0RJOMhW4mcwnsOeJh+HRvTSxF1aefayA/Bj/ZjdC
NV7aWU3Pgoui9ql7NoI/JyoEtZM4InOpkQlBGBNhXD7JXb50VY8XRrms7vMEfb+edBhu4wCw1Cxf
RyB03nfsVCxxeVh/loy5qNUp7n7UC41gN8EoDntxQUIhbP2RlvW0Vfqy/PvBAwboEGpk7BZVlDXC
Xj4VYYkK0YhANSeEQMKgnsCEi4kdXygU13Xy03AELLmmW0vgKcy7rSa3Wl4NZuGsWOngBBvOxcBy
wkayC9ugMlv+XyGvydbRvxeZdC7pDIh3Q4OHrg/a+KEnjqfD3pWhElwqGQh2g8LM8g/ZQvwURiiA
EimM+zUTDnQ+zFc4SX0sDqlvAjjIDNeLfd/3alg6ijSWlwO88doZ7iYMSVeO3Y0+vEaZKZxuO73v
WVEYo6zPlbHovjyx5RRDL6uFIV4mfF3LQg7gkTSHsbjyVoBDny5ibSARfVtq2UPZVULAIXMgQYuO
bKi8KzW6G2XeuS4lOXo50XkbrxdariqSR2PAYnqRVxlB+h0bR36b+6vEuO1ZX1jX0eyoDCOMHmGe
FMSCTMTBDl/EpeyJRUcR8PypzOgtS3OwCSRXoTd9N56t1ac3th4I7/6sKpng4ZiqPCvDbHOL9fCr
eHrHuDE0wSJot3m7u/tzpzA0BXoSeql3JCVDCmuqidB5To5NAfcLd0dtgyiCufOVKQptu1j925s1
cTpvRMbt7jxwzPTEJwmNQTO/g89UoSMZUEYalQddmteBFIa2rl4JBmXhJn2t89A8/W51Q5Q6laCz
05gLKykhhIsd0RfKLAUeWJ2Z2p5YJe4HPiuvfsKMW9flkodFRCDoOxwKN0ohquDVj0DAIEhA8Tqc
qIM1+9V+Cw7j7DxvBBr2K/TLPibYNAWEh7nhWUh8TOEqNsx0pbLtDZRp1vcSe+/VjtmwGVHaJur6
QWcIvMQJNaQHDiIr1Yr2c2Ofmrb5R7lfzwOejLIsCZMGnGDeDCp1dmqKqtVTAE/dEs9jH9N3kQ+Q
7xxRqkTx8XqpuezV4hNsBnOVIXvTR3Rez2lipZ79gtqtxFCrA7vTh52iF6c/9J8Kb77eXv/h4smZ
oHYX18/ilRbtjXSOEys2VrY7W9NNvXrh0ZEJYh5KIokIqL7urmZIiYIWsOU8Cb4y0hCIyI5bEUZk
bPA21P1pxfljY3DiKfxf3lmPzq1mD/lpz3UI0KoIV0xoUwGvEp1kgruhmkQzD4XOZmJpRXT0mU2A
c3O3R13NyKgF3oD1l7iZcpsWSGK9fLHrSZu96jzQcCcY1a49GHBC5KSwpMWfCcrXfiRSnSfRnj8l
Qu2b7GD6t6ZWNjqSSnDl6y+EcJxWzlnmR015+/dW9LbzjJAFhCStfW8+cvO+QfrlSva+k5H6NIix
hw8HbM2WgLm5ylpKt0BgLCrBWESAtMEBPP5NaJbrF/r2AFrA1GoYAB18DFW9ZyfeUbcVxlgkvGvM
0AxQ7xM9Y9vkBOWTk7h3K1tbOrwjhwIKPkeaEwPqDH2b/nVJJw4SA92PMNIUd1k9/azMQH0C2dlj
PHWIh0neyN0RFzi2Rqvv4cCpsXtPOcszZrbfNFGVIAIyfEzJRScBJ+DHeqWcjWGVI3QPff1NcO3S
slDSnRUpqOJuv5vdwBQMrB5CCEkiqS/vzxaBIjc5k1ofzvkofvEmawg43jo6H3tYEZL+v7eaCvKf
CTyH057t+j0XdRliCT4o9FhkqfOZSQ/rjysQkz5Rq/gLTRLKbOssZzMzI8US4qIcl4Ti5R39F0Gb
ZyLLSTis0UZ8a6qExDsQktZf4PR7Jmm17A+pGRSbdzGL40bnnG7KiEQPeG050TvxadlI7KlHPjWx
BopTWC9M02MKdjjAzHvNXRJYFE74lG/3Wr+XLtBiGc9uvCflos1H+XzpHpaaeFgheoAhVFWGfIff
ffAB4IdYPpjrVLrbJ4FAkJZ+3vgO2P2T5mBnF6JFEkWci95LqYU7T56pogXhfw2xc/NZ6s/eNiP2
SMZ2w9aKtS8qFUf3lZClA0/ZCQMbG0XMGZNcUBXWbq1Bm16eXa0nAbO6nHOKCTPUm0hE9bUPVKhK
zPSG07chwSb6GvL6UxfkUSm8N70iMzYh1ryV64QiJBAwXKvjwl+r0PP5hQnMAtMU6HrUtC2n9FWH
5XOd7ENnUIzPIcKG76oED2zngWO2xj+/ATTm2a6ScOkaUISuq2lLHGlde6RbQDT1EZPpiSkM0YzM
vqpq48ehNgzUg+2eWBcBJafEOMF5VoFH1J+3cfMEhBxqwdn20yN4fsGAsqmS6iQHN5fyvI7Bkope
TZHtoKgqoN2rLNWq9EYDLZUzmzr0V9IdkjszoUiVKCPCbR/71mL5P0ZrfAueMyG8F8pT/xGruwuE
MXYmtyFujnawWak5d9SmJvFS70NRuMz1T70lL+cVaHQGMqQIWLPJ5LvHTWcR8+Iz64/Tc4ErZMhJ
EdSZ73VcGcI/MafCVhiHti6UsDpvo/6q1ZWHx27kJSxmte4yDHG8NGmfgm6W1RyVUCuTyi6rSAHz
7xrO+Hvvx3XASenjMush+3CtBnsgzykckl/QBorkHlgT43NSlRfKqNSCUsU5/m/7YinEMvDk3uFA
+vhg4qRNUOp4QcQUdqsm0nhW1OB+CsHbLe1Cfhc52IsFYxjs8hwTN/16NZEk7O/SMf7CAVASkkh9
3B4pNBX0+hjDMkaffiEjUp1rHxdbH64c8vc+U+/JvwUsvOlCZrEL269WpUv/62nNYVeLoWf3p84w
RUYO9/2SJ/FbejYT8zPEgzLv3lmx8regeZea2Iq60MYHF+C3qWLnikmuB/XxXaZCZ0xa0U5WydnM
NlTaMLk2ExkagvWEwC3H/a1bYX4XnWQ3byZAUDUy4M8LOcP/61ploBg2TLAPgSwywjxTN0L5+mqf
YLTq3HSyzaiS4r+z4gEi6HrngXO/TuvYKumWn58g+NohFuseP+EL9hdxrBfrEkolkgmMQefBSRSK
sRSvb7SEDJBuXq23GyGn44RO/OCnhS+Q9Xnp2JsgIEk7MqkdJi+A8O0vGZQSso4RBttAuYxAUeF8
cN85Hyf+z/tbtAJfsro67cJDwFo/Z4X72jDzWKove58N4gBQ4kGmWbjjwGN9qiHrvclRUScaHHXK
wNSINZU4OxliTUpbYYJbYf7vcOjHjOMXe73ngI8k6bPP1EmTNfjq4w0D2M+TOtcoFu4I9qfxNuym
Vcdb6IunFoAg4tO0LQzFYbbJfqQ6/JYbXChxiSTO8qcwTObnnT/WL0JhiAAf8symJybKPZ8HqZKm
nyT2PK5mep/NP437oWIOwDEtTSA7JYPNR5ew37IUCX68Is8emcQGzscffONiz7PyrMomlmt4t3hj
PaY5RsfIUgbkuxEP8hm7k/3xdn48LY3MSDUiheZgubty8bDOwY9F6N3bPdnJ4CP1Qs8S0qyS2DB8
eI237ci/E35aE7/qtEF8lCHwnAxjRq0D05U7mfB+t0RMtgcnsDoP1AtrHfnLQonlKmX5w0GxE9RK
8uRZfIlGiDcOzCjqFhd7MhtYi3LYkAaWwHibaCvZF+6K1MFSCZM/ElHk8kiSbnnqZ/BU4GvoMyw0
elrKSHSm2nXhJ5DqiP2DKf95tjYhFmtIx1DJVo3zIWjgE1G9Axjzx8r+T/spAhRG0KjYQ13cwqdY
wdxNDLbBFIuGOx2W/dwf+n6YVD7C2pE+DDldJOpqopMGCmlrY5Wf4y2kcvg8iax0OhXxYEF8cHQn
2dy5teYaNxjAwBxdA/GKd6XfkJ6dnUdLNMEFNmRwk82CqPQAKsxzmMI/knh/HAHQs6SDQqAvae7h
0+KqoqzXbMiJY68U6YdUepUgc7VF/PxWcGODkbu3ZW6BLOKBMpG3ITmSmt7MQdn1yDOSbeuorHm/
UjeK1ACgoabQlWK0WZfZI49ScDFWLiA27EWnykc7iI4WCio0iwsquKDfiqnf/GKYCd71zCYFBRG/
20UrpErvfIhSqQTgpi8GigDLz0Z7KW5heyUwnhxy7tMr+IqPKbFOuzm4pBtgs1JO2x5ctP+HLXcD
iCP099i8UhLrW1WCSUDzFcRazoI2g8uY2gVTYcLhyyDk53kXiZ2L+XqvLPP8wu/P8H4YLvio7yHG
8TYBK1CRxvEWPkIQv5ax05N2PXyNxYhIvbHmWVCztr/UOTqvNajBirGV3N0nby4cYTl9vndam3NE
6krEHN50VLuMW+/UYOkQYnm6AKUW9T0rL/8AArcgfmSwCKSCIhoq/kX14zlw8OMaWBf/R/Pq4d+Z
Sl+VzIYz68X8a5MnyUvqQPpe15rQ89WRySPvtAzMX4+WgU06nJhqS0D/YZLPSkl6zCsqVjMTspi4
5SGZ5NN0YARSKSXxNdXi01YJBsi5kpIrV6nDKunlTQemVcIAmH5gKg3g0JsJKOdO+2o6mjMOwfWG
mevzvIvdL2p7m0A/4DjvJN+OCAn9Z/2WhX6hwXdyHsQxQpEC/HL+kykU1lW3nHLq6mD2WuoeqwNo
DB+zQxDLR/u8CKY7zyDM4TviZq4mo34W7CLNX6PJfGZwes66SDL0oRvLj0VQhghmkkL8fS1ttEp1
/tM3b+ifc46wxqG7QKP53jJXJ0ltM0kukwtLNvYojBMSNi25IrsL07Tc5z9gR1QjTE/nkoGAiZhX
ypjX4j2k+zO8xS7fGYGM1vBa0/3PsLQMnaBR4amAnvh7oqaT1Q8QkztnDdoj2NYt/pR33kt3Z0iX
g20aZ4zuxGhIoR5a9YEceDiUi0ted5yk/Y02d6fBbt7p54oE0394xJgrF+RZ4bDcoZ1JnJy2iJ6V
eVZw+wDqsixMPF3swy1u6zv8+o39MH+/aAjbd6hFmXyMpURM95oEV5x7wiODf+VK4w3JL9Tu2+Jz
OB1CLvOdXO5C1A9x6MxvvOlR/6aIQk3QcoHCIxakRVWQaSnkudlrGZiYDla5WqGyrm0RZ7LhwR49
cWWgoQAGDz3w6O4S1v/Me8VzMsM4RolNRZdaawjn0PpFNQwdUZaWnscFfDtmloLHzIgTfW1Pd/9w
ED7ZNVc5KlCCTO9LNwhWoGtz6M61sQhi1KRss7gplvK5JEm+oQ/xhagvh1uGipIJ35vd21a2uPaB
8cRkAk74s/U22TfOJPoZfqvgBBqZLBJoCHCEb7jcZbhvlBRuD1kl/vsYLhUja+jiQ4G6smNzFXfK
Ia9AIbyZ2PHg+65figkKs8J0pfpFnwJ1ACZShk5Z3W0o8XuuGKtcbqyY58UzP9nEEEp0K77MvJNn
dvD4mGxwCNGIIAvrZTB41ftKXPadwW8nwJeFx3qm8ynHe0iIqNYW1ZHlraihePTSoXO8S+E7vfwb
yOPfgbr72fLqZP9XjsOho2Ec+KXxNYKW1v1LhmQNp2F4Y42JWMSxQSVhjEqxfSbS/XrBlb49sMvO
AGrx49xSOAneHsNcI3nzrBga9xf4PQUwzb/LwgL5WSJ2gyhRh7DL9K/dU1iIcsV2MYy38BCsw3Xy
huUYymuvDaHmLY8DGeGGG9OxJKfZOIqZM/ULqm+93St0BsBc4nPu82yUYN/QtyzwkYukqUhAKIm6
P7Ye38Gcgdu3kbUaRCTz+ZVxwbChUKnb/78d5mZVlltqCcqsL4BI8UDQfnH33LbdIu8qmOv1fg7o
NhAqyESpUQ/mSg2AH7lGQnvZfvxnRiCwuxM9OfwveMUD9jdbir5c51xEj815POnK07tFurUkBL8W
brZi3k2XdYbvSqNBVlqDv9Rc32fZ2BFCCmfCFOOVDWNJWtNGUfUsN5FNP8uaYzcxZq7JCUsheYXq
Rjlb1hF6AJnGuoQNkZyyvfZQWnPJRKlXH/3UaqZf6OGPlTo3Wc3bk+jO4RH4tnqOI8372tv75yzP
d37eL6tVvLSmADzJb7YrTdqLv7aRIATroXoiY5mbo0j0EokvrH+4p6E98AvKn7FUhKXTQ9D1yrG9
k672DZxqqfAoMw+eA2LCrCdEM2gNFYo4i22hP0p4B3ZU7erfP9+VpEDSJxJvzGbVwubSajDhOPT/
r0rbIbiBRF65GZo/g9BSUw/sxmtpxHoRKhr0IaEqQMBY1wsJo0h7wQQLu5L1GYZe/RObsyIw57df
Bhii6/iSyaV6iexZHWt6uuLrUihW53p3QS9EN4HAOB9g8UUPBuLLMqUTs/fs6ihmORZmiglyXjXV
Txy8EBMSpQP+XE/JT5kpKJ3hIlmknTqUsQKYpT8Sp4hPJbCIirl6qbt0zIxImNSKA4hrjpQDZE8P
gMDBNjjB5sRiVYVB+OYYJVa83xmw+kzxdrAAlFHKCL1UTCPCjlI1oR7yZNq0OfFD19IrlZp5kwo+
7FadI/z5/GBs+KzQW8Na2K3sNjSEUi/ZNm2I7RhSDWoETQhOAsJ5tzcnMYf+C3IDHzSjfb7nlNdJ
cemeZO20u1uJlKfk0kszQi8glvBNYKzTfl0D8tu588HeddQ/qEankHxWHv/cRg/cx6fkZUdRCh62
PuuEfjObYrcb2zFfji04QAssd3L4uKzHxj3i9PdeIavXPQKoXP5YyFJkIMd+LPHOFPCnU4jQGb4O
lYJww59TSPGyjSEdTwYmb1dVqiCmgPGmS2SNs4GhPOKns8sBB5ByLRG9dUOmaFSMxnX0duKr+lGH
LJTMV5dgPSpA3rv+X/j9rQ+RR7RAfFlN3hV1npXns6FWXPz4Ne7TlmijyNEThn3Ri8dpIA4g/c4V
1lT9DQjU6+ETLw9r2ebvxxyXhaCn1E1UA1DXTrSHvtFAN70JMpZ+Yl6u8tWY7tM0F5BOtKSG1+8r
2/jtA9xd6EZH+xUcxvKmDxQraHxvjLW+Pfn8xxciKse7s+qGC1PeqWkwsLR25M4/cV2uN8KsLUev
rpZT5tjcgIpylt6c2ULSZP+qfLEH3sQ7TfFE4erxfRHVWCaIo5Q+bQi8DU8upJuLu7jGccy/ZrBm
O7Ke8M29fUpanph2oAR7r0AiKEYmo0p3En8llbYtK0TzvGv7eq4H8RZDvwgW3h615t8kM0ti3br0
LnKCsPjipKMLSYkt8zluNsm+qXwYHeJAEPm3XdGoZNoPKj0yOgpcshpeCNwa20kEoVb4/Mq4UQu3
b58wcVhFC45tkzJ6gto8aPClyof7sVytBVA6VxUBsUNoJq6dQeQCyXIpTld/c5z+tVpotaaiz6tO
m5SWJkCYmF08E3zOzcABKlBZN3jQqUM7uc0JJMeT7o52YquCyvxRj/xar7xJm7yjNtPcx2MZYucj
WhCou1I1RGgBjgBTB7VNHQLECbq8HkdfNtQYeFeUO6qfaOGVQxvwAIyoNWO73EYVqiT3LZy8nX0F
PmOUc5hvhHLsoIETCbl6QvQ5s/1cN+d/DKsYkwSsg3+yZJqrOiviZWo4s2bhJu0Aor/DMiHK/OWO
hOlKC10itsWogcqDu0X7/hgFi9RXfVnUtuX2gBroW+cQvYY+WHwpET4nTvdoPLLf4AQndHd4RdGQ
7icOuCDrePYrWF6mOMTKf66LSboPx4FopmsoDQYIFbsb2cK1iiN/hLRdCM4unJ6alLlxoHl+7Vuk
N2KMnQ9/WB1Pmte65djcCNX2MSqHGBcFhxUu3K3Br8lYaHPSlFiHgXgSUGAkqFUJRjdKGsxlOAJB
73UlnrHu3wXfbMZNp5taASAymhzRk1iQLDeKX98EG187jGx0zcM5VVKjeruiQq6ynNQe25jwHu9l
7nKpn8DpywDkHXCtshxkwt/RJQXf/UAK0C+GdTpQfk3xf3L3taBuRbV5nMR7XZ6X3+0hgvXmiM12
BtRVQh8sm3EiBMxZacjXKsnFIYyrY9P3I3jSw6Ht/X7eYMXvNRrqHaQbMAqHChKHBs2Q887AjJeG
fo3z8pXVw98A0cHyZIyRGGAtexjI6sxDO9EtUoK5RX11LrFR5Pif+F5btBYV2zcuUXtLoXi+DdZK
pELzac807tpSXcHnc5o2RKW7ep5poY7XwhbjvRkFl33JzhAEAK9sE2yRTRTPGkD10iXIprDKjCdT
mV4skaQZvSIBDopSgxzOxEgWfYGRdyALsHcHhVIXavK0WUzvmihm9OKJWxPWmGyXNhzB9fuHE1HT
F8CyvMbkWCoXhOMWpGw0CZYtUYh829YuSM5nbhT2xXSqFZWSrPb+5gjzPpfXDBE7RGBUtSJ4Nb/D
XJv434ltWBAy98575a/tnjO02/GHadj6fZSVT6rbeDD+VH0azBu4Mi/1D9KlLJb0ghSsGgd1tHeB
iJMeo8KMw9XwD1WzNfiVdal3j7+fYeqXHlwT3yBbzQgjKR8YLf/K1ZQc+FSM1SRWKm5rXUpOiVTu
MsUPgW8brjoIRtj5LOz9bPr4EkGF3UisD4pEl1bk0KPnN1hFfhx9wcg3h0k43zMno76LSAs2KoJC
+Jjny+hc0beI2eDAbTcdeaVW0FXyeKZDKTHT+0gS4y8EQb1eCNxhvn1Xpjg6ENYtj7A11Y1/D5uR
hPkI6Ov5u0exCOXdDAFzd+kcSze0fYKJ0Jw7H0wvnDdYgOaCmt/v72PUZ1UtueQjtEXdNXPXicIG
ebfmcy9W5Xfg76iRbaTe2+FB0KBQG7bv+IQiOdMT/5SPhiSNdt8IhAxc5KNQilnCBalK+kAr6dNr
CMsrljVUs8hfQHucpqD10mJtgNol3nt86JoW+tFpUlfrfOjNIHjdMHWycAkv4kKW9gNayyKostdW
P/qKW7i1/d2e7zWTPDbqb5Y/XaalWz7zyNR+dVyEcGnAkBngvRzPzhbYMr4iMEiGLPlLHZBxhYgH
+V96zjGZcmrW7FZQuWvLQUyYuWhx1itbUcAQx2m4GP90qiAX53Uz/Nh5OIcae5PYF50mRXz3B7bY
J/wZ8jChaUYW/qllUrONARW+ULsCT7SnMFhgduNUoJkRyA1TnaRsiykSJKGWjOZuIeHJxLmVU8DY
gTqWIjdbnpbiFLKGH73eO076wnt7YUchEBwEa9jr2rCg+geWdEumM46QP/lwnD1beNYMB1q+Cp+Q
NFqTG32f9XnyECiAGfqqc93cipi05CVxgL6bhoC6B+Hs7plQzCZMwWmdy4VH62qSJYd4Qv1O/g+/
bH8FDlaX0Sw9ZX7Nh8HQylF0q3PdFHv2vzJgHCymtUK/4FKG9CoFaN0TmQTJndzbHZFL48/haxif
SMWxit5ZwwvHBw/717PJI8uwTXSf0cUrYepSLA1jYQSp4i65koGRtWqxlOtTFM8iOZjLnPJAQkXp
iWp/8ZK/IIQtUw0t3Tc53w73hnAZHIBt+ud7hMD7FgSRqLTLSvawmNg115pTcA15Asb+5/8xx1nq
fl7bhZDPyTR0OFTz52OPHuzjR6XG3y40I00iP07EGFZHNI328PaOClv3Vm5u7h/FzEWdRePj+dd1
cCsiFZA846tjJ7RbvYHCbOOxz7AsY1S6QC6vpYq4ixQUjrGbqAumWuSftWoGIb3OMonQYfPV9KeS
gI7yCtclulZTZ1Dn35ZVMHYz5klJlYXfoKS2ZngtZuQ4FbER8/zEcI1NttHBBnZnf4+Tzy0k7RCR
yoRpHiQ1tYeScG6RPYgJrOipMfVMED5WO2pXuLPOBvt/Fpt8JUTgKy5A69Te4tuiV6tnyYV6rF07
QqZ5DeYipO7sGsTKFbGEQ9GJ3QL855NsFjC4eWiZXvoQp+Jy5XezMVk04JAMEXsD9l0MdUNQTiVb
swYOIfYBRnQeBF8BV9C/dSOuvLE0Bzwh2Je55+r0lF2/JNAyEfPqQs3HqJe+zJnbZfK0+iLn1dW4
G/bLl9jlNgeOArAL375KCkh1gWb09MJMEaymHhW26z60Fh8sDiYZTDVtj0iSLOZpYaA4sj3rfHdX
8ayA8V/hP04/o9OpA6pPBbER0brDsf0P5JTnEG7I9y2mfuv/nR+P9S3bRQvU7S5EZY4pUndMqpL5
I1NhzvADescWI+qGkPvkhCoINNarr90ngc9VdXVgldDETdQ2+VOaGM9wqaUC2tdk2gocICM9WxHx
MjdpGMOUTVSef78vpLNHJOTGZZgGtWDoz8WMOQu1dU/3Ak6zQF+VwNmchxBxR58OhlQc2V+IWqOs
k/2nz5I7wFEg0NWlr+GeYIbCqo3KV/qJkNQccH37XbpFp6P3zGawJR0q7fAmWHga5QE5KAo64YHn
NQEnwzwLgEIadwHhNrXXs1xmaGJeAqSbYOR4nDCvATie+dtvo6kHZs9mJtiAlbE9/USgfE3+bKLq
VqLUi1tr7+uk2/gp1veYZvrkc7EEgRvSZkDJYmEpRRHpvC2jH3OSlG7h4JS3mynvsXTiA29l3EYL
oEjEs2iChSEL/f2bGhwNk8jsfoPeMcDE+RgJk2uvIEXlmvOJewtbHoa9jznWZNT9aA3aV4y7oxXa
jiZKJDxFPd2iAlhm5+OF241eN0Vqr6vqI6VllF4/OAopyfsEYnEFJ6YALzxMlvCGPRV1KKMAaTny
qv6ugZ6GBAi0BQU2WQ7Y4h6SAygLYd6qHCMpN2PbdV7JoHMMW4v3azeod7YFNXczBg2hm5n5qbIu
G7ZKIBVUGeeciLFNQp84zD75YTMa+P1HaKSLuQeMtj4nD6id5AWl0tcXuTyesABcGkAM4BrawAuE
kdDKVJwEcJsudaPZUDKt4r3UGO9ZgcygF01Eiw67jR6UDZcv2xkZsL9aWtQWFKhUV2+WurcsmGyR
9LCb2ZuT1w2mfS2QQjiC3TVfSdrQoYV3qGdMRYflArGeRwPpRrsdckesWTEXFDdoSYGcQd123PTs
QlcyMOQZt+p5HDwK/kxan/M/ybKN2cTphK1VCfbzyC4seC0G3lkvGmEfz2dZaurZt1G22YlYIGcg
M4XRFOwUTdiJXPE2b4C260MpvjtPY/gxBUVIymneU2Vsom/JTMggpZYuqO6B4qq0Eag1qj/VYHDf
/IujOxsFee32Zl54RRdkNiDzVfDE0hwsna3RB3cMaRGVWKAjheH2ie+Dxqw69I3/a8qwWwNgkqzF
Z0aMj42w5XviSyUKsShCUMY5Uh85ZPKk0cy8HQN/bFCZkD0bjB2pp+dtBxn0ovsNInrkm9jKtXxh
Uprc1VPnzmopdDaksY1u0eZCrK+QMKHGJ1SqfhS/GXiS5QThLcusQmqeu3fr3yNc2NWKFUVlcofq
9n5X1YNYJs80yErmMevTOwO5ppatKQWnCejcnHTZonvkwGvh0vtil7qkqF0myyICd3/c5Ayn/XUO
a5hAeaDchHRJqGRvlTYDKuhUn1bLZAINWBQ0Wt/N7W/3sgT5JmlK/lwN7WSNOhIJ4hp1l5tCsvxP
QEPS0u8RyKbir9CEgn01cO+tzYQqUj0ATzP1fSNWTreuiymGlUd8dAtUNViBqeqOcl69Rm0xuK5k
xN+e3BaYNEqBHUWs7FQcQugS85Kr0XvhyBR2gH1nz80uecQaVwf0RzEYl78nF15YmPqhdSXjIQIL
JNeXslLCtCC2pvX0LLMdiWD0leJ7RvzgcRiIhrO65ZB89nqOztAl36cKsKJXCsd/lr7hGQDGRQf5
3bC3yNRMY6eviheIQMHkAaW6g4oScumWnywvFhrJfKmF/91pAcHxr+x2U29uiB9D47BaNTjv8x4J
Qc1D3lC9CTOi9+4vS1FXtcBFq4sXp2et3kghTRrbqCOXFWaQcJ/oBOoXZn8Cjv7Mw9Bd7F3Ri53P
GiKtMZv1gjwU1+2eVxWV/imy4p1oiZ7mDQW1hnuscHVlTq0N6z//+RD7vRDUQz6AuhHdNN76Frnt
OyAnoHCZwORypweIm688R4HHtCcK/NlRi5ABqG/o0riZ1OpVN9dsMAKW9js1HsMK/Q5wANQxzt15
lPk3O8xh2J+TN2n9/hXIxN5HePQPHt0j+aB5ZgDf6Og2gArANNhjgLJ4lF1BfTKUPK4vdM2Q9ToC
ux2tbcBIc2VU2Ph7mLAvcblkSPSHJFNmw2Ykf64KCHCqt0MEokstV3I/I9OJpaCqQD/e07uN9Y8E
+R9RgwpHQpVHvb/AtsRKNUzemhX52srK34IuwafHz5vie0Onuu2Mt1XoKC7t+53w1S7hrt8YQ6y6
K+Ziek/NezOwjQ0z7nTUHuMfrDjWCDQnzYvAUhLvq93xDNFeWjlfAlBz77qGLZEZyKEMgZ7i3+Ix
tv/Pk5CkA8+EXz+qjXnpRLd+CW6dA8/GKPPD5AueljxY+loobqKU48anznGWv7Ewh272ZY8SWrle
FqlTsyIkKd8jj8pthSv99oK/dGe7GE8WibA8DzELi7LKL+fQwYfAFeamrrTOg3/B6Jubfwzmvyy3
RLUK0JeVjvy2ETnD1oZZOcw/ow3lkgnFKGxCwN7yXbUf2Ifztqrnfr+1Sqlvtkki2zEiLHrwSLl3
lR9Wm/esfNZoshdw+UIcH0rShFPHBqKrkHVwNUtaucVJyKs23kxufzTEgfi/86zD/A6Gfi1FRbfT
ALd2YQhKyfqFtGTq1tLGmDTLOiPqk25wPERtTnHlSoTbXmorExoLaOPIqmkgMO76wQaxfq37eFzy
Cg+RLt5DOuqm3Skjrj0MlS0rfsx2IFt+ah+SSmazzzzNbHqzji/2qhIO76Gt5fPdh8xkwbjxD5jV
WWD2+bzIvpIPOOFbeNxsahqbwFhhNN7jdKXA76XBx+wlSu/9YjiSRT/EiXGNFaDx9Ieo1KfXPOHm
TbdIa7vfU+GGjkYVtGojWV7z9olLLX/pOt91bP1LQoAZPS47CgysonseC6q/xceo7pWa70GwClCr
4TEjk6WYZMA4E7mSyvcatOVN/Ng4KxYFss3wNDFusOL3vDgpaLJLiSekK9xoODggUncBsv+PPYMs
r8n/ESYoqf39KvzgpKJR42uLIowvhQUCKtWbIXaDXfOlzLZW1hXM4MQ55+UiH0gSHTDykrnk0cpN
FhKLS+sTPN4pdEgNeM94g1GBrBnIvpTAaDANRVjx16ZovqQs5FF5EenexcphIkjj0NhYqeCNzp5R
9swQkHVPPcemfCC/WQkD6y6bpYMpkQNSgXhD+yQRwJsBfAj9GxwBtkKv5BO4kdgG/8d0vYCKq7Lf
1A6WwsvSesoNJkeK/R/KoflrZNKOahp+P633X0o7K0PAiozdVf+YTgdHptpS8Qw6hI9ABAbQZqNY
SA8BdNiHuHWy1v4QOQK3owGLstP49VcB7XuV1maee9Zpl3mTi7w7no455iNHF71TGtHfklNmLQ8s
cmLpbN9U3xdYQZB7q89BTmIhRvAAPwi5RN4wLLGWqsCY/5ufkdjutAs+PuufRIDGtVc304QQltOG
uuc4tALaUpoysYtxIVyht0EZwbespK/1YxZtb3ixtkkNt2ZjJybFNbPmjd76P2SR1TX22CS/NSmC
q4UMZvwECqg4jcRmy01PBpVqYvhkYwREMSTrJ23i/ZLyT1l+bYOezbJ0XXIcM8U/TS5XoE+qEXlQ
29J9UmBc+fwRNBkV3ql7yS8/Tc6KAZ/apss8KmjFI9jqNkBMQ+ZqM99V52Fdt5bNOpx+LHpLalNY
ZpRb1ezIUciZLNVZUcKkmRRUihp2XZD9nkKtRivaTTWxLzThlgTtPGo0BYv7E3usD/Vo50bSs3YX
QqQtHj8cNOEjMBTmVZ+C4icSM4GuHUcmUKWekHQRtyimE1auShjT3inrmanhgVjedK3bM+k/zfOr
cyDLahfmXiMakkPv+vh8jccDgfHghi9G1Jtc+iAkN0RDBesZnHQFinPmvRHWNAMsXH33EKdGPlxG
H6D+WZhgCaWcl6xYMukUgM+SFJfKnew6eCXUczLN5H6z20oKxEmZ6wuuXZQLewwJKfRL8HT2rsBx
GRxMZ8B+hWHDgwSuWjNvF1AN8UnGVHbh2t7zhqsqepZMFREjlLwfKlSdpY6QXWp05TeMYsATjQc2
uMG9JfPbdOZSVZzPZV1KBELPtGJyYrDo5HFerwnXaQ9tZ7DuSZqccUwKFTckEbakBUvcocpPxOaT
dkGlz8yYok1oHAggyel7fntefvym0CfJawBvP4qIivBcRStuAxrIn+5G5ihOz3yXQPJVC8YULjd3
ka6mk+cEwZtYAao6X8NQ9gxzMBC42ZdqIrKKODHj9AG1ix9W3stBF7fzGSDudlTRCyh4PEIU8rS1
PnBtxc/1D3fIyjFFA5qkgWvUUr532dPli+naHkNfTPjFsjuBSgi5BMZramXeJp5buWQZy97Porrn
34dZBDKCcg9nCzMMDuEzXXeViYT188wkvLC/LRnFy+8sBVZH1hjRLCyZwMNVNrJqqn8OwWMo+3Nc
lVPp9yj8dCpV45skzzFHVg0ynTcwam7M8glmwbxK8iDNk5v8qf+fuVo6fSb6DhT94Hgs3c22owAY
AAYk9EsI7uSJKJKvEosUzw8URMa3qkkUsFuE9+TcPFlMijewv5eDxO5Z98L6v6mq8+uBkVVa1uLb
Jg6EYwtzWF8RRoXeMGzqnH9EYrHgsqVbqR0WkQiNw9k/Kn48WM1VmSiTiwE6bEqwKafsqdE9mdg7
8UvKb0Gx7vH/z7v9AJeEKWM/bHbMi3pXsAQzvokVf8q+L6raFY9dribcTuZ+94O2+4Zs/c/n3NYh
9IIXye7U/LvrFm+eXLQyegXstDQ1GQ9C6UqRR4TpPzrTcFS30mo3XzjGf7m6Vs9p/1ruKEiUo6GE
PKNMJCBKbSM9xMvKRBcklezEp+2SfD9dl/xwHZJ1jhtUia8MLckg/va/RPFLfwCIlgZk/5Aue4uI
kY6ba+AsjiWU3J/JxMMSPH8bL4rkxKla1VNJINv3KuOY9K6spofo6ybs12Cn+ltRy6khvWSDnZRf
tuleMKLB63U7b2pGnwXELVgrJn5AKo6lSv+co5Fj2cSolMNAlu7Mql7wAqyIRSbpg2+93RFvlPPe
jLjfUW+D5onTFJBBBC0tIo8glHnlO7Cnq0KpbakfA9VpU9truERSGx6q7IGXtxdrj6IePTMEjwNc
6VQe2acdm2Vr/J6IinuQhhTHBJ/NJYGoIffYSortUI3ecca/2aO5tbyZE5uE7ijvyibbX80Xr1lU
/QCIWbmnqZXnu37mlg+wn4v7LGJcGLAjhckf6eDdnfwOJWtQV95M8g/2dxWZ4BPU8P+okzYr19nk
hqGeUmuibsY5B410J4WVvX6Vq2/xrmQ+IjSNvwPL7g0Fh3/evf4jYwPBUsqVK9xAWVriSFYfv0wp
aFFU1u4FVyhuXuzvO2PDi9IFZvWv6XE1ee3VUC8orEs9qGhF425CTwQCbrH6R53lCMSSSgwkPPbI
9szhDrLgUSTwOy4/CdknJAnE4ioUDHJZZIat1tVwJPcXnCs076y78cXa3yGC6aO5rd4xVff883Yq
JmlE1fLhf5Z/HlckLZGFpXw2XBTbNf7LFcMbBVR3BKmA4AwTsftAg8UU8mEGVwSOyotG0Z9x6xo+
kUQuT66iFCm82hM4VS6iTNLzQXt+fgksd9cNpSxKHvAS7LDInbnyS5fUslIG9rxQqh47iT1ejXFw
kmeAmZPXVop6jSuZUWgnw052ISa/Q8Q8PW/t2R1BF3tdP6u5UGZ09lK716YEFI7gjsaK4y0q7bPE
tVR6MuDTQMBe8yQCr1C8b7oM2otfG1lRiTlAnfVZYR1ZBwse1om7GA5+ps8LnMpZFDOUuvbjwksM
VFlpL7wDrtjrySWxLnfJ+MBLBtEjI6VBnAJJzOIddEsCAyYjkPoiDmpHiMmPWlerKahlEvCHwSsH
QSivLWYSyoZbK2TQpvNyJmj+zG6s2BTjfWLVDMIp9+8P+pwdA/9N08VqEwLWKeEX+/ffFgbnIg59
9iL9DJ0zzSA1xdZr2fwoNuo0zUwpWUR3F2qbCkFpAndpuUWx2J5lhs31D/xy9YZ5Rm1TIi5BmcAl
cjRFhereamm+LCw5Q5Ckn4FVmEbVpHfp3IZERboeN1FS2T9pvaf4oN62dXnogSUCn3JowOqdZgPx
7P308NrbfXEjBLFGmGUmdwvFAB5p0yegRJ2bqdsd7+NdoPgvyLtiG4wPKKtED74/95jmRtARKTx+
Lne8ubVVkb0yqLy4wRDKTdUhdmTzB2QZqZZCrrmKqCoxseT/9f81M8GCvB8Csj7Fr/WWfxIzw1wD
ccLNF5qa6sm5zv6JWcsgb6kkIsQDw+++aAfk2fb7Z8Dc4RGE1+9nVGLqkz5XBwantIjn+024U34z
Ky/4bpOWocu3PCEoedafn6fPkGcd8fwvICY0nagfoccOklRowJEwHBfXVk+qLcAoywbnwoDspY7f
CqTv0XXwsTKf9kTpVv1MlpBZedzLnJt26ItCNvKgF2fSdIxpvSvSj1rn1+bNYKAqzfl63h4zlncj
xuQ8JTaYRG9MDuwrBkCy/cIPu3CvZRY87TjtMc2WDRquqz4f8gy/HDZiLY/eiDDBNy2qwXxx5Ykl
UzpAKbd3Ev7x1uBcKtETEo8io9/iZAnDJXyADUODJLa7VybVe6+T08GtIooJ4SSFlW4RGcgzmmMP
akrkUBIrdc3SVGr9YFKlQIQPbeuyrcBKabnJtTKjKKryjvKZAAItkAgNhM0DeAwoSjWcLjwwUmPy
dVf6+nyMVQK/9NS/pg1LVONDT5mH1xFmP9kNSRita70oR+moziJVXbugLVLhETivQ1rMIDeXaCYJ
4cSuHnJEQDd1aHnkhv6ayhxy0fpzUNvp+e7cl6ld6LrQTOcD9sc1WjuKT/AsylR2e4hZx5wnLZ3l
ADz/lMEvazKLMEdIkw/MHocvtOxf4qCfHWFd73xpVh4WtLoiSbGLnLmSxHCatnOjaU5G6dHeJRX/
m8XtXhm/1OrAWJQtCLQaTn5qELitt7ZMZKD7FyK5RT10E9NZd743fBxGfScyCYA/1JPh9cikiFqz
VBADH12moyb8qb5Sig07AwXDUV9gAUEZz0nA+4+fdsFEMAlqQ+m4XkZ275jtvuWPaKZhPnYPO5UZ
lvoJl2hDunir3klP2aY9rGXUrb5CM/hRtrQGjPocITCCIZUtTa9P5QrWmYYPAWICFIgvenImsXLT
62Zy/f4++kn9+eS6fB6iVPBvE+DkRBfCrHw20dRo3AgOx+I0jveoab2xAqmwrzrJIk66OA92CVm1
pYof/x5K7cMAzb0SOEAJ+lu12+K3GhPhZO7af0FKq39ZsW/1bH72rtFKMKmgeSFPZXh/NUI8Se5h
/5xzNiLtxZvYfjpRA9N4HTOV8nNwzZI7xcbYqIkIbhUo8cBP2S6ENImTI8PQz1i+bdZaB2l8JypY
LrH9Fh3zzZO6TQCa3UiVRTZfEGABM6PYbSEE5PcQLcXrZp5NT9UV8KXlY/l8K88hwuxK8TOVVL05
R9rnuFnvMbpNjgAHMvFEIV5M+KFSRxE6ye++Qf/tuxDbO5yDzB0bnFdOS+v/4u6YRgH9FH4yq/nx
7yIp9/tjxs8QD5SOuYdrWf19fYi4SpQX9VDz9l6qmSffVf5GE8O6X39IFZ/K2JdKf5tGP0gH7+Wt
VKapVRpcN66MvCSRnIKeBVXcrVCatuQlvSHeVV7P7I+/GRLv/0RS5zGS0ShHaDciELjISSNTg3e8
TCQzDgG9scsexkX0ZyAtES8XZClyCslgJBOP9AQFUBtkc5KmCw/rQasUITc7LRHB0WwH9Dx1RXZ7
OJjN9P8Fj9S856hvD3LkOHGbdPJDdpPKbgaKpVo545FWN7avVNqGaeQtp3C9EHxYAAsbU5bZ4chi
kf1uv51qNLbDaxpd3eWRmx8CGD5p4EseQHzILLKSVM1o01c3TrjwuxweejSDuRclb8bUqzoRcBjy
QbJluM7JqgLx75MIC8ffpGLS5QRFWEQ/C4F2T3jV8GBn/LlFdC3jPRNvELpMJKiR/rRp8C34W+gH
f+AtlIDfKlCd2owB4DsO+TX+DzRLVQjOO3ox4jpPeZXZfqPPfELb9GIjCvPjceghn3yCNmqxzsGJ
Fm9IWKvw5y0F7oVjZNBcdjAN4r+BJLAP+HM6QCfaPsLoY9AIVneqCQkxNG62fpB6CUSkGc+hh1IP
rgFQ4JNJCJZM85f7HNZyEczBwGgeyfy95Sqv+gN6IS1adZ5qgnSGC4DyCRRn7Fp/X3qrFe1DBbtO
8q4PKYRBuAWboMHHefBCkUR+S1DGoXbu2yMxD3PjhHZOIq25lq+XzbI7J2eG14+AHnrHqucGUQcc
fZwEg9Yy9S0t9bAsiNAcCqKUqt1DvhaDlO/8tfHvH+OCetyHjrlKHahg1R/UzlxUnxaeCpNwX3CQ
ks5+zV0zowUufF9U7ja7whzQqyHEVm/8qVxprrhv8E0xU5M55UjMabewgM0ZkQJz4Dcy+1E+Snig
x5lyLg0f/y2bGsqsCZweNM+nA04J+TMt3At3lvn0moalydjA7Q/pDWFZ4UbZXQL6UJYZpdCzkonN
aY3GxJusJ+3sMqIw9SNPdGWwBpvah693tEfXrL6eNDC+8jPHA0smT3Vvr5hIV8IgZPDSr3YNMEOy
XNTpuYnpFL0uyuDT08lJUZcNYpBR9X4lFXNWpMI6M2/eyAXdVF9MFjdxFHfS6roZEbiE71q7A6SA
QDeBGbC8cxzkXZ0DCII2GkuYXePGU+WR1Fpv/Ly+hYtANIJ+s1SqJzQez9WIUESEJV4JhSF2XM4v
M/h9uQyDtkg7T4DaLYv+SxDsth7hVRondZcsMvYp5jfhyD+dzqwTDBtRhP15XtdYkgi8yRkY4Cg7
6tEb5quNvx4q5y3KEEznvph1lazntclxoJm+2hWWn66wKehBj4F/RW/5LOYdPs/3DGLBnYkd94E3
HgM7sFHCUbY4A/yGRDqPikB2DBmpw5eSyJyJSgwe3tZf7vMuD03sNv6Zkg1OU9t6B+yYINKlArPq
NrbBWdIS0fxjLHcNtoNWgavM2Y9UoN13kUd4RKCGby9jMJvzI01/AQyzuXMYPzBIska6mzWUWvXP
f3o5rIrkCSxbSe2oOkxTGduU99YVXOhEJW1vLCPFXevUDlTR9qEYcLt315HE9PkC+57tyy01W6af
7Rt2EMBulgjp5GrlQJQiV0anrhcb45CS5xUOCfB56dpf5lm0fl15N1Hu/TQ/u5l4SfHfynJX47aW
++w/EImMKeXT/pnlyP6/9cdWjELcjzzkDZUp0c51ql+qoezahy8B4cugqNvY054ACAOdKu0GFElM
8hmhB6tjR/SpqDO3UGxolwfiIdBibxlCYGyBiJJlW7dUkpQLDlA2FvHqnEH+jit8lK2HlKzSE6X0
2zzyM4O2JFesG86n5GSxY6w0Uiz525zmY46Ay8qg3lsUOk8nQzyXIUB8KRLJPi1mM2sEixMKH9wc
5Ga0wQpDsIrTblBCDZZ4Np7vmXIf2BgWu4XdQQlLSyYOiEDNarwO3z4mfd9cVaSIE9TX0jCr/Av/
xsu7J4rA/U9xT3IjtRjOZLhOcQSvvWmh4FLqfYNhbvZegIq3uWOe7f0Pri7O4gOTacPCOAIteAAz
AiW60pVyfg6jVp71d/fRN2K2QVxP1338PYhC85fL9bMuNqtPyiuGWbIHnHYebXgm9h3/bZaFHM/8
B6D+KtheolRLlDnlJimddb90slxVvwRbyfkPh4JMo3p6d38ErIIxTTe90ftiIgd1hkdiCRFXbcuH
fFOleZ4nHFC8Qrz97Be30PDWym0eQWAWjNcKT9NBM4GxmHMlfyVi7ep5l6zB1ba86pUE/y84JTqL
F2Y1jjpXfDbI30wFcBSUCELg1kK5PRImVkVx51K9GOQqXysdB0p023bZUpNcdk4Y4n27i7D6x7M0
AxorrqIxZJcOlJAnOoch/Xg4RLIf1UAs80P2DWBamAm1SpgFpP3e4rOagkT6Q9xaZzq68wSQn0/B
Oc3cDKgQ2UgGr35xS2TKlWQU9nltvSzO5bfplUmsz4s7cI1MNbG9zEw51jmrkbfEioUyPwSpXt/H
arWrs+XKMvmYRXnByMS96TY5sDsM2/UVy9xl7Wm/KznbapPohC3+RNf/4vh/Ack+DgnvppnMPhGo
Rjx9nb8OUqYx/9VJ7C/gdMFkBH4lF9GudHtPo4LdmsjGm6Z9DbNmtUJBMLZV6dLuEMgDo63Hh9Mf
PFm6HWjL7LuM92zwX3G5P1Y1eqVc7V/Jr+x9rd8Uozp1/qh+rzDqEc5NF3IMbnA/lVnRcCiNUGqg
wh7tbdSfoA7t603zw5Wug+zEpDM1m4KGsMB60ViZ5fSq8lOlfL4sm/vvhOWaVeoVbObTrJWlzLcL
qz8xkTAKgn2oVQznLX4c5MKQuAraN40Kx72o/80d9tgweRXnlXniQl3HGFRQCnaNi2dLnMY9nHlu
L+/y3UA2o9/4w4ZV0iYd8jHY2qUTZ1lU49ijThmnJQ0zCCFis9rhFk3tVvFUnyR+LXRH4z7BloKY
Iiqdy7WGZ58RcWyECEXAoQyibAaZEhE+fAiDUvxP79zkyWquotWwzpyj1O80ukBJC7Mmj1IhzU9N
AVWRjFPgoGbVDmdk/VlXBG2Gi5HXWSYzOvJoQ3THNfZseeqtYWt/qk2ZKSYPcf0WgFFFZjy9bwD1
sFdzrUi1hAR5D1/Lo83NgUrmJhe1hG5VX7Hixkyekab3YqkXrRK0gn6jyAGsOMowX0ZP8/gU8guY
lQzKOlYdD0vKxGNX/qHwnK3BI156R3qDv5bKp9ERPsHipeHYPLz5mPDfXufEFp28frtV7p+NWJqH
KqpF53dQAqTH/TShRbEaCITE3sGTIKAuHz3zZJMj8JCfDd9vJ4k4XH9sghgMQv0O/9GdDvW2esRT
eOAIEHz3EJlR6rFnpS2l7xKM9vW77igUr1nKjqIhBGodRVUVAVBSnt0bp5ME4XoYed2I2WgfkRGv
VniDr/cC5VAJ1hikW80APeQbSsk4bNlqMV0zndWWCAASeVbHWV6KLiXpoMZMNzyWJj4NGyForuz2
SUifRlkZodX2C0Cn9zz9plPrBwnUBGc7yOebZ4ZOZOUxHVbG69ybytz/TzBoLc2+TzyauKI7yLih
JDCeuR1CQWXZ9nYqZrBcoBn6Ww7ufVdKYKCywG5Pnayhs9ZYDbl0eb68anIftmNAORUQWL3anM8r
tI403g+efbDZdyJd1cUpVch5aDhKtwuXVGqznniG3eCWr4v/MLidr3zqEmfNLXhaul/HmY/WaibZ
Hkb9w/5EItLu70W4/Dhc9DV7+mGNa33uv+pKaveG84gy1vblowvCXzS6D2GwDUxhgJ5VUdTHHn3j
n4h4Cb4Lr6qB/vb6xRy4HSdtaqG3e5tNeVHegeGKIlg2pTAjwWR74fkxbtFhFo/UGUCWp3Uv73Xw
2ppajYWdF7fM3sOKE7p3ZJ7XPCS2uFy+RFxuf3JmRMEl12lST1ZN0hfQI4zHQLhaUWIfUGQVqqeR
QGRUjCORpHSDXCAzPG2VPYwms/8EfZ25RLlTqW3DjFeE0ymX6/p5D06zY12CKEEgJ+cv/mRs4wEl
Ya7hiVmljm+mOq/2zkpbfvbdlSKb3CsTomPz9J32Ynj8L5kSNoRnJb7qGFCIcQA43N7xurVtC8GB
aTSIa/oi3YQ1Lvmzc2CBBpFfOWMZ3n9ZVmwsA2zDVE2o8Ofh2vjSl/l+VL2b4XXuN3n81DG7D0I2
9hMNanzh0mmH6ChwwT21BDxKoLMBQ1wjxon8Of/oCGC6nyTxQO4d0UbFEOlpmFV/gTA7fv5GgW2U
AmMjHoZl1cSu78uO5m3oJcfi6zNCeftjJj17opI1CB+ux3bVHpNQES1xFC8VAT+SBdI9togYzH8M
/3wAxRS16jTunJ+yISc0obdRZmbQ+pjKAAtoCqJHtzglq7s/puA9/jF/eBMf4za94t4aDr8qa5rM
P7D03TWVnbD0GB/aBcBbd5ANsAAFi2xp9zutAyuAE+Z3OX/1ZNWtgvnko9JRGStClqckfSVFIdFh
IoHt998h/uWhjv4Rq0fNQ1sFtREiVEWzLTA0HeFklyD2dUS55pP0BKDkSLhGoqjSDmz9zjbss3GY
uo5f6aX7bE9bgHs2KDpYTQ5qyoXmdZC0gWFybubc7p/w3uo7JOT2+ZB6xusXXZ/4ShV1y+6MmHvO
KKV251Geu2CgwH5C1OcUHMCIR+CHBRceLatnPvrfcPQWjdlm+OJw8CCacn3iS4/QpV+uuPv8vAIA
635B4hdTx9VeXhTHQTrkmdH8zIdZ6FfjBr6ZgZRbLBR0nylPhmfV1KmGjORe/946sudKm3r5W5TL
0MaIfwl/YcXt/wWabvcP/9y73AXzS4717A+sW8tOC2H7i16xCo++W+iHUileAJsrskGL0Pmrtte7
tNvtsLyj/+1jqaWVRYJakYIxMQ6+uOFI8cF80Bt9JCFkjdpBVtyr0xYNvYhmsgvbzbzfaI9PQ6PC
Ce+otbrBh5FJpiME9vjxux7BLXw5VP6tRn6qevITsPr6LT6ym8D8WEeTnhbWlsMtgaWRprF8pNM/
ER3hA+9P/BeKNg30uEHVhY++BtVUZeYZ8a/00O1EzI/oHdH2syFCISn2NJNv6qY+W1fzQF2nnPly
O3ExzkI13twZUJ5WX0BsiQskSrBxYC13zE6Bk52o3daqHBonZd0msi5xZK6Q7Vl8HxTo7uUrK5D9
wyreVEWc0F7FWvcALlPnqOxm28aAlgh6RmQ8g+rzfgquJCUxY44X3U4g4ta+VuP9vxslW29GoYGz
HehMoCtz5TmA9y4+80O8Pi42pQRYW/PSxY/coYKRjLfVJtcIlnrUAbKt0Wt07gNrfJw4pgW7HVsv
qPXhYy19NovzwTUYiA4Qo1YUVxVR8C0BWswXhlnzzsrXSjD5Iui9q7YytyOzNMsgbbH5LK3GiqKR
V7u6bijO90Kb8tFbhJJ0IvQpC1TmUdeKaTLfgGoSQ8YxEkccsRTlrCbx5SoJJ8ypvRanWQKUDLan
U07Jnc9ppVhkCHfhPQD0Hvx0OSYnRlKUu83CB9uyjBLPE8f9L+9xKQl9BIisc14j45cg6kVBq15Y
8+PxB6Nh3P6GnukPQevUJTTOMcwpAPDhdAIIFNNpFUedgLG9Yf3w1TJUsJF0goqajUNmZUn1A+Pv
8N3RYN9MvAzRft7dNNPaDF8dB8kQf+hsTMf/P5GXJqLKBvirIaI8GKOvRWlGasjcg8kLS+f72kRY
5F3Jb6L2IiaAIzS/XAGYF0Rk+HuTPlYVJAyHeGFoqgQCzU9iD14tSKVyAH9mo4CYG3RQK8ayU920
3Ybb6HJNy8PIjy4ERkdt8Svr8SQIhDaBirn3Pu/PBjHePU4X842xOrVNvrvEonT40X50/SCiNBrZ
H4uNigMOcO/v7/EQpMWaLM125VXA9NS4lsgwvoefvx2ZK3c72Tap2hSn8eHRlqeqYbBK7tjwnlSq
D1frUjsRqFDRnL3lF6g/SjLKG9AF1C/dWQQI7APq55HKmRq+tVe/I094H6OEdKDh+Nf6l9e/t3/P
bdoP8MgAPXm77FEZfCRNGWX2by1hiAIcP2XDSZp2AIyrbqogC3sBbmErcYung4kqY2DcNSjgdZ3L
thDA1twhjKkcdo1N0AdvJIoStgv1IdEpDoBT4+fl1FLF+7+6RUcnJ7aquDK5BA31jHXwyhVUy67h
Ty0ka3e8nVHIHOiWXsW+EdfO3hcfu4PZhxqYyCVe6wELPu7WynBS+fjm0JcFzqEHvrV1PhFjnGBV
ANXCu+0JQ0SqTn45Udxx6c3Lr/RaTCWiU+hb+rkCCPYukPUh0m3vd2dCI+ddVsG2O3DQc0x6whde
ocWYOx4VbAhZcQHTyDEkj/SyMGZH6yu0ROPF++y89bEZlnRJqY2Z9iubhkbC0y1/HAKgejZrqTT2
J8QFK8ymGJSlfmw7usg/d89Eq805oJ9YETlJdMI1iRczjZk2X2c/IcrpXflEdLHRAtMPfNavDUMO
3jYgtwnhyABNDCdt4YdQWiEBdHRIhUgCjkbup6Hv3N6dXwCvjBwdEKVjfZ4ssma+lk92V25Z6Xf4
NgW3Oecztsh0UtG0zalDPL/R+UKozuglLfdF1Z02RvYavcjs59mUHO32GmXSSbu8OLanY+la3pA3
C7avMDSWcnGFpM+ce79Cq97MI7FvKPHiLx0/96H8WGYBcrPQVgBq+B/cjP0aLlJBEFQCJMpc7W48
BRmO42dKTAzEHMgyHPpAwV9S8JW9l7VAXObAH/pZyexpc8KGMKYDjBOrsS335oDXtUk+ZkMpCAU2
EfgE4Okm2B/eDyjJrUOIGEcMR1j+razn/HAgCJdWH+eU+ZcoMtfQXcQ9nGI6o9FGkV8ukoJ8feh5
2j+314iNyX+8QIR7lDICVVnUxnPi7+n8+QK//4DVoQcTfe+4Kp5PE56d5l5saOJ5fRWXdEzQQWZ3
elg84RdVPSAelIYEG2BX5U/Y45akX2AVr6ZYXd0pMDUfpqTzGW/2eSS00G1lQPqQQTmx/q+IZzuh
0r0pUsZZSzrFSWdxskaTOW3C3vNYEjBsxMcdWSJPhFbd+hvle/U33ItV0nGZG2ZVaUpNBuuDuugT
w1d/KySKgWVWNLzGpg5pER60FVe1Cqo3Tvd2p5tZm52+5OjGKqG9FYOBVi26TqIx/L79sDEF7FAW
4kIqIIVfunLyFhuZeXd/smDXEkWmGfBsrO40ZZjpVQYWb0u7wt3HzoHQa0rB0HwyEsvoHyRSrx+j
CsVzV2lfptIppEo+PxNfrBiP8T52ha8vXhz4uQ0+VvyLETaext7LAyEwqQ2upjEzyD5NlFTZRkJh
ljvJ+VYRpLFTf0J8nrUJRELv57nbr2T3/tzbS4NuMThlNNV1MSHGDcpft/XLFHGXp49s1DKCi8G+
LUO/M+hTaUJ16LG7ATBQ1xprlsWQq8o2NnNjZryevlqfnSnUEjW3bnon41W+FTu8PobTqDD5UnCk
RUC3xZqx1LMVvRAALi8YJgOk19Ibpxpgl3aQQ0H1IObznJK0MXir9xABDx1DWHcYapw+uEm6Fg08
Q7qxYH781exJ5ewVhe6SS0aoNpUVkkTfMWTFnTthtUa0a70JjiH9lz/96Vk+MS6uspo1D4m9ZJ2Q
udjs5AggjeipIbY4YfDdXwP+0Ss6Y16bUnHzxfC37XRPZaydFMpHK1Mb3eHRkk47YKLSka5lxpPa
Crtd9flJMswVGBZ8rTXeReq4b4qw5wT+gKtNC4xOBUEGD8kUFzJU1eJ8CVh2ogC7IhoOl5O7hxkh
6XUriEN7I7vaH9n3Mb6K+2cxu7bi9Plq4feUJedkUVi59RQs+eTsOS2C+qe8HtZ+l11ImIZ9wbCE
+m0msOeoq/Z2xjeS2NCqLttBNX6A7p8Xfs/oKkECAJAs7UsOJ/L3W2lZmu8FopsP4NjNx0B5f+mQ
Ftd9tdLCB5KUIjHZvyBvTbX2SQKGhJR0ewAJFxOtWbGALrYpenM+g8usqX68LHruFb8FiL6tiHcS
ovVVsbV3JM113rLOLf8cZnpFuUiE5eKhj11OgHVwUjwhe+hglTCvXHNWm+lQupmy+jrs5X56xeVa
JlFGLBKgTVO10DvO3pwsDTqUEFEGC/Oq0sUE3TiseNCwGPW6q94VdoFWvI8CLNw8+tYjZPVkwclK
PkGqG+1+6TlMb3iX6V0yi1S1L7yxAQLDPMi06s3q9CqQoc0y+g4Mta1XmROalkmHsmQjDHtZsiwI
aHGj3fTZ6AcX+A929JjtWufX+F15zEy8FqS97CiSBDK/EVOjpnRj8s6ygmfhdDP1x53N6gRMsilI
lAbg1FdNyTP986wJBeVv8rFfUqnFvRjrfJVrz/UbFI07qa0GWpou5UShHSZQw7ZtX2ihQGlgmKG1
XdsKOdJp8LFyrvRZfh0h/1b6xrTkVOJvRrZJL1QevQbuqc+p000QP4PzsMVbW6XW9tmwfKFXRcnK
XAilb6u8UZ+ZjZjpaJOwnTbe0P5G9ixJZckroi0MfWn10ONMh02F6vpEeR6391PQuCVd6zR4PyD2
PrrCJA+i01g84pPnT/yJeQrVfzTV9yccLCxewxC/d8Md6NAMlh3tZOGXORezBnPSugA7ULURcdLL
NVp/RyyDVnmB/z6qKqj1nwyjtKxXZc6ZvlRuPtqKWFZ9vQ8DY+BAijBQNconzhzd5J70YvLv0mYX
qrIEDgpqmPEo9EF1Yop1VMdjevawltF9BpKkmQKV1aIV8EoJ1eLXXA6AP9c32+tD15YVJwU5jPUq
+pQXnR4RuAORUNI7m1vKkvZ0oZdKp30nWd0Y369RByp1fq93tIdIxL+qolGAg3EmXVqVSgBa5OyD
5NDnpOVkSqxTL2F6ejbsxw2tIUG0oTdIIqUQratNoRRYAmv3vDQ+O+aoNQnS1fVfhTAECQ7NNNCe
oucVLbyFyQnwR+U+/pRzlKvZgngwNIz0fs6NJUgVpor3CJZWwiRTxz7wVQn4uDQwbyaI4Y+TWXNc
G64dHcZbE3HQzYv73wPNVrlTyIiwpYvzs/bExania9Fh3/XTJVqUDYp++0xEG7CfDj1FG5nGEt+C
Ias+D8ScJUPGUdHqNVkpCUihsaOa/CEY02jqwP5tIxEW7WTYf5Egzb4O/BoB3s6zvV5TuCcHJIso
jjuz3EqfoWE6lNeUkIUSDUhoLnGOnGS+Nk+VH/B38IL8/YoTpjI2/VXQeMSGe1kgMpdnpc1JQWZj
Cr3cq5bwr39gh+kTTmLtc8+aNmIgtl+v6mpQkx4Nz9uEQEWywtDMWvzjpyxngt8hIaowiWMuQ/YJ
wDIrwD+rlaEyx8GMAoVMBksusSaHmXpOUlhx4IHpKBQkH+Xpi9OESYMde1IUBGV7A/vejbwvatEB
NIxFB1/mziCdo2StUNTu9XFCaqrCkUpMm08bLiPmX8jXN+2i+gi2FH73fBlydGtlmejsbFY59vI2
u3pk/K/aknQ+Lo3KogSF2AH1HR2tAXYG9Yf1KI9nM0NOZ/lhwmXUGgE2H7SEUzMjvLCeqhMhBO/z
6/lIMF+7/bSbeu5nFaCuR3y99msRpX/CveIDTdKDcXVwj++fKOECiIpGJ/epAPITi3ZRgL7jt7aM
amZY/Wp4hFmAgBlck0Z+N69kWHDmEST9XAkfh/W8rinO9gFawixrj0iz4QTQSbbOKjSzbUQttD+x
Ufj6d63MJutt17YcqTxvOsNs9xLtGQHqOqW+bMhLSDAwD/FASccznk5pOG1uiFGzlbIh6AiZrDJJ
e3nRjcoAmRAn+PavB/QKUpcbXKUBIxlaCYuHVKpFHeiij3VlQd/KI60DcfwgdqjIExgKAXEg0mbr
/tVhT2umX7XScTYB+f1zV4WuHvfJChIwzyVVL241S93CUSXhOXtFoMGc7bLQBdBPk3N2YEFaDngN
xlgX/71pRSVXvq5sJZhOm4k3Z4u2ISSDmRS9RKY2eQEt1OaVJum3KPX667RfClxCMJewbdmSvbm+
WqXJunIVS/GJ0WBYZXx2Syp0WvBjKCq7dQ0XemO2y7VqpW1dS6Xilvy6wyou4yrAXnvV8r2PyuMj
u0WtG0Ji4lr463ixs7ey6NvFSczqvk8M6nCTYeXPJJAJyc1UoOkjgAvVy0XGyL0bBX9RI8dftP/c
yIEW8Xk8SS9AH8GpbbQCkswF6snbRzA1VTmBvCR1ncomyL5jqxVTAtDHZPVxazZIXn7Duh5TcSvm
jYQF75wUiRvOlIwSHYz11NB+gb8N4s7DMGF1rOAECXJMxJE59xKboIMSa6aWo7804kaa6GCq4IYn
7R0wd/z8PJYlsmduusVzYuXxUqZzsWhWlrrwvM97WfETiADW5cG3H8ajPha9M7txriM8GVYwQJzA
ZrG6Gxv8fCuQzphXvkUwC2wi01uWrItODUU0uZP1Kj5DWB0WTdO+falB7m4glZbxFKwsYJ99YyqH
uouoVJGXK9DZGiQYS9K2hNdHXwXZ6fmwxxybd0fk6I8bsoL1MyW3xOAQdraeP8y0BWTRSUlZoT9Z
Dl52ADGxIUm0O8vJAh0f6sViwxAyYx0JuiDbfzDIFzQ5bGFTX6imUlyA76b8+5TtjuvmdMckb3/y
3J5qDlG9juxkCy8b5gziAulrZeUs3MJ7lgEEwIlg7Ske7Ss+JsvqW4dQdfIYJ0wkX7WTAdA0wNIy
2lW5Pzem7g7OA4/yzDZ3lNmGK9TJs69d2MrMfpnwSNjCXOQGcZyTsc1CSvjoUAvRMdX4/E1d1FEL
InNcbxnsIKkrZHwkDT2P7F30SR80M0s2lwGL9T2zf+ry1MiTL7OpGvdUu0UKfaulXRWLYsU7tcME
RdmL1iJzrV1Jmkr1aut0VqZkghp/M+UgweSgrSPReO74Mmbv0NTg+/VvLUs5HM4c4gZSvGk+kuwo
XHzHSvN6Xp6wtuOliF50+EMva0kTkmJ87DwGBQgjWhoqnZq46Uxl15RA+emSA7Zcy/UXZwL6ujSq
EcG3SznwogVunjogr9eQp3z02YPOddDv6RMbRRu07yWouayqVMKH0SdFEQUt/QdPAVnQuDhqKWRO
FzxZa1uKTRB4XrL6zB2YDZJ0fmudU761k7Cxkbo5eF82A88bGRPAP8lEnZHuxFsjAFytgz6P5koV
L8jhbVd0i6h3lfgnbgQ8XFIL3rAJ5TOklYHGkdB3hOxrnjmAWUI2QkNXCcCHW8IBR+PCFoIjnGyL
mDhtLQnhI1AGZlu+eRXdQH7xigtJfysfvA1YdUdKz5TxfhMxmvYg/nyVV0A3XK0A0qqCRoD+Fgll
48ak0xkAc/K1tseHszn+HlnjLq3XsDNH03cHnu/2Qh5Y9VX/NvUyZXeFIc2sg/zA1u7rg8E6iJ2Z
Ia8p31VEyFTRrefIxN8bhBM6Ttv1tgOlGo2M4UQJq/OS5E7nWZ/RVyP2EwLJiQRPJAyY0/3gHtqr
u2bXjkyxZAXQNX57Ds7i8AgHBDKhyT6+1/9+6T1oWYMCa4dBztqgWM8H7tvS1iwHUG79IcllqRWz
ttAhnZIqUiPsDZxxRCZ/GcH6kSI9pXCh8xCiGbHlojoS6wuHFMFK0i/UZVZ0uKa3qzTfkSzMAnne
Ic2Tdn4jqX+OoAQX60ew/m/RkcOBHrEseSKFd2wpFLAplEP5L/IxfKJI/8tw+UWzgh7ldR4v/Vd1
t+a+aMc0KMmapwzMCcHjxnK7/hBknolWzS5auu9xg17KIEIPqoMNInfPBwump68AJP94BhYipnIq
cAXBI8ex5hnuOBX1ctkQ9NXJ4WL9PHFYyfx8nKAd/9PlNQPFymf/NEu9ePMEqKFE54mbtRfv7Xf0
yiSN5Q5sewkUwM8Z1d242/XYuFT2aSZaldq83MwVU4UvSt0ioXBLPvVtM3N7FvaYSS1YsCxfCMfS
sk/Ngzg22vsAjBAx/++L4jOhhyzi7mQLIFfTUuVFG8XV5jfeY9zef+szLcWBvxc9hEsBCbBQy2QF
TaCx6axFD39eAKeBvpmGzZRgUcuM95AAlmRboWVGijUrEjMEZjb8fD5bIuRHTKciyswEPmQ/HPtx
eL6yPrTbewcJ3JSj/yqq879X0iuNKAOapX4fJ7+TSOrlbNFBdLwQBxjJa8h2nS2PSzrnL5HN/o2W
58IwlqG71+rhGuf188s/hGmCQV/B+QfAD58dOHiodSymPjqTUmWZIN+NAx7+0ycCa4JqymDGaNtd
zZoUrJInr8l8jv+adimfY9wW0AJiP4GE0x77tuVvuhT1Xg7KYYCBUAxKx1H3JLv1AxSfjQGWma+2
5/r4BZN8Mmwi3IjsmYxWlR60fX/srkuT/UF+bPs6gx+bPrYPF+jahS1qwnV8WMecOIA3nzuBbNAO
jdd4RbIYpY/lgSvVpv9j0aIF9JkBU/Yre04xXjht22XMhjjKwRsKVtGrb/OzlyWQjB/CJf8/18zK
ItFWoSrfC4GXD9qttXvFRCE0bcz+4fE0pxpNOOAiC1+6pPaQByb2mO+ei79C25zvzfxKTOguPaOb
Zr33c/wmKjDKUIkx5cLPUMhASGxe7sE907ma6YDhGogVmMqVu0+CkiP8Do0ZAUul9T5kddWF0Kzg
VdcXzgSbw3wHAQfqSWpFogux3XCsF9iTcCZmsNJEMLc5xiTGkD/VhFiw1mrYq31NlHJRpoOS0kM1
ohPQM82nRx37wRiPZDW3x4qD31DsqlM4Z3wbJ5VDa1ZlH7CDcQHvSrJ+EhqH858IQGx16HWJGDPs
B+5vCO8jrbY84iCSFBFLf7Xi4qApPT5xFcilggTqewO9AgW1SaBUT5qTI29epS5EIBa/7/SrNrUP
paebehJVQb+2HVT4axQ0xvHIRdbtikkMWFdtrvDNF7G/KvFBQGroBAfyOmBOpVjSrX1/aas+QdvJ
+iTFPL4OTiVxTetOk0U5A0GZl0CBMvZrJEQVim8oSA09PB7awoPWZk4mUlM0QpschmuOyVVwMONk
CaCMuh55BbZqOrTMSPs1SFjOXWQFBuWTGUS+enIjciGMQUKnVvhGWON5bAiYUbEvHHSZYk3dQK0Z
hdrtLs0SgQUezdQRWsTQA8IwYNFZmB4LSF+j+i8eaX3JD7d/d8q/sqpgtvYkNhG4H3vOsgD7RUP6
rAkjhfNwlQWJITnJKbNTRAm0BEvHweXBo7WjNbxqDRamYOcgyeV8IM7++KW3ba3w9ONO31gdwgLF
c+H4898tmfdnrGDgqrBvbjLK3ma+2ur+XaL4H5NGYBXo2TUhpzu114IO3xkBBUYwj1kfV9IfTYcK
x9N9Sts7WP2ixhKv5egz5EI3kloNj9dKAMxUsIK/FgRPhNQO9O+RMS7eLUwwOjqecATz+1BuXdIh
9FB18jHIZxQoAocFEmWGWpCfr3NXURW2BjoISgTBlFfe002buxF0TyhQgvtqYn4wqQjY/WHTlmUv
ZU8uKFhJpg5lYZ3ikBDaAraGN+cxDjZnzk+PsD4LwMNj2mnJ6LNpVzxpjKkNDCmaHMDk/o0FPgo4
fgTFAp/S7F6KdSPxUGzVjEbXL2ETuo+ixpq0tElMZQ1+nxZXLeDccjcGkieKvDHLkCk2gfm/rNpC
7s+N8kIKo7Ug6K2u0VCzFyzEjq4YNwAdRzmwj2H4Wjv6Q269BhRrAQO2BfMN8jvn5pqRB9UxKs+j
IK6KAQZLwlBd8LIftxoboDU5H0swiVJqXtVRNLbqTUfWW8gVZa66nSA2FbpWt/UykkmAvEFvK564
QiUms/t33Pr+NBMqgKbax4ZaUrnBAsHbQ3tGAsN6X9wFOsCixpxBQ0OpT9LDKbp2u9vN58WdHJDK
Cy51GguzPpV1CyzCkjxa+isq4P185DS7nglsfr84AUxsLSBHeXHWxVH0ScFC/4GlF5k2e9LZaRT5
EJAw+sASD0amSe3v64r1Mr+YlYqRCfrggHYfcq/840u6veH6uMNWtnpNcQvOvR7ImM+ovYe0bYyf
8183xnnFwtJBNcHO/d4dm1/bxfIRaa+VbCKvkmbqVX8NiNbiSAMws4KyjF2UanvROHdP2MPpkSCt
ufbI0xW5R4v6ek6YPgUJ5+DBNY27T8ENMicvzhGX9NyqS18KrpuWdtlTsuhgwIuSRjHz31PtMvlR
zTaLbcDMWZLpGWig/t9aTnFIE2zFdL2H+V5TnV8wM5WIHbuUzHdsqv/uEPwEtGZtmXuX8d9zER5L
VRSe6WxjkfTOcdChueJt4V3GDg5CgepXMiGtt9meNto/soY/8Wct5XoAqwnmdraEncZyR6gcoaHZ
xRzuoirEvxXvd1EGTgMc67r7iqG1Sb/rufoqcDn3ok/kIDy5qZge0RglWT7+bUhZ++Y0xPG0KFeN
/IuteT+FLidu+3laUkV2guk6tpZEgYeXs0/UfKAnf0QHy8s8gTe0XppgGr+uZmZMexEcVowhfYBn
yzGAc+a20R0qoPqFBKzJVuzDeYOFVPA98jAJ8BV+XXkQaZjhzmG9HtIPeVZhxZ1nUMZQy7qzMGFC
Gtn8oW10Ldt9lVEv9w7+Bk3Nia9ilbjI/hJWZmfNfzBGP4EADppdoGrzY+5GZW/m7dT7LfBDRdd0
MYUdgDMum5aYjvB1FZcefzWDixLMhYenQesTYB941cfZkSEL+a4MqwdIs9MvAwFC49F/wI2M58cc
muPyO7h/fRrHgZeKKrYjA4ZO7yJyj5VnJIM+sSxS9TYMNNbxIfEyb0Wx+QmyBqkri2y6em4uXBU+
AvEW267hLMcghWr95Q0jitYtBW+0LSyKjdKyXauJ07LjJkf3/QL79yQeLQWW1RM8HlNEuhbVc/5Q
BJ5SSSMzHQD/Z9eBup6BMgsO/WuA2w0M6c4cfGhE+n2tMrQPKe1TSDav0dC23AW1Y6gGB/Da9UvW
DgjKtD3SP9X8waSs9YkYiCNH9Ld+xS4p7xQg+EbCkvnoqhgob0TT17gJTh9Ch4v0rIbUfZcnue2O
5pr8NQvDTNoFWd73kou6FwRcQml/fbCtBlngHzdrFKnsjS0gxrWZ7fCAEY3RMhvBAjJ6MCOmbjwL
7Con9b2XNwcwP9lJrKnz8EuNMf1zPGBmjfvZrsKPFlbBgabSPjNchxEjnuLa/4ULGb/HlnUQdilP
r9BalsFhC3jRZDf9qnipoQpTZbU4juGCsYtutk0ZHejNPmUZYiwANfgQYMhP+0FZtPYnU/QqOOdW
MUxS4E79v454XrQ7ke7GYPAJhj0iXSkinV5rw6pJLh9FBjwGJqZvpPr8NH2K3KLuV6tp+eohwYoF
m20DZK3VT8zvfr2UwW7XBldhOHP47KZXGPHQZrx2uykFsMtHWRBQaiLPrYkCEXDrmBAIpefXLkrQ
+M9zkP8M4Be1QdUunDOYsyhJFjxE0Unku+IuaAQdmtiewQx8cW8BS0J8U4C3kgcGUXkxHy6DX21i
Aze8sV4SIXEjqTiSEP12aYI5MfGghT4aynEVsrVCiELiUb8MlLMoufTxbT1ELsDAMqvTCFeCRm4m
JeghAc6rNYxl7IEnLw80XB5pS56Ri5yyk0Avh+SNLT4RIgKnZ/63F49GvPqMGGjVfR13zYLCZbg1
UiOSWkRV1OoQELB+85LpP6bmKA5xBY1/eX0sIWQXO8XTheZT4RNqqb0+TYjhoQYIgR/C0oE1sVym
WC4pT+XsD1hZ/Ml4WML2c/zbQfrEMHHgfbzqsFgsObx1Ye6KiX46tPB2pFCMo4M5I3rud3wqVPSD
Q0KuzQmskKHniM/Ug0Jg6T4iHxFjxL0zHFwQc3Ewqlq0BWOglHdAgr7tAHcle1yV0ar8JZKKenLz
d5acicOzM2x1Fx582yhtUGX5FhT6ffYz+AkFWiCPSHvUmZNASrJVl//mYPp0mE7CX7mLfjhdwmf8
fJIX6Jtm6DMnMbvfP4b++Zkibwd7knhq8Tg4m6xOADckX1oWWEk7kyQ66ultoHlLf8++W8pBPyn0
/imuhJsS3/MG7rhiQIQ0NUjkUhG2DUWJ1pRpzQUQ1V/A5EM+uS4ICxnImaxo2REvPJ4KtcpwtFGP
scm/4A25apqD3dwbF6BXRkRuQeLUxLDBGCWqaJ+NpalwSt35Oev9xW5i0AmEfBAR1KTX6SzeA6bS
44e7XeErW6ZqA4wQaCGkWDYEMMJS0JipQCzZlyCNnk1ejEmLw8EBSusWC3ZnvC4AQHRa2pTfA0Fx
8OCbm5yxCamEWBPqF9aRXW1hxLhc1neBEhh4mPjWwiPedKzFP/QvFQq0KVi237x6o2egR5dA/vpt
1Gge+PmoE4V+qyGSRKIdi/v7ShNzppKDt12U2fSwmd3aipSIItz+LcfvyzFV5te5zecEQ+v9Wimo
uoFB+alF0Slcs6D0xBIqqlVgK2PAIW9gmBg5yK2oqLllmIz41USUcjKIQ8oN7JiDOvMMEAgZMBT+
rzFl3vcF56YaKsqRCww2dRsW6Z71H+vx9E/uyciiCM/mmTQ/aJdYGOgV2fHedM3mQpy/b8gO6cKe
Qzh5HSYf7If5Cp2wofHSQyI+FefKMB7bhc+5ewx2zw9ktlKdymELPARFOuEeobVX1+B/Ff305Emw
X055+0iyZ+lc89qov95PZFP2dgQFQWIsApRbuyJ+m/9O7jKzUf/VOMavbAd0NjShjlKvZTpweDQ4
qgDNdGPbohnlO3dZ/cnzHhn6VlbXyyV6VLu3ilsrD5k2afvHaOchFEeLxKl8H4n4iBHCgk2VcX87
zyM5fzhmYadSLx+b/RhoesyyPg9YzOydn0vNimr1uqYHbtU8BNxYep/xXwpsmrZHgqTAX8SixU8z
ZTmNhkAHjC4mrhs4+walBYAY/a9VUl9JOZtOlclQmWBdJHGZ8RbnDnEtyyGvZizLWXbK65KyoP+x
1OURLgarrH5pr+2/IzseQ+Dy1/Zy0Q0l3/bcsUuGl30PMMuQ77GKlnZFHyWP1C8YYz8dK4Qjls7c
ssenqkuawA4TeJdu0Fk+Vst+DtPIFs2Rmls/vIRBd3E9v/2WcZN/xNr/jzrSM/XWlSCgvUqiSGXM
UAFOGMcvqaokUay1WVNjgmYG9MqkYUifcGdP54tv/LY210z25SfIMfA2Y8qjHInVaZPuP2C3nPxi
6IO5CUluspl2PlgWNPj9b/Q9Icvz5mkdPohffgPGnC2TJ9SVIQW1W8iOvavvxHGqC/bpaiF0AC+g
douioOAg8IQ53VJhYLTRuP0Mc8KFTAzQHpw1Ui1z6M+mOfR14zDaeF9iiiiNxWXg+RjLUhuuyWY1
rGTRcBi43zB9KJskSInEORymGVaEXcqJTYr/ogc3zPjL5WmVjucOBPU3Y8neDSKCwyIKXb1Smdgv
/hW1kZKoKAfRLy/5W+gR7ROGXPkEL6OHMm7P/7MXGLNZdGOierwtqahCu0skWLdgFz/Mq/BaT44+
UCOzzH5emmepOjF984DPenoARJGfp8x5AdTCsKJ/rTaqJ2efzSsXi6RcXEjjRCpPg6NUlrprHGdu
bLv+2p/YOJll8oulG8IrryuyfcuIRiqxwCaWLxFShnBMK7ZIfJ42jYsvT3Omuq4UI5E0wawL7U5D
sQHPOO6tVoTaExlWBVtnhU+/iArafVD19f46S6rPOzx972xL2VzDHOjOtujnLLEK7SHh1+vvsfKl
WWq1Zb0zY57D0fvserpfsKqWpW88EcMQD2PBP4WRtNjPTwHxoKepivfvNOTSFaYDG7xaCbOPuAOG
y5c6i6w9dFML7APNTRA6oBEpAghACaHBsCzLqJ6spz+3DvRn8IslykACdvLunmhOMIzwCw5U6id+
nes6cbAK/Kd4LteJLTR0Sc26OW1hjk9LyyRCvS0E9HHZgr/XoK+bbioTjyA77NsFPXrBk5Wt65iI
VJDkYbgDdZRRdNxueuNtH8cnCqqmHV7OfihJon4O9p6tqbHzhs3WvykNFe/+smAFmhqU+VbUa9Xu
tYPE4p/5SQUzms25efd8Xr1W0KhSHOeWcxtyVwLw49TcOaUf40dBCguBri2Q7jAeBfKBEMH8BLvL
Wa//I104rfK43lnyl1Fnvv9AjrZNCMRzaugp71Y3AQ5LEaVABdpjb+pcURZFyEXbey907sDTGs1C
BZyk3RwHhZn/zrkOYROzObFPMk3TndS6433brXb7THivqkUJ8TPyRfIzIMdiFU33iz4icdeBc+FB
85bZOxY0/SnixwXQdKPJwg9TvlJqM8uVMqKXicvO7NkVEAAtv527IulLkt3xC0TbTrnxELs7Smt/
SXSAFdZhdOvrQOmmJhdYxpEmtYauZaybvEWeSamVse3b3J+9qHAlLWlAF9wUzqt2UOJ27vdGQYv8
vhUf6FZFhihR32L9gm25LONY1V2FSxqqJUFDlG0dsbj3b9sN57LwDgMckNavMH7nucHLAs/qGtA0
ks3goytWuoycvckZSAXksAv6mq8Eato6tvWmDaXk25+VS4Wu4yfidQU/fCZwnaX2F41wYkZ/NJMP
9/VUy8VfJ5G019X9jNolYqCX+VhkR9eUwgA4+9+6Sf1isaVLBjOCfT5bGXTCMHhRTZMYtZ0Syubt
mpCgWKVGbDIjk4P9DHf+BrdtY6abwB+LU4GQKacqsUj9gnfQvSFEoUnZSopEJkgWtCNe79MReSGQ
wneUI02F4I5jewTmfHkpo0e3Q74/vwWs6UbUGgyxiDrB4E6U5/Fup/9IG+zfwGLojfo6gF95dYKB
q6VrpQFHkaaOuaSafflNo0HwZMhueJ47QGMuvV21dYIFXADT8K1/sq9HrGQPazFABgXYPijRkkEE
hsl2frsKNFpLcreU+zb0PH67PWtx4ibp0PySMTZ6kJv/YiZqSfM7Fm90Nub9+dKqVTmmrHfYlLHO
HMmEdcEZjU+/Q7O6fcws7qLK13z6pQFJZiWcZiMBpwHTezb7T59qbWA89P45UX+KGfN+YlDyoMul
3oIxwTe+xtXCDEdlYO57diS9xVyEDP92HuiOIWHt9Q80hee2Fo9votOfYGn/s/zuqTz6ho/Q257m
DBruzcngiWjyYwz430qC8RonGjakyXbdGcmkiZtsGN0WIx4GMVLauQeXql3TBeG0GukKC67XGZ5V
Lyhed/3yo4Y5jXbToIGmfaT/ZDGMsuIxlTbEpIzuZ8kYPprrrJCd0i/6cp7TX67uKIOHb4+BpT4I
/dVnpRgN8+LAjo8tBpzi0dmdCSwqGhuVvv5aaaOiFMzg0nEr9pxSup+LqDOQHizQ2KZgaSY/FNHn
s+tbYdhr8pCea+PhW3ZYQsMcaiuZa/jMG+B6IGqCUPPGSOi/IUoHiF41HSHs6nF5M/SrXzQcgIiC
/qSMo+nkC712Fx9rqE5UFh4RXAcJcHAFeAlkQjKYp+W9NGo8PDr8evn0wb//EMldqMZ4HtPiGlcF
5Mvz7qUs3hCf8pXbTk9JcqGXMqudy5xorgl9yRW+6vmN2TJiD6BcY8bHifvenKhTFUQaBOixflsm
lGeNoUOVVux0E9Qyrp1zGM1QFY/0aHvAIN7TU8LNTJ3NFx49FD+akJY4UKHtiGihgdQWS59RfJXk
uFIOpAjlgMU/yyA3AklJn/M9iM3urnyf+GYZehswlMzscQFmnQVmHmDnu0ira6dafIVlK1EkorEW
mBH9NS/pS4USH179d+kltlNQaPunLOOy0fgyz3GPpvivwj4yS+25jW9LHXmR8RnP45eZcBka1bwm
jxXCR7x8YL6lGbVN1vplCg8NzBrQEYOfUdcule0d3StRjsQkgM+Y1lAh8UHmDGe78Il/QI00nf1P
VUDGONoSykXtpId6trIkEllQXUVdxPzDC/F5iUBRGRor03xuXfuyTvCihrNcEzAyEf2QEA2hOFT2
h9UDEbgzSZCtaExGYgoRzGoX4M0fdPEF8VUZja5FR5ztVoBQ9vbu1NDX6vDfhkKHGbaQqM0BXMO5
1WIr983Hv2847bHNCyb69Nilaa8ASbldk/oUX4aMZOeVIEjed/nSm2EcNxIkt+aRyCyrqocpL6JV
U/dOtTQZXM2Pw8ZHBcIVY86aGR45BcSrBxJ0c9qbMis/bK5EWqaQvPx9u6Ka+AFucHofem2jG8AJ
qXKtg8kKAuCvN4H1vZquEltFFm/v5zqW7wcjjQt0yTwcjcNYuCezok40v7BFVqykThO14HsL8+CE
ZN3rehKRG0x7d5369IBeN9GQ8zvBjWezK4D+GAh38P6nYUeh/fnmrdCFGA5WYWEY5UwfuOagg1Bv
PaO41KO1d5sLoW2rr//6a0hdj4xpF2mAIQTUb97S6A3ZM9KdN8pD4oIoWAhANF16qwiPYYGC7M4Q
Wzvh7jQ1fSzT/2kqQtGIU92OgMPV6nggUdNExaoiRnzsOokMNHz+1OLr/mAtyUIYWqmczcZ5ZeeH
jxE5J2ehVEvaAOi2T1mEuifKo4OVUs3eYriyWtsyNfGoFNGQHCAWy0ZxVmf7+pZQ7mb8XotfOOP+
B75X3ROOjFT+a40oJpwgeV7YHg9rWJsmoSEQMUhST6mLek+bX2sluRcmvY73S8HD6mVFXQBtCGeF
TZ6r/ElSaQ3qMk0wQj0wVJ0Q076O1+0dk8QDaY36KbJr5ueb97oqcZlaWDO+rjIMKSj6TblkzPcb
DwC+Sv7agG5l3VNAwnaQsSzFwz+tjSb/ZZehtYA++bzYeZ1C5f4MU7Q9mDxrsLukhHrmh34HLuLr
3A1AJwBa2dnQAYWgI29m+TJo1sU73i9pCHHn6gi1DaI4uxFR9EhzVbVKrPBUTQv44qlSKoHuUurX
tur6cXHw3y3KeCxzV425ZAcOoJdb46PEoaPP9a3jq8kpZh12rrZeoewUfcow/QTsnureEC396vWw
wJgZUjuvWs77+p4RSSLKy/0DAog9WqpR7j2Xgg4+zI3mrt76OpgFOflH0QAlXBmjLMp7Uju6SGHW
ITqQVVqIi2caXQKHPJaJ0DS5H2XEGLmBBjHIEkBtBz9i5vlX23FvubrMZ4KqZrMqWomVVqXaGovx
47KAuG0lyf0D13E5M0eKGdWvv3vLNWSCFw6jj+MqX752zsko2dJTIJEUZD+M80pMAdU/WzS7295L
QnJKO/KAjhS0fpnwFwY5sTmS1fIfUI3cOFBTm6kvBqktBREv4ozF4MtlUhfA92r+7k4G2rNBLhiJ
s3UnUEbUUMBsaZt9sR4ea7mCJrZJaj3UF/57nJFcvcpAMUUykluF4JLKE5q/Ig8rVW02k31b9cby
fFw/gukgO9Tl0PtI5M4Eak2u17pYmd/JE3MwkFbBajmkJ/l8gnB9zfOgVzGKyZDVMydI/5lPHHTF
3LIU9P4piJcnaES1xpTR4mskKKdKskh3XpyMTlGWUQtb7MeevvVpnG6saM8JpqN7trAJDjiixp42
M+qh3xBmriK7CRob+5SydnEQlU6zX9NIWyLkwX0oDcJ3xELKzL9DZe/8C+O27BytW8teVdKRJZEh
7eBA4igkMPs9DLZdGpgdOSeWyUrK8HGKYTpqvaibWAJg01+hQTuZucXGFZmZLRqDaoYe7fH99u65
d8RELSz4KSYJ4o5TmfRBOco9y3Mjyp5bzRnWgddip+t21MRKkHiPv1jD9wql208YgbsLDqyTFZfU
JPF5O2CvBZ/R9kfNj2OwTgrvADW7JCcqLI3er/QwaXeWDkSrqMUZXSEzGVD4M48lvvTI/IJcUKMK
BAlqW7wciyZS13tnpFnLde8a/KgvFKB7QidnA9Idyh2vjQHKJxCEB8J7bHvn3YrFB0qWM0y432Zq
PWO8QLwmVqLV8+eAlMTvgz2Z87E2aaIM3j6UZGAR9r5v2oe3G/fv0wU9Q67cRjrYBJQNBxj86/n6
B5wfq0YTNW64333pHGntaj7NrDDloA5iFmTCfYLnoaq7DHPBQQ2qq/+uwCr1cUhMK1a3pZUSiQC8
GH2RTfazXyf1rr3bw3d6VCC6ERP2k0fkA0j2BTxCHI2YfGNIt3YuZ4b07lxq1hXLhBVQ9BXl+nk0
AoxDqGBrMZNjqQ9pqx+s4k253+yKGJnOMkIlq4OwoIdGbFdHrvk5CSEod81iHizlPjCFq8skz4au
uK0vQCVcSFh6mfszDrV8kZtsvg3/pkf8kL7p3pUx//xmTN0rZz4cAX8uqOXqj4TaRU4cy+W7tZS7
CJgL6tfMDBhii/qYOM075PkTgVck7tu9GXmP4SJSvqhprp4MevALeTCvn4La7fLMw69553ibquDw
4xAISFISWq+LTLn35HCbraYn8VVy2sUkR6hCB+zpXZ/rM+yQ/nDfhrWI1ht/hSHlmikoY+aaheLD
63E9ExxlEwXJov7AHHNSkGCHNrsa+r5l8Jb4UfPiyBKMtiu2RlXCuaCHiS7A4eUlkc3xjTMPacek
mYQrLq5Su7YPGObcZlitHDTadAHztYzJCT5kuuyK11M0GKhDQC9D5iOrvtxRPaKpGvocfAfdLs+A
OJNOBjYZY7IFgV/+gBi6KNunIU8WeJ0BVScKeQFi4r/V0o9OzM9ftyHOPa7a5N0mV4saAbsCTbpN
299bMRtDohd3cCyWDBhshTT2dfmLf/CVIc4BmclxDf2GsA4OaYalgTWlkHijvpRFDzG908bWBpXA
E3I9Yz5wkFt6vdlx9rVD4daEZM0XHKXaY59uP3S6iroUAQG/nKR2VWPgMwmXpaFzA4u7a6FpVNpG
Nvv+cU8f1cZCd9SuKlqIopJsqBu//n4u7ilHsW7bdG4ZlH5Lbcqx1h9ib0dgMjULTwJ0VV5cPnkZ
4WJeWiD4UGTPj0yL5gHQRkX7YHCrlH19SllEQo9OXlkbLPO1GHl7l2hpuAQndu4Qe3y4T+P5GzSP
+s4fkFVWGifGBOaH/uIJlBJ0s1J9Qgh/51GJXodGJAR3CCnv0Amj4DbgSSnQtIzKvUpRS4pSE0EV
sIvJtkQvx7V7pHrBq9o/LqmZuXb84AbePR84PAUkYV+X+CIACqAIGgKI5iJKsaG6BJ9uMe95gVMU
eJH3EpZ3Oq6DsyFX0/PsPAl3e9yWT1YGq0FoHZ6slDJUk+lviHm8gPzUFOPvLgrdw1nXWGTTlNxT
L7Upki0/flO2b76OWz169+P2EJxfy3miEbeEC/1Nbpx+kFBKuJgAryr9/e1Cgk1Qvl0JmCMKTCJF
ILL/+0hG52COD/7iIlYad4y0/INzTHKZ4S3zZ3awvcP12BMYHQMDS1n+XkNRWKXyxoSxc/Zt1+Mu
0X5EGEYEIMXzD6sR3+Tpihfw4x25adLLO959S0GoUZJTQRUYBitCzigTuxXGJW+1xHqx2Pw870VV
8polNTtBIUjXLyakgOJvv1iAxHuIWiNv8f27MyFoMM8xf8WusF8qe5eIDvnRsbPx2yQU4eknMU4q
6zV5gKKCu7MoRM7iwLEMKpKmdZ7l+FMNSIpEpjhW1nez8+5yboDj/Pl5N50LYuHNbAtfpLm9MZj2
JyrqlYc/qQPLGY/dMXmcaq1bJyiaxYr5KBEMEO9aqJr6vJa4hEW5zU4M2r4rEz+TcVfGEBqR/MD2
UxKLfWgAGz0p41C3cxaNxjwEhLQyEmtcQ5roW4hqBPvy8TiglGOJNh0gDeSeTgJfMjXhvMtPp7EI
oaIfvqP/pbrE+bzd5iE61TpuTWfgpw+2Hj8DSxlKYsiGsMyMxAyzocCNF10kIn+QwaLXLKo0+YiZ
6pMXMbyil1XUGaiT5MWlfMuwcK4TlBhPwb/LAbLnwQ/lQsd89UHwnMZEmPNTONC0rAV10DKN87e+
A30CwfqEIPM+sZ1IhsFbLW5nz7x5Ym23h+iBLmnNnOYQ6nO7SIAieosq1o+xHNUnOrKcXLaZLT7y
C0O20gWBrFZvWcoa/3wzX5FFwm9A3VnXTKRGXJUnzhQDRNMB1lX/oEqTZzWg6nS6zEF8q+O9KG0v
wiH7HLbT9uSUAZnHAkDoPbKBdnHJLa5dK7N3UPKjNReQUDnZh3d7bMgsowmQ1kTu1XO/CmZNwaLv
nrspFVuZsJ/2cLCl6N0VTxeKHKD2Th/5Fz0WTuLc68sT43hcRZI7xr2AUFwzgK+M8y3jM89NGkXQ
ZnlxYKQmadw7dTqRkOqAXSjxoK3Tlxjc5K/tyzYLsCjCZr7oi236KITe99vVsur3qv5AaEDhoK01
qwYVn+MnVZxxFap0zafttPDpIURfN1ujbk6J0/tW6HojEpmnaJeQPGMM5j/4I6IZPO9AjNl1Jjt2
uXOU34lBdfM2eXswrN56ldZ4GCs1aajTbs75SDz/6sBRHt3NPkkCzxkE2i48bnJx5hSXVJw+/Gcd
FWjJx8LUfpaLqyIrSibpAmKDiOODTVCHIiLjQwqPZdDGrrAYjbVKLr6/s+81fZv7ZQ22CHYVMts/
5G7dEBDxOUGQSLk/fmaQldUp8z9yR66438iNBLNk4zP04SJZuuvmSVRGpaHSE90muQ9dkWYegJjy
cVIp9g7uPCnSrP+0uMW9kCXZh1WQLPfSWBfW4cHJiy//XcPVQBY6cmtDlNmAQJKJdr9StU4D4O6H
p+TCp7HskfN8H8XFOf6wXOOf1CqRuBLoBfi13bX36CN/OzTKnsGqDj/1+rlOVWw6k1TcoNWDq844
2LZwZeJTG87Zq7hRfgTUNXFrWMu+WLQ47lrHZ2oxHUFqSE9KlFXWEO64JrV/TtzdgnavsHWD/ETB
Hju5KQSAglGPikxg1goC43lEJcBgcr8ArcE+iJXZySZdA/e27Sb9l7IEaSLPgVilUfkk4ogv9NQ+
wu2SlWkc86CTbC4RoBde+nYUw20rs3ObhIyATNQO3fFjMGn27ZLEb7qw9O9p6XPJhgS97vCL0kV7
fbJksFQ4hjjYxZ93lYD+LIztlsIxja4HrVM1BlVOC21+NrrlLRASNcG9TuCi06PSBHJtyydKmBvB
ioGx+xycTbjOMcgdIX3RyVKsvU10BqwEXvlwKobd5viOvpDifA8JlVlKbMs3T86uf1qgyIz3PgbH
pP7D/BgrQaqZ9qVYWc73p11K05ECWXbAzi0GWgDadgxjekhpJAANnxi/WT3wqcUF2PLU9jfh9oTg
6m+ppgvQQhDiKKVp1/FvALttCCea5SvoKD0hZ3FmLX7Npta8ne7PrJPm32h9sMx6gQx/HLphw21g
PXbxIleurCMIdmRz9kUh++KYi/twdWpFG5MLS83nTRTjza8VIZzJfn4rzwtlBbTGMaTNpzV/7X/I
K1Ojj+6SarFfbkPoA5f/LH8LMwXZbIYiHK/SRT0i8nx7/W9QgxFusjUKwbeIaJ2ytkjyGN/OPNJF
/+izgEjjCrmEMYiYRTID7GbbzU3XCnXKYzJzvE/udSFpcSXMCK/J9+rQ8F80tJakEV7b335tXV4a
MSgymwVlxHCuAzq4A4jMNJmaEknLdZ6dJJJc2YZLSMNdhgWuug/7kUgUOjxPzlyFkWTSCFlv2OSp
QfCBw5dWPOcNBBE1rfIEoihbxsjKF99kqEL60FOvsRVBrnxLMFnVwvMcAGvqJ/+01wFixjkKT3PT
y/A1WMgeBk76Vq/lXtlZVutGINWQkTUg4OjN3RMm54aIWMEY20e87dYCSo6EKC3awwH9KkevsTQO
yNtbN6kUAJOMwbWk9OVmj1tQyYpDpKjieOLmfyZx0yxSF+yfrh/4YRsEa63W/gevDE363GHG80k+
LN3FOYWufjho65+4kuVHIh42fbcH1DgKE7WS9+tUJunmVWNOb/Qsvbrhv0+gyCAUnqiqXgFa13W5
sQmSBodUbntRmpvu3hPV0XSwHAmzCKifY5SUl1uDmE/WRuspCbyk1T0Shu1sFbG6QsOxzzdADYNa
aSmnwGt0Lw6/rFhEiAtSe5iJoeTXbZmJstN6vgY95qQ+XepTyYK7n0II5GPtfOG09u/qenQWj7Oc
Gvk7+S04u4E80YDCDd1GyvPY9Eifd8mICSi54TiSV+sscWsbgxKPF7tAttgEJdSoUILzdTiJx89j
CPJ8dwmAHH2XVcxiebOeWQ/1ZjGtWDoTSxPgKgXaWt1nxd4e2UJbHMHWi7t7Cu7CcdUHKJ6Z+A+k
g1cRqKAwKfUjF4aCTcYLll3q2awzS4H4wxWaEMKLFgkmGJq7FotcuoUvoilMKtjv3r2TlqcaJ3qx
JD2Q5vBSjQ9YHaxXyaHAj6H6mc1CY9ziHSLqOWh2mJ3FjR9XvzXFjC4tyBfVofy+1FOeUAQNB3hN
v8qsfHED3m+ArnF3W55hlLuDKMxcTFJO9mszUwH8d8R9wJtmb+hbttYFMbc9GjJj9OMWME3PBICW
mEgqZXlaIXEq0mjN77bxdfN1ySxkwWGBG8T/qWU+Jp69/1coRMhzwapSMPoMHrJ7D1VZsPm+CCKe
KyRo9auWBXeGdxppFfT3vf5mt2lSYjIBqRh6MRezvQsvWOE/7ADK8/xRkk4yLlo+WqZJ1MPl+NtT
aHEZmz7M+3YrBjd1ATGqpoBf5W5Y0oWPskRBASdKpT5LAjfp1IiElLzXHrFrRYrfzvwPSXksaqWy
1RfjabiKXb6FVdgqhY5ZruH/8aOnfKPHf2/uPwCe7CthXCEFNRz0vvZZ5C+yyhIjBz0cX6EcLobd
JsZ81JaM6P5b0n6WYClHZVIUeUATiW/ZH3cV1PsTTzrqTjPwcEx2+9I8+X6KgU166WjZpvn+ufiV
grgM1Op9/0ihJM9A9vGpPVeF1AnrGo9K948r3O6gUSOB1hQdaTPC3EyE9BhpbjnMNzSPcmrsRz7l
dM/0o67MzL6gnjnM/Sfoz3dJUtoHCu4u7BNiKzXU0gRy+OZdEAR0vr90k6Xw9o/fdth3NCF8VZFs
w1LsoXJlpFVWojToLuU3Y3s2zu3hacsTsPhMEMtafel23SUNLTgC3wl+rgmlUnYFiIPMUO9VjqhJ
5YKtfJQmvVi1jMUzMCRTMS4FeXgDkamyc7o3zgplX/Lx7KJy9yY3KzYGUjFmjANx22LKV5QNPV7r
GiyjeV7bEzPN/0//feOTMjeB66usixeVHm+8nqmxZBoM42kb2LMQs39AMhR4a5J6CTuDFwpLbhCB
lqoYN/XEpjnbL5G2yy5jscCYr3xkAes+MnMrDqIIOaX5447ZPAmOEe9b+C5JzrXPhwmNYSJgINf7
/jRzgU+Gp8V0tyIPW2oMtqKp4xyihnucLvqfKiDni+qus5O0kmq7JOulXqtOoI6ApQkPuxsvNwBZ
zfqa6iYOvV3sezS5bkljLWa/0X8uv6psi6QizeS9P3zP2+K7EAGw9a/ViHT4L37YrsaPeE++rCcw
m7ZtR0ogFYqBfiSewYgB2HD+/nFffLbEqfJOi8AEVttXRS7t5/OALgDlhXUXB50NF1c5ubpr0zMn
wz5jJ7jkmLZtIBfZdTi1HVXKIX0voU4+PiBk+blc/BbpSaxqrrglkxBQACoiIBG/nMIPn9IPMER0
cSHQIUqaCyG13OoV7WbW4McA9OBAGw+s/ef89lxkEFZOlPJLvxI6kLZGa34Rt+NQyP7dM5NpE2Jx
n5Cw/T91knIX+z6bxrKnYPMjoGjkECwyNQtJgN/x7EPhYwj+F1jVuaYBv++zMzrRK74c+AqxOqsL
0+YsuD3D+YnA/y1DVhGz5kg8i2ktSrbrU0DDutjqK44742fcvWvERtnPnQLnxSuBSFdc7K2SpcoE
5/S2MsV7tSUHGayqi1nVuAQbXPlOwB7cbAIeDEoWMYZ8ujCE1rh5hmvjmdJzB+AzcKoSKFjI0vWM
iVwLmc+oqRsg9cwxvcZIakl6/VGZ64c7hGHrxmb8l6LBTdU8tz8g/NcEo36/KUBe+ez7kw/VPsNg
RMz5nxzm8pIc/AseOI6sr+T/ioebS+qJu51kuuCZdxK9TUs6S4xEtE2l1vmxzDEgPxdgizBPCE+F
r1VSDlVH4zzmhfIAC/59UES4G/bbAavZgae+BIY5I75cWBC5wBHcAnes+RxuolOqeSNsCDSokOLA
rDc2wDVVC2GlOyip9mHYWydrlp7AsstuZ0mUeul2ovXsJ1fItRm5atEK6HZhel9X6wTYGtWcjWps
R9DykyiBzVzdyHkY+W47PcHe+dTKx2GQW8wufAOYKPks82pQ6nXXYv+/MLcnXUzyarl8j04Z2L4h
RToJAKm/pahM6LVcj9kVAhFgv0nUtRbNtCGFEPiSmnxCOaGLQL5tVLnn2mUvP+l5J0zZZ1Xp8+3o
27q50fyphBuaUUtiwDOtxk0Yqrn5lgLwZScWKmDJq0nWdWlQ8bSSPbndiBPKDVW+q2MnNguBuyac
zRL7AfhNLVkzqdXFJndAz2y/VIPKPUCCv+Fy7t8pgdy6zhcX1tiYr64uXP16dlSUeE0Cn5o5h4aM
aC9GjKMJIhxfJb8bDdcXPr9Cx07POJzn/vWHIU0cEDiO3k+F4wLqQOCmZCqVS4aaYk6q3VOdqS2A
+VImCRpprJ+dwksbvZ8XK97Lihl2UyHWo/8SOpdCZPpz1alKQMtoZiORJD4VSJw9uxs1lDXbkGuw
qRHEtmvUahor2JAhNa3mMnBKJqwODEU/Gwx7bEto7TXhSrtgSX1xYTuGtXMRH4vzXVI0irk9H85m
ZrGgxtx07htkxi7QYVkJm1wPXio6JlF/V5gea9qcsi4CS7TtMoqxYM6Tpo7Iz44EEebWtoCOVxPV
qwSIjgtLyYawPuBcJg25jbdrZYec6VorfukdYXACLKhSiKddJUZpUiaXH3Y6Fa2RrhYV6tsiwBAa
3slLUOoQBC9Z8JLBWDJgRg0xxL1fourZ+sjSoHtQILKI8xoD6VKsSgVadI1c9UK/csMVHjR0Pn+a
SSEktjNv5l201pgXN1irDvlBRGSW0ViZJtDquYUSgLa8EZpL/FhIn8bbotQwvKq9jbAEbSF3MkEd
CScZVRnjgLhmn+NFCcMNusV1XSo/Nux37jxp/cTPvxZZ5jAQTzytxj/6z3fHGrlHuVQIBn7uHUA4
+gM86r2Oa91DQalybMCYk6cZIeowKYDUoX/Z9m0pftZc5+MMckxpPHMtzPAEeR21tVde1J0WVkkj
WYraWvKTNEMf/j5I/sUUUFLpWGPL7L9DwNluSh1Tv9Wo/QXSQRR27PtJgRLzfGvRoTFHbiLzV+SD
CcN41uR88xSG06gkDvk8LSjyNBcVqA9ka42sDiUl/vpY2zl5qmMes8aFhua+vd/HH/QtgpZ5zAYP
+7PMoh7VepU0DEA5j4dq91nOD6DIdf5loix1Ok/yZCnSLyd18l68tQpQaAA2HN8hJas6hU3Nl0BR
WIkrhLJBEKtiFnIeEJ0SeuKD9XlKosV4kmr2Ki29hZN0d93lQvKENLdXUbKP8edpixKCpFKn646A
E2+vBjNqRXZP2WA6xr7fxzRpfYdb7QF3IQg680UnmgJSHOCiGcl0XaDFNV+B/2Zp+/LGAGdBXQaB
8fzkhSWAKbBemkvjtMUQx3+ypgtq1Dw1TqvXt1ZSdFVMiYtKjP2OjUEK1S3flJjC/FWg+VXxF+Yx
5FKCDE+AKFkqT78evrQ9RBa+J5mHY48nycgmbPfJX9EjhFZhVuJs+YVrn1Wq3CWutMUIgprKP7vb
caIrEzKpDUbsWahFiCPGH7WAfY24vCFEGYu5bAgAbR9O4GLu7GBLXGSbxZLdd/kqsMS13sv4ygzl
+me5683pqaYIti0NcuVrn8XcYO/anVs4xCtvNdShKktrbBpD4S2XDQmijqdWZXsw+pjpIwro/SkY
4f0fThJUfUaP77nK4Plg6SJeW6JyDFHOLbwyltC4hQnnhGUn+og6gA/O7w+JkOTF5Y8kPDll5MXq
+0+9KTigVkYCyeGfL0r/uJ3XeYWL5MGihb1BfJnOjMDuk5ANYwFl6Zi8PAkEpN6rzbKXu+0oT5uN
h0+WVaWJHQJZPTCxiHL2cCUwjGnJI4QfFfPkyqTKq8Okoh/yKwYv0zaZQL1jTe/njRhcy8AozsgY
kEsDY3JRBtRpsxk7wtdcJrX1uw12eghZm9pvCslvnPf9UFF3kpPnBQGarM0TyQmXZ20G4Y+eFR02
mQovU4f2wxe4Ul+jft8qA2Itfnt+eG7ywbMutBICsEor2iDUh7uj48NPh+31XOB9CejRfJlPhate
yUWQrlb0uiU05jXWZeW8ePrmikLDUIL1twUIHlJYMocwOGJNwwcKe0NEpNzO0rrAx7QgL5SylS0n
ZxAFkWFJJZ2OroAlHhTQqMtAEwIhk+jFOGPUkeSFEV4ELKyFtp5IzZnFsfqm8Koi5DE4J0WylfNO
Z/BuxxJf6lYRfUcooHDMTppzIO2a/s728cRaoOci7s0/hHsKiMoAXJZar2NsYZRyF8ug+ZZJnK4L
CF/2AJQ5XdbH5EOvrODw4QvfoKsjwWfP9ny82j3Qe5J9o6/c6Bxp2GWrvrulVrEI2QcUWMkLJFc2
NR2NUR9Hxbpe98Wpa9plLk4RjcYXKxCqKoW7d3qK76GPYTCiXV/ASbykwYdKZ0uISOm4KNbb45AV
qBXjFUiSNJPEoJnEHG43FeHX3AKqVmD8b31LuV20zqkLAGN59V4bX6YLQcK+TCtyR0sK8XUQ9+I5
IzAriu7sZCCdaks68HL5aABrlPR4Wwf1+7aEuiZbJ0E9xBo9cjMDqT79cJH/WMH5c4H886ufyQzl
mLT4Rer+j5WMF8I4ieVvpAdKtRhklF+QNr/If82yUqhmE/XJXPK8fkR86Bu4Gcp09whFE7r2cTPX
rwN2rL1sNdZqhrP1urh9CGRqX9f2U3QPofqRCvcfOUIzhHtWsuEg2xbefSYVDXhJO46uPMqNJqvI
qvgJJC2KPM0vI0PG8rW46eJ4ZqIgE5CyCGSWEJtdqG4XCgUeMoWcJp5oMGnmtBAJ2rPyyr2xzn9E
C+9MdJdZz0fvMidHF2KpD7ImdtlU/IgbuNfa2JWVhNZEWGMkXjdyujmRDYaeh9hXes03eusshUJE
dsipPZB3gi2GKwMKlApvLKgtfb61Gx0whHK5GqaBDWXEhBtikqpftjuf/q1gaSGxklhOqTxdCsMs
g/2iz9bsOThbw+tmEPUR6S4wUcHxsKHcJv0aZIsekV88quYs5i3AhtOqHc60H/8f6z0RpmKo8TqH
RM9spZGqGfEAZIITJ3S385QRCRdbyh2L3DdXV3LM+FuE2xY6G5cGQ6Iv+cmNLohDLW/Uj1Ir7sae
9loMp1gv7/PO2yq9OHJqOQJVoRVorIUdkDaLbiDDPrOhUNLR+PBcPAlrdjCgAD5txYisz/z0H112
owChTiPHsOfM9xaUDNArFO7McZtt9nyRFra/QMdRjufdX6EumwEz/GanrlVJ7jg3g9Dwipvc67Js
s858epLZ44SDMff3J0Nzu/nJTmmHsURP8v92DHG5hW2mgVEbDPt/yyDfVoAXXbnx64zFo8ZbW3F9
9Te3aQJ3i3k+EkqnLavrfHYVaCfJeu3O3DK9owULv7b3k4LsQPpIbinh3lES7r+ffPv1WUjJFQs9
axtkbreKK/6aKkqh37UbRVs2zBcdTxAkm8AqS5Td/JAX2UDytR+Z4pdIlUllFCRXtJc3jqd04Edd
5pWCbiZW7TmisLgdUpUcmApLufV8CSishCGLOCCbwQMBaYIrekPbTpWKwSSRtu+zB1KNW+4tElA6
8WU6fZJ9HbtG2Y44ZHQ1H+FVrr9948BCJ7MBB6bZw33gpqaewRdprASVs4bBJEKsaJGfxCtH2V47
W4ckXuVLbEaLMj8DFXslMp37dPZzQPUcqmFU7u5ZLvT6pQKcWtuCmmtLsXgLcdxLwJCD5hL8W+P/
jmMS8HuXlJ4s+4z4JwAfIGF5LBGDHi0YAaAbtJFsndxDAUIYr51bgI/ADPpMtkTUpEIBOdZakUEU
xTJwckjPTH7c6DSUBSbcEuHQIBXn8WYDsKemt5SDqaMW3NtMuqYM7cpCUALBXaOq++XxJpCMdwys
Viyq+KtmzgW5n4TwyphwnUsLcusGitVwckp2ffmB98GGZ9Q6DBZVhdb/5idkcZCftWXAXw05k6+u
NQgj5qrOfCVgZX/xP4Asj+SBKBjS9sIE47rzSU3McKGW1ReI8iFh+dT2/ysZpJc9lIIatdoe5VV7
dXwjbXp4DuCmkGP5jUCfUbnxQscINYc0c8nIHEUWislPuwrVe/wptJAf4egXUULpnlcIPig5BxjX
pOUWZ3f8nQAY1PRNOgD0JVjBnVIXZkkfoez43biiWxvQv9OmKGnOBKLlEegpwzzKOBQLUYBgaIi8
E8UiG8oPvRAgR4mcMbw9icrLgmRRh+YGaBHjyaul4hHx5oMWHktpxmlLCNhjWBh5BVUIHcCkoVAl
1Q2iwhn1eCPrnLroeV/CnsOCLyKNsDwBFRGFfopAeV03DgSNYXsFIlMzd80CljFgVZsVcR2yw9Y4
PsTdIARvh7H6KjS4pxNp8nlmrcEIOH/Rl66HPiuSoVK0RPnuW3qz+th9tlQCKlIJ/26wZtWR5rWh
mG4RJd/tDwJ8i23FnuCDdloUvY7/STi1GeD1B6IY1FdeQ7VYwOIo1MEAM5Wbu+dKj5XUqdCXS88K
ZEnv/vwVMgbW6FHBabkCb/8OpfXUnp4tJGm0AFkBjOxJdkea5KksqpGzFtjZQF6icpG7LcpuE6RW
7humHBnhs2y72Fl2QRK/S4dNofFRkqxtU5Szz/teuCXcE52l5Ms24Q7aCb4gZr8L8Tohy75NWnY6
2u2wkjVMJOYuVOJCHnVKL9DPhGExxsHDnbIRtnb8EIE6UYXa8ESldD2EGGNKGyiiVPDg9JtLMLO1
z2/Gu6dP51oH9T5Q/3o/t+q4zX+mRkqptnApG2dCe6WXcORSNatnVGh0dvIIZvzLT9JVavT/1xnA
S5oL4EJG8/e0ojo0+OwWrIgKecWKvo0jMBKZVGDSbI04dDk69vsO7qE0RaawEim+hi4kUy15+qSi
wlvZ+oEgtdlsApIQGadIhT6IuFB+IE7vmE7gubgASgyYlQazHu0kR4EoaCwKnq5WJRvkiunWztQ5
tEA60DjBxNwe0do7Wd4k8huxrAVz8b3l6aQpJVzVFrExdj+FKIU3LoKRUoEDLlMRukiU8cydpjCr
H2609aI1oH4ZMRwwD8dkmZzlmKiKitnuRb5wZTpe84MhaHG+wodCBemOveoF8VWvcg0ad9cfWSxN
gmLsPnrlQXoynlpJQfk5IoW5SYjR5zlHdwmPcwD7v5a1YKiu2BSZ6k4AVAmnhufWCEDJdi8NjYAd
kVrNKFZ89H+sdewjNx1kGYsxKvCagiZ3/R75l9NGfEcjx0/rmIRJaiQN0nGEBtEyCa7bj+echZTl
by1MdeX2pNnyUCy0f7iTApH/DXG2Lwu3haB53+/6SHzKCRFI4Qm9rrJRu8u4YaXON8QpQ12lM+pZ
ABJQcEVVWe1yaglJO3/TARAjKK7y9qfDKxlKUuCsoK5tKiW0tRPGKU4x0Tk2ehlaTs+KmbwgWQRK
NUuAgFQeZRHxnTB4Mtyx8+9iJDgJTlc0ySMWorZ6XUp8PAekyxbp8qZeKH2Y1WqxvSUQ0JFFzwWk
c942CiONL9dWmvxQI45FBQiLCcUXClFpXwCJGHnAhPkYgGX4CsusQEjzO7auJkTBfRVua6ob8jk2
LaaaVy/U6dUOXC6wiFx+Iepr8cRiZqA9Iwf7ZgYRY+xH4JJGfKXsWzs3KZp2hOrt5/fBNXqrlrzb
cMRNTOanDev2EyYLqHwhcTMirqObeq6QD4kwsmyM+J9g42mkAWEbaU4CUttmnnWqa5zK7yDXJUtI
Lx+IFJEBrAaLwjN6rU53w8IHeW4In40pPKzM56d53yxL9jPNmKpOzaMIwDln3XUkAaz0ZddqkY9E
B+srh8SCG/cBxVEoprrL6GBGTwVltqNfvRrkKLSuhuV6B6Hrt7+Yu2nIDZX6NUUmz8QHpLEtVHla
Alsa/+PYrGxiyfrFKNo82fG+UCQ8DsJWjhE07MBz4oxGo2nOf3tzp8D6iDAn1nrQaAWOgN/1hCFZ
bXWIoXqCnhrG7BSvyUaKYVBWQPTIdlNTvgTkQFtSDgGDXnOBtX34fDOB7NszcPdtegxoe4vc4bdK
Fsis0q27A11St55Im69zp0k1PkCIGvvt4YbEg2KkKffx8PetF1PdGbODuJM0vZKOMVD8qfqL3M6E
/ke+X1uzGSS7pvopH/yUqpxYcEVFhbMT5tROTLg5u4/KUiLlDKL8lBOLJQDhHaExDxBckSmvJSgh
kXFSytAmb3YJhwBl8QPQPVdqmhXvB2qhqk5bmHwxgDHF+VPgNYvRjJhuT3zbXZJJp3ne4CnQnwjz
+hznKCNAFz8O6WY/TDtYo+lFi0CtC/Brfi82VqAMwnzRmztN4IIVlM1te1emlv5LOADaVtTplZUb
vwG22clj1A426KE/S08EfbIxxVkSu1ItfuGsbsr5YOeItjH1SCKvu/2VdZZ6wOI28H2iO5+ahs5m
GMVSkT+4qwsls8+dNCJR9ujV3DuUkge+lwqkiQSpkSBXMHsY/OUscVCxCOYoigZyWO/kz0kLI5fj
+qy1K0KcefV03wkbCFQ/3PMBj95Zyzqsq+4V7Ss3vG8uv/ckuTA+b1XXcwAAHmOGMvJDD3O4LBkK
04+VDh+foYl1Bu+x8uaK6MYdvscVMNpWDQZNMH7dE6ShrWcmPT40QiQ+9OKKvQLj+114td1r4Pg9
Oko+ih6jsOg1OKT8/scsY5QxmCJ4lMSgrvLMm1J0muzmThQc8sWe+R8Tax24X3APw4SSj5eR75dI
12l/v8Zgmq6JgRaJyxqHrqH675lqsWFtYsMo2h+l8lbXjygmGRtT9g3+XlieG4Q5D6UICT5LxMbf
4nlULkoRKw3QNXWm9AgwXYGZdpFG7B12sT7ZpA5MS8kN2a1B9llnChCuDbQjdWMYBn/6KTangSUM
c0n26dx9ElzP8337OzXeBlzaHen5pmIIn0qe/53nYeBTtlBO1o5mqOGkWfyuUdKqxDy+k8BQxPr0
Rozh4cykGUiBiEV1LjGaBN0f3gBOX8tnMzn/QcOAnx5Bz4NO6L8ZUiY9PS7CAJJbmWXAwtpsn3Kv
/Od19Vs6NbL3CnVnpOyGDfVKESaJwbdHCug4AeKLZLDCeeDAFkWSHmADvZFYKpVjkhek3wUZiBdZ
6Bp3+fDruM6CeE1v4W/3UaBld4WvPv70eXa7Ry2gz1StiHwlwlF0+32r+Tfq7fUwjQ8ZP129AA9q
kX/SJ42LaL36/Q37qDyGZ2cCAvXoLLl/MvwGSbV5CnLzm7pnhEyvVReQfz93yVJGnwx8Nj/9Kg6y
7ANzcvTLoETQq0uj+oJOcp/mDqP0ZsoXi7DuQRtlo8pe0HJ0ROFpVvDsT/wjOunMkbUg/o8ui/P1
/GxSz3fADY1Rhupki43aXHWA0FBtAZ+EA5odhPJdElvmYiXqcxhc0UsoPbuxrD3+eBMP5Vv2QckA
RoNIt2648iKvemYXWlUBbph4vpAG3vR7FLEjrFYu0+Nud/vtmBZdm2VmehFDDvIlHhMhXMus/yIP
9QWbL/8xt8I1Nu0jGpu7fP3TCHsFSmJm/NVyolEaLrMgAoiVLGUpWomiXb38L0WZXcXPFMa7eSKf
GyIkbuMT17ERgkm9EGGf/Nrwfm//s0+lHKfNb7iHcC02xptNSuEdgWIGMjVUJudHkPX2FoAopUgg
v6SE/REQDkZIYjgUqTtOUAwZ8PN0fTOU46SAbJDxMlWeDziZ/0gUyU5FPaKCa6HkSOaXf+iDop2f
hEdWzwT41bppu9fh3aW8MIfRMDmg6j1zi6s5W3L5tRlzTldfMm+C7sbhVs1Iy8HeLRkf+Wp8CBX/
AmmGr8TLWdM2bHQwl6EALiquFc+mED0GFqSEoMZMeXTTNGkJAD9zaH1Os7XvKNpLZWC8i/bv3Fds
ZOHWbRAy9ntqKNpDmNu9vRmFGndcsPu3s5kXYCaoE+xBiWeiEeWm6hyCafo/W0hdT9mycipSJtRv
lr0qe3Z0Y+zGwv9958YCL0Dg1p7vhkYnyK5IXXEDoWclOYarbVfjJez3Fl7U/Ws3kx2j51ojfLlR
zTrr/sx+xA5xmfWgOKQ3ecGgddcT4Z4inWL4DifEY7OEcFyHHeHBIiszAbTH97uzSQ6mkm1OIfca
0FjSP6VuwXwFt1aF0YyL9c/t1cuZmfImtW0875mWgVBKizBJEvi2szG0jppXu/bUrO1D1TvmDGva
mguzjBHSfmxlk/zDmwb1ogBXUPMyA0AZGUGDRg3T2PN+UK+ZuElq6/wKyYleBhm+zcRzYFfbR7OT
jCNRmj/EWiTolvC9Hj1GlC9x7sWOj6KBJsxfyHxPGW4SOeNs4DFZVFw+CMOkXWvl9Dzxde8Dvu1m
oD1oEP7PHrKPFD9dHS+VUF7DzVaYWbBFo29QBM9x8OY6Yd+j8/P/y3Ygmf9rw89heVBrEj6p3p+E
NoF23DHZ2lr/aVWXR+GuUKio6XF+jSd7TgGpLuKL1ZOERlsO9v020aH1GztaDiBx76lwf3AysbTc
RDRFbmcN7EdTbrTTquExhLyKZVDzE+BaLTEWwL+t2UCRHP6tDV6MxQYVwGXzYugrLSGhcv/Sp69T
YzPIQWF9wLtZWNisUFEZBr3iyiJ31vkuZ331E+sO9a1Kn5pIFoJB4VbhyodoJcilRXn6qs9fF9lB
kZkITezGS+67BfA7mUtYcVz41pdn66a2vnSy0vbQDzaqZqNP1LOqQONqxTRbqdjQ4E5wxSb3da7j
mElAv0qVu6pHGW93O89JJfbKkBjtIqPhNb7uMew8b8vTuv0oHuTL8rQywnClYtpIxu84JYDuFS7e
rJR9X28puTY397BJIR+xh1ifSoVzYYE5TZkmJNwiMU7lySWEF7ApPN2gv1aX/aeHZaWZGA74Ijqv
zwsKJ7PkLIyhfUQC/XaYtBLnhWMrXxYTVkixlG/G0NACOBTABFXV5AY0VCJuMjId/RKZV3MLB7vo
076mFpZASjmoQRVQnJFxuVbynIJ2EyjN9IFL3xj3o96/w0T5OoNhvlFt/1pz8hbHfc8iTe5RiBP2
NF/D9E0W2mDr+N13PVcTuUd0LuiQixGofN0S2RIt6RfA0pBLTdQJxRNAAuFexMqboUo/0lqCdu8O
eKHuJBJyZaf2M8vzA4ozGLUaXYYGrm+Cj50jdHXQfUKA8TrTuP1e/UmlPTPstwuKPg1/KxowFiRG
JIDbjJgUpkmf2MLQm55eewQFX25gsyKgWPQ779GZnk8/10YI3IoNiizfntfGgiSdqQnYOx2EYmAH
OFsi/34GJlJTeTySAwIZEAAHU7mLKwAL0M1gZSl0UBeqCuN1aiZxcdgqh+i78YI7fR2zQWoxMRqN
3NyhxrLlBRyUwwqcqHe4QMbfBq2/Ag72UqURaxwtPUyNHT9GAb2MQ0f8kbZkrN9tqb7jDabgUYv7
C0epNkKlOMynYzJzXzBKO2/hPM/GBUyKfHiD29urFwWNbseN3iLrL4YDMhJJTS1JqGqpdReyyzQv
YOl3VFVxPmgwoKCd8LGuB55JE4HxPnYPK2OUapIW+nXrByY2TsYBYDgur3OaC+G8yAu7ma9jlMPr
cBCeW3QnDUGnkeDP/mw0XofQC14ew4ArVoSBwv4XOGMLpHC4dxF74he3JOVdq+kXOH96EH9GRtYD
SgwKttU3ISeI49FTysGa2toe/ut+XYN5mZPeybrB1drYbIacclI6ogG7S/CaRGbZ2lG8ItfyRu6h
30Y24eeJHY+P9KIc8oI29/bNv0PhZ5w5tY9i56ZcbxGmBafg7JAf2rgrhyuuXc+kHN0GB0rUJYFn
MCyroAYmXs9OxgpbonWHd5YGIn7YXHHfe9S23Gm3TLVjVyUQ9L/fgCAMDnHXLZejViU9nk36nNkt
FaOz7wqDM7z66BtzM+FY14s3lv5pCgTwF5FJCq5yE15tsFHawvPFW2qi484xGpIudYn1mI7rZBGs
MKtuvLSWUgfKEiUoqM9V96KghiSkaEV7b/00y9RihUfCQ3ZqmppS0LntiybKmvdoJANhdu5gtgD9
Fwr6Mjc5ZHiY8V8RGpNOTuHYZsLhL12obhLgzh3YOHV69UB9YA2qmZuEgGxY65E8G0Upa9NzExzw
teq1uav9tngu/aDDJeD4/Ax6u87RfKIkiir9QoTO7p+epNCRnL8bkfCCck4/ydu5IPp98usU+xNm
Ub30pZ7QyiKgqvX2FQxaMsDgBMaNSmfOsXErtGW+B5HOuFYYWzhUvihonjYpvMpU7NDyolAzrYTt
ZhjAo6dr7n9qhm+0DgZcKKYmiN3Id9f3mPNRBG7nEB+pyo7l/r6GdnWyd2SIkbyPr3pkaTpp0eEu
Td1QzKsr00/4vRwhGvoBiJ72Zi+Ezu7XxWXdQfR7n81/LJRM4QIdgqteTvYvG+QcAcVGu3SP6Iwb
TJXLbGu33HJ4pNwgAWdwRdIvMPh4kh2JMJqQUTcFY1tMNliCwQlWitE5p+YLGZTx0/5fcRFlR2vX
QXb2B8eGhMzY/KADDjz4PL8i9aAYb65EdhM+YRAS3WNtDSaz0sVCK0FVuFbb20ern5bnWvqWQkM+
R71tTuVYaIpbJy2OMpG3i5hAdLRQDixJGHVFjczVFMZk6ELr/JvRh3p+90WHBqyRT0ndOArU/2FZ
Lvz1E2Eb7doRuJb+vDHC4Pm+509jq1rhr7PuDparah1k8UKeYZGDNQGOUyfQT5hPuYY5sJQ7MpAW
ft+D5EbKdEhIO5DghJR2gghdQ9w1cOGE/DuVxxF3xhmtGn3li6yJw65btWbNcsCdKz0BXzUfAWgV
Cv34IcP7KJu+HL0cnjQns/EQHrxEaoJDL69mMLdviLkIZlKJ2AWRTotwm/uqSz/jPH5eGTKBmLbs
dZvhX702nCTdrrhvBzPYgFhj+jkkLvPuHpyLRf8GXwwUsduCP7qN/OtqGv4biYih8WQ8I/OT+l2E
28s4OQAaIhl/qCwF3WeceDAmxTygt00sGjueqm/feacaReEfFBP5CNTcSkBxfYvq98CjcZ4Fl2pV
j1e881puW4DZ1Yi/UKGu7cnHSkPgh7v7Dq/ucEE8RmO1DSsmytPmzPbSmIXCWzUPFbZInB+WONk2
6/AkEuLUR2nakKBOgFZzyGzrgo7CmxRWg2ow2Jlh2BDep1x7OQu+MuL5D3bkdgi7HfW2BgwOwWAI
cYLi8exRUwUQgQ1k5IAl3oiIZNkODFdWT2uC412RgRZqwLdI/ugNVV04t+roB27205K1Yj2jP2jJ
1w8it/4q8RwOEyXP8oPnkPBa1N7/qiCn1PdsswIGwaI+6CKlcYnhahmQI2dIjrtbpqLbsTaxA/y/
JGWJkN92J83zCwTp1a45xh73gAPCf/fipS+GKKaEBVQG/srJVXZ4OYfXOlkkbDVnhTAGorh3Vv8r
Htk3bag8Mc3xTvSu2PC4wqmYfd+289SxI8m4K3pDEH2ton2HSB05lZcclWtHQO46ZZK2whfTmEdX
YC4Q1aHwJuiAjF2nbaRxMF4GXU8BvZahkzRL/LPFIILO9OUDJAFGLUCa2nSDj3Kd4eZw99/1ulNX
fuKvYGQbFlBBMbkBBLOkL4Oaa0M3yHlq592XGXNcaxb7B0tNcRgOXfHw1EuF4y/ao9TyE9APk9HJ
iTTJmU1rLbG57iKVtV1040I2Kqq4o4Yarc2KExH3Wh2Dswy+orI1g+D0TXRFyBz4epOVuSzNwPKD
TSJN831PAaMx5BCGceNbxyNlZ4ykqqbmEduL5JY17V1aX4PDqigD5MhQYuaSUh3kTarvqKiFU9rg
ZRXrQbJSDTOyyzEPpbkBNbE1UHEUhVBmQop3w8KsZ2E8PMA7giY5Ujrr+o1jG5dz5hkR5XwMTXNE
ohdCFYidvvHnKwg3IFidcQI9prmIt7JMyLftl786Q1viNJKjfqOPo0M+l7/a3Z6ZlrthoI9sIH9y
5EZBRx07kraRi4ATsSu0CXkLLp2Qdwn3fP9M4c2uNIjh3UQA8H1nQvKB7Quj1J45tsIbhYLq/iNG
ym95U1Zx7R53I5pCYfTR+Gl0qGV2C/C4uJFqjcg1cD/e7zPwR3QpaUPq4nrH+UXnCR9iKFT1J26L
cJwnbIgflda668bo9tM14eM6VXvb9v+UBtr3OejV9fsQ4tYjgrV75CxjAHBCnEIeMMS9hQR2RZuW
MtfuHlN0dQBceBposDUyMxD4JcVMET2cMHYk3+e34FHV7Nh9rXXqMqc8Mbe3i5Mk+Vy9cHgliga1
ftmaVI0+TDk2/vLMoaddUp9AqG2tXNMpnkIpsnxrN08Eg3vRreUPc8SkH1p3toQIg2qEPg2QMpeC
+NgbqIGqpw9XsrsSHLpv1p6W/wKsWLdLAcBXrDSEcy4t1epHYFNCcSaSmSBpfEE8Tc21pIlvA3G+
ujQPDRMw1Wc4GIy2kpU1EhGjsoVTAJ9KGKaKigohByOH+lCld3nIlkF14VuR3hAIES2v8QUdfzof
vRzunJ7bT2vOKZtah+CdkjFfupPifhtsXWwl7ha6jNeAdfdCHo9az4I2bho5U+8aGQdnhnrtPfRS
Un2sVG7e3DhVtWS3mpmHE8SSGDwYtNot8s6WPjJGMVFX0Q+wRr626d8DELwOVkdrP0fK+o08vtHu
69wqAcRr5qLgkzp6g6VqduA6alBR9GZuf0Db3jHDCGWymsKw+AVGN+M4vfhhFptRiZ3QiCEepMFq
aGQ62NJy1c34mB9YsfjdSR5ALppETWYCFMDEhMXTlL/DXnMPsHhRYdCF1yjNmwObGYeqv72FGklB
R4Bajy8oaBL8ScYkay/gGtESgdLOXb2voUV6A3Q0NdBoRO2SizpsW1H1VvnnLpq37V1A0Cwwi1ZK
zux3YkHnw2d+V5T68nqt7GOkgYRw4m+R2AZzN6FhHPmPkpN+dThocaJuwnnEs1YnP2P9sXTHpUMF
fbki0JKptyjVvHvId3an/sG1/ntVwNwZLnq8KUvgxlUhGZhSC6ommVRwFCwTY2biBHH4078MiNYj
oG8HV31ZiurCzgVTyClFRDwMkgWtlJm3Q37peyJtJLi26L3ZHh0L7QLvY80g9UQNhpqKutQpjbf4
Rpnf6g8Bu5IrkV75GFiCfY8cbi+M6OAsgvQToH0gBQGXc+Wg8igCaEmJbKZxc6wH6Dg4lyXsfbDs
TBzFv4531PsbjzlDrq+Gecv+zcReK55sVn4ZFRfSoFiRdWcxdIXNr99AP3HuXnEI/0b/G+U8IgYU
BUv5Lwh5HEzVDuewzn/XEnLKKcKP5bl4I5WXCEoftHn3OA7sIaPvLyDoKNFDKFCvHs4zbUUaUypP
9z2VN8lN4hKtYpWTK7NzXKNpJ3Tz/Wwsoaxo7mf5uld+RPh83+zd2dXwfwzGQgH28A4wYqNsAQ6w
lqA/4h8DYg9y6RC1eS8/4VtgtIT5iBi1di/nYSZ9KeZh2sLHa5V1uUu5mN7vh2bR8BtXEoue1drL
/8BOyk7Llz8zbrc1Gr84GE72FjqvNt8wCEs4Yo4L8HaNRM2Vdbgjb5Y6Pw2Iw51X/awkuFwbHDYk
T3otDgKJ+rWizMRYDyHB5kH6T7jQBZ4ot/AgN8ZaNxJf22hEH3ej/EeVYufoYVMnd3dLCCnOXDI3
KwPUYNox8uPYXV9EysW2WaX7+DqxYin7q7gwalhCyz3fEwsQcSp4SU7ot/gFKYbcLX3/20Bkv1Z8
OrTCYBN/8CtEpp/ziSuQFPkvYAEMt0chWknOuPgzSuzBteYn3SE2b7wP/7QiOp5el2y9GwlfGl6C
L+uGogWYUZwkjpZn8EV0v9baBDGn96udPVsA7nUMEcgnWfS3Q0kKLL9w4PPW8M3mk6YIAe8KKlSs
I4waeIQvLeeALZetIuG6MoKdOFb8mIBP621TwBxyBzgKF8vk83v4m1O0tUxbhqRasRo6Gue+PqYD
YSQR72viGPHCLQfrXcn2nC2e0mpNtaDPKO/8fzgqLVHdqJsZ2D/SECB2avRUkbixoTGhnO53vSdc
AzttlZ9sD36QptLjyN7i9ZNRo+RBYqSYWqivceUfK+DlNBMzGdFJ21YlDaOA1GfqX9YJ+V2/8+1j
125EnUV5J7Ahg5HTxEI7jBm1dNvdO91v2SMsn8tCE+L8uW2NVTchuSGyCXNqpO3cNcn4lTYrO2Tg
IhhbcZ9KhCbyPRf9RGZ4HauOGcOp508RCxV2hZ28PmKeWeX4Fa1s/M8Ud3NIiPztXOD/Q2BFhKXd
yQIvKmCrgC7FGgioQF+V7xq4hNHkqHS032N7+dqDla19idIgekTZpOvx07LfLh7sreX/bkCYYCJu
9DOLSJ3AND8XW7dE4VgyW8GbbncJ2TVeqASBo2qnXuWuGq3MTRAVI1HBXOgN93tw2M1m5eHLPq/n
dWM2h16MdtVsz7A3OtAFxpOsZV1QU5wSZLHiLZz+HXkwEBrBbHPzmROkzZHhn6xf5MUUHcRwzJi2
Y0W6ZNfDqTEYGYNk6QflOpTm9OsuRa/VaO2/EaFrMT2a4wAR+FG4ThQ+h6q+bsSV6qP4kD6cDKlD
oqGTzKyTUWwULzEponq3WdwKLVNlK3qfN1NWXAzPJ+ynKpHUjo0dqyCFRI+VkrQlxotFADsI4ggH
Tg0EVKn1JygjgtiYsLlwOrSCymaFp6uSXBR9BTnVbjmZyMVSpQCjpbts+Yc5aNc+Riqb1BL4FssA
ckzHWiKWPjs5kP1TbnXI+DIVoqG/SWkuT+68wyhf5y9XMo1d5ZPFsRDwJ3Kh5Z4z6YmR4yRdQJak
W0E1NoLnbtFVVkDHrgY0TRr2Le4nrysXn3Dx3wnBXn/dNdl5DMAOgqcRQMTaWgJw+6SkuQ+maWOs
EdoL8KJD3gpL3Xaj1kEO+vlUQ3hZDvU/9/koAaOmlBm4G90w4gLpRat/3fA3Ik3TMvVFOZot8pj9
tVULp8mxFBAwDrXznDCRsZE8TGKW65XxgFsF9UcSKueY1ZR4TicVoxiX/TOY41YfJaQvzQ45F+zS
c6MS0143prPGcXZAzGYR6sMGcy9YIB3WynEyytwg6l1PYRpXOQz1JM0Oz22EYvuRPlv+aasGvIA/
rHPqFNaAeNQrMkRBfUfkRHVFW8wvo89sT7zNi5cH2gktescjSNznx03FoIKS+PXegh4x74VJksLR
ZJkVBZx/teLzpF8l21OodRU+1upJegfhLVXp4e/c2I+Vti+FuRpk1GQs66keFYWNwer46Cjnxsj8
Z30NKJxCFHlmiXrgM10y1kGEi94Bfe2Xdbep7rnfmZupCyn4zUxCzcdcbKWeAHJCz7LIhvkCBcfC
UY+NoCMTmN15FGeR++XPpAbMWywxo3cjrvhrzmnjZ2XqfcDRL6GqHqar6uuzInBYPRYPqod1XIGZ
UXeFnR0pXjTyYJwg0+sN+FkLy+ZF2X3tENKAJZ1gt8MEWsfGxNYbsIQuZLZf3mipKAy5oL1ztI/p
VJYou99GX59/CWrpe29++J1cVhRnrOCRS8eyAq4KAZuAV5Ro/aW30w7vGNxfYFOHMVijRzaSLRjX
7PpcHMl44an760BoR3RjWL7PEUcScrrTHttRWwm2NxmB2OrNK6x16vC4AbaV9BldB2M7p7GieIgU
lRc/CHrHlKdqz9mY2K/h2JeKRRCuwXjDm9hbHbEBEBYEyu5of0KO+ae1CAy2o5yiNJ2DeIF4e1Bo
PPCBi0OmVe6b0jUtQW0FgT1RJ4s74UTyK6427GdHbY8c18uO/N7d2+2L+Qlf+hMplBceQnjTrK4w
8mMN+sIFOuqHWhGAgFXa7mrKUHE93CiUtoTHc0H5MkDNeckfj3qw+VtcTLOX6LEWVfD5Rv9jgqVx
NgLVYedLFFfYQ+T57/s8v9PpNdOAgi7KD+HppCmDmPAw3TcSzeHpNZ712sG2jgNs9bcwcjbHy5TY
h+PwjWoBnbIOya2ohLxalgJBEl1dcibMHk0ErZwLo32SblH/3H707tSjBHAcU3iW9T4gXbmtHWzk
zeb1VL68YZd8L2h9GOJbD3xHVuduFGr79Pg3TYk1ZuOEdw/dUoyjGrNx36KN6jS2Z8qscduCjALZ
BymZ+o/WVf1MK6DJjlnpz9DYDipDgD7qVM2QAoHVLDYVdns/c9uZxxs4gXDj3Jvw2aCYpb+5TPmt
1WTMkwD2DBmzkygwX4rWOcu9YOCljX0rNrOqQzedACyfZS5/U/aTNhqOnOMR8NF/sKmipplGxcy0
tjG6Dad+opti+/on0DEyB2dnBCGH0W8fZUxvuDn8TRqDXnp+L54jHAUkGCQmm2Rgq6lc+A5anRDX
6+tced9P+odYdaYVAQ0D8ullb4XCrolr8Rft/c2h5EdKk2phm+UrNIo20hDOCO/+yljM19xFMIrA
3PefUEsH7jbgDZ/u904DHrSVUuIwdDsIzqFoKaD5BVwIDWxzbQF7tQiee7VMYqgpuOlAcw57S43k
kCnpj8I4MpsxVr579t+Slp2dgUTE6r/jlYjk3Uez33hdM3SCTnUsll1Hm51e4dcXp86Hrp/It/by
jD1j+qGxXqGOC1Sd2nhtar5OBAPmsRiBiNRtvap+rdmknlk9rskqoBn9yakG9ViPmMQgLrOBf4uU
1X09bM3N19NnXBLbKDuodSdoTdjjpAq+psGwgOMrlpLA2U4ZSFWg+79ycIw+dKMEbjXrV7OUDGqe
M7HAQIFevr54nTeByvPPvtsGLKxx13CaYVsMUM32q27naV8nSPM3TjU+c8iIR9IYYxhWzPyJceZE
On+2eHgT2qnwwV2/VGOT5+d/M820O2yJIVux+ZFYrUhA8yyKYJEjSyId8Ii15s6gWZX68pn95k4h
Yoji2xW4z3YSaWMWgQkPRz5SAPNIaHabxYRKydmXdo2Pv956BrV07AEjV+SWTzuwSD3fvnTvnwQh
zw54zpgEHpNeRQ7Z179jLxI4OwbdXJQWURE92Vwo4NBkZ9u5PhiY4+MHKf8rO47vtxSC6xHJ8GZY
LwFzSUnrkBRjYO5FhkeeiFtuxj1vT3couGR6kGo1JbBbu8iuuZTWhdN2tiiGy4PUa469jCE8J0Lm
jO3IWwH2B5EXn6vzl9HuQtHmZ+mRapIvXPPhZcmdnDdK3NB+Yy2rTU/YKqacoV/ma3Y6wF1puOb4
6zy8jrz4TI3Bt8eI4kTXatmKTou14LwdBZLgfe4OOJP3JiN40gSqKBstqKkZ5qruwdA3KOGMY42N
wxZCgWmdnQP81uiaIkYCn3b9RfdRzY3a56LsRF4pwgpwvsH+PMNdq6OhFDO6pDvFpE9/ENJhnVXk
gTvrqLb5AsY3OtJiYDwKUHl75oZC1TLBBPwM7DERpYyQlG4nLvWD4z/vqhDa15F9oLp/1tg+6P13
R0pB2c8k5SxKK5wxMR3zadLePNdnr7viKS/bBjMY49TC9QFmboKO2c8vR+Y5mHVvsKy7buJoF9Ka
ZUkMo6riB4KMRt8tLBQVCdYv5u9y+81ANO5nMu+xRvp/tAk9FLue9gsGa4kDuKOUiyZFZyMtpH8n
zAWpo/6h9KhY5uN5tijMexTeHBYEc+xRZBsYmAp6JDORGCamREPp4WC+5EkUD4g968mibiNJd4If
VMcsWvsUd3uAdbT93oJ6lweMzBX8S7g5R13mT/GcLnzOFWIuNQpWS6eWj/HyyG1ns9itrPrrHztp
u2fIQ9D6k8FmxIgtp8zn3GF3F4Lfgh0jmU1nztfMMLLxz24q1EQ4HRMUPg3+vmi9vmjFy/BuZ9cj
qYaf6hwVsEYCvrmLCnlDtanII6O3vbhRc7XkgCQ92atXqFwU4Lvd3fSl5MZt7zlrpG1CNIpDUpr7
w8HiaBmMh5d7fuzjtpOEUED6wePofra4SntsVrTBGgHn95gWHjHNh02E8C2xNhnkE6lO97gevulz
L/7826CfCLjmyieWU9yKtxMtR/BIyxW3d0MUTQN4Yw/C+4zmTy0lo1fJcKDojlydBYvh60bsbb8w
uFjra40zH1TElSE5zFizkL4HRZqItAucCbailzEnj9Z51oDJP3dbJ8xm2b9XB8efJS90Z7NZjYOr
bfpI23HRsEgyL776RNrO7Kg/YeZ6caD638PcRwLj9sxFcXZpooIrrpe/HagceRQTCwFvxYpeuhgy
pUKLWZD65ENiBFrIq3of2hVdm+fVbzG1m4mFLVm3nAPTh2rB+c4ZrNP9lIFSZbIXFE/9G4NFOorS
h18qlwNx3qctOGsNVNUMjjnA7jz6gK4q9ahDwHVFQcNgWKnw7Ayk6koAJqheWKQpwMwHi6wljC7z
nJosG8UI+lqKe0e1qNSxys9Kg/CUw1uSYSGucsIxr/9uOXPI60AxlQ+YKHWTKDewTVh0F+gdhfsq
xgYvzx8aVm9nnH+cEKQNVZV4y2LnlQ5wBu3217brOHrF0ZTcgTfsw1ENPqgL1NitYEAHmVWNDQeS
IfPJeClBi9WuEWN5ujXG1X3RDBwAZd3VWVNY8eluaUGL65nV0p9rdQiqW4YzxhS8666ShGJyCqff
jc3VgYtvKK/HH0oUyYgHzLcgDg8NUaI2kPXXCli4SFGYSmWL0kt4uKn5lURW4hYOdntQMDJ3FLYj
YEUtUYKbpntjxg/uflqY0U0Bik8wvSE4e20Uh2r1RsKSE06yHw4/3UoZ8w0bA+0B5NwMIE8NbNSC
T8eC40mOxnsGeIlF4bld/HqJrJecIoKJMfdlxowiOFpFu+KmRx2tcIKXwmIgi5Kr8jA9lrnLqTIh
fv39LxQ/aoBKynasZODpd3pTJ8i+sM10UxtKiSwGb70mgHHAsTaJTST4++y75AavsTi0cH2SD5dS
4iDPmV9USE7dHQvbi0jdNoCuRIuA6XPYSxergYOZEb/UUYr+iC6cWJ4AdgCc4+1y4bHIok7/K6YC
rS89kT/Czwt+BEesQ2Xu7vm9VLGBkYex/tIn8XUVQ1rC201bX0OXMITsyoWIIeRByyuoh5kCpgwb
HXDgH5dEE0A+neMhqOb/7p5Z7BTqm/I7gvUtfllzFcIxeP6hkw4sOdL2GKJ5ekU9szUkM3HI1Ec1
Oe8sfr6ghtiOuaF8uGil4Qa3z4FIvSWbHZuLYFeaIMx+7tTU7JQyVoaSd2QW9Nks7HGj8sd0kqQH
2b/snz58cEhb/CfGBt0OjSke8cDndISi9UJts/sh1EsuBNnejXiWfN4l4RnXcSKe7i/F9Yi0DDJV
1bB+CqXFB0HwC2r1pqSP30Z8UfHqY4uLGT1mYl2O+pkmGtrVV2TdVyRxgCt/rWW1EM8Cs3LuEB2v
r+dlNMWFGGSbJYiTUY72mklRJYu418zDjzCaeW86buDLWgeL5o+EJLqrDnnGoNWQmai0whaiWZaM
1ZRy7eGc08MveBiZaNX1kdJYX5w3hwRRp4hvJ54qoAXs2MQQr1gW9z5OFXPMYmKyIceiU7fTqKML
mvDIFjQLNbWF9VG+1RPbtejv+3FOuH+wi3ae3QA1i4KN88BQZxRoT+hXTpIo5yxQFNteoNhKaQeF
6jkRuzQWJchtsKDXLdoSGBgOoq9SMXliiCG2gyM2f+S5AdckW0fnALmwrtkPXZzdQ3ZNd6rLlTpe
THcW/900d1hkFFPv/u8De9qH9HbCbnzIogFoZNg0npqaIxkbrGg50U4ZQihMvq8E843MIJIWCEtf
H1nQPpiPoNabpneoS44aH9B7XCJcXtJ3tXaH7n0T5ASFRj+MY4JnqWVjAoeUy2Y3NkvBC4P83hwM
77cWu/ZojyXAlaDm45UbJfDZh6+UdcFuRbTXD8ffGNBtmmizkUaQxSG6t5TARtLP25Gtjod3JHjD
DGycyaK4IgEzFZK6txRGsGdgEF37OP1F6THhyq6ZSMTsYPSwrGA3bcLXxNuOInjiTnPC4dph7/+e
jSkBgQDFlGYf/wFenu51WDKUoyInQAsRQwhMUfAlPO48z8qMsLdZAcjdQSdQNzSmU5FiCxHKDaJW
NyjMJ6PQvSwDvfxcd1fZpajtGcl88XOzU3S35DSjgHodpRtw2KM8CZKOmptRIB86l+375F+Y4jZS
ZpZS389FAG5koJrdxkR/lEPjA6kJbTXmyZw8zqE4imhfUw1MuTOaqE4nF3fSr46XiSVvKQJg8hP0
eddg7QzE4Xyr71p2mAvsPPI4JrWdfI8xegPmzvo88hSWlqM26ZJ0xTKjZuULEglJRSRsG8CxIBKz
AsUhDlrw/lrsM7dk0IM/4troeIQbTA+RTDbGMP3wBwdzgSttDIIM7FZP+CiLjxP2BKzuq63bR8V4
Z1Z/V3AHjwfXFHNwdaYYnNcVg2EVtnbcq5DkRC64KlEQGtaXvh0R5EiVFw3Z7Zt4pvORzm38ZaSV
JjI8yFxxbLUsOFTS/9zno2lzI+fHPzGWUhIdDKXJI78qH9r8b+NMphoeGLZfB5Uln8PTqLBLcd2/
OmEyent8sJrYl+dkqvgXXcJmX+3xRmEQ7TYfhqjQ4AYUoj/wZt5RlO2yVgNWDVRj2bi6Nrgpn4Qe
LeWkTxppQJ3n5vYVOdQhUOT2MOaICF66+2Zmfjhn8Jw4RlfU/3MdDDyLM/mojVs9nPWMb/lZMjT1
HZhsu8jo7PX8JUv/atnMYRLbUTcesCwjnloTZCwZltvHYuNS6ICw9pntSKBHA1V30lHRXMFW9a1Q
wTGgXS/7nuniPLE/OoMv7bXMy77ZEAhY+NvtRhc5f5wUXIvLa+0hK8fU3tDpBhkk4onlXO/WfOYG
G3IRZrYYkTueiW85Ig77vu5G5dqpQRN27ocD4v3Hpy2ckEIZDpbXVHGLWJpAdhb154ybOI1473+x
q8zXktLjT0ogI/HDn6HDkkr2WbYSBPoKTlFYYvq2h41TIbJmEhalCoFKHH1ZgTGPUjp8KkA0G9lH
XwzaZQkHEXwxFaXPTdwQLGzBzy1bdNQzO2pk0x3ZAjIeSNjJaVQTXXH2q39XGELXpH5NpDVFwoDG
XC8qnULD1B86Md+qQ1SqmPIM6HnMUcPDFhXtSoMTub15/v3BWzRTDhtAoE9qcMV7oeJdEjkSan6D
0nWHQd+U6wYXvmbxti+rH1IHaHLy4ku1EpdLNeOn5//iDHE43VOg6NfZ6581Gt3E19q0JSviMQK0
/pq6YPKghG08o2vhTTJk1p2+EGEzPODeDU5o5jAgykmIzm6u+Mhb+THCUUP3bSn/+5XPp20xRpHe
jj7mcQPe/cQRyuhNQbYMprjINK8deOWKjuF707A6n1nyFnDCJ4wyXd43TvexUXKVMxsFesASg61M
T9QXofM2JUEVnYGsVTGthaVzZvO2S/ZCH0JNc4W7VNvMQpAX+GOq01IpfvINoxpuRiRIo2qP7FAX
BdZc3D6t0+LpM7fnP1SZG/wbYuLWnqlQR5MW57E4LjoAMmq8WgJ5JfqzwjjE0Iv7jxRyNMNf/foP
2hwap6kjHswaiHNFuEb081++WSuYsR6hssyG0TFV34NzVKv4Rznn6J6Sh2MwWXrcJ6qVuTmzlp8Y
FeSc5A9ZPizLtygvBQ6ztfuOj9DvsU8bK6I8icQa540U3yj95K5n7xCwtln0mNjSycdZQ9qzXyYK
DA9ND6CYMmdnPrmHiCbEW7n8GwlIHxDOT6BgmbT1cIcSypFMDMGm/V9QgC/pWa6RrccX0bVYgzyz
8t519mSUumpLoDHBigRw09QuQRXurA0X2j+adfafMFBdIyoEjAg8CubWY3DU30FIHbtA9tJFPw3h
6p7Fo6y7mG8rHN2MugFUyEV2/Z96goWmddaiw55XdwsrcCZmq0SN2QOLoctltsO3Ly8a4IfeHfOZ
PpATKO7YjI4Si3oUpSWB5lkZfymV4HLz9qaUurFhWdbeQeqCE7EWX68kT9UZyB7yvJ7KYlMXP3tK
r6EciHE/3WJhxwS8TaD5Sm8Hl6LXw053uPcT7w4qUClGSCjWJAQyV4fCJaL4znlUYcDj/051BCB4
Gn2J1iO9Vgx/Z3CRTgsDOUcwzkVBwSTlWPwNufL41Hi3E8HDkFWCemW9ViJaPQIT2h5Weq8kpSCF
p9h1O4HwWniw30vryVgUcLuw8/CxJ9kX1SIlSIaRslkHYntbThKCY0yyReR/TcYOT2RBWn/tmowl
RlRbMebv+yquhJPe2qEWKJycypCBqZylxMnYF55EbShYurM5eukhA9IBEPGpnQT1MsibQ0BO8Fhg
NWBkb9fyiHSep9b++s9xszxg2u8p8FFrTc1Gjh0nwEADPSs8e43oNBcOucqI4v9Q5GQh/EKRQbuL
Y4PcIYF2a2nXkdAiurkPTWNYots2ugZaN70QxKmujn9KWWWzbLexH/DujAaGLGpYyzUUEhe1BMsN
14yfptwvSWwEj2UALv9hH0hbgQZrJCQzzyVA3Ti8JlwQqqmBErlNlvZ81a9k+jibjBrwU1bT7f57
FOvHLDtnZVTHaCo7HjUcYmArdd5NZqrcHkffD5bMxJd3gfe8YRE9mpxQcJ4KZQFb/pjN4nd6mFkX
c2zJHZsce7kqEa3WJ70YoB3LhiMNGZXs5fg0MGCwZoiWdFWuWOfSRWTWQ00wzSHFHXHF1eApT63i
Zcx6ytF74NPIg9HhuqzigthdPuHCU/sk3jGSGBGJGdpyawFCcIoY43u+QWJYoj+lCTcIkEl07LT7
v869pOfyB8SQntGr7pvJjkJHcy8HCRqkFKwIqx5xZylCYWckNi+iXL07HjM+oziVkBkT3fNLAkEr
eAleZTpYWkw8A7RcTqv4wdwgw4WI2G59A60+Pnfnz+o39bivTc0P8YHx95AirI6/2QvPTuEhci7d
rk0blfaoPSOIL2imag5l56e81uoc6SZmSpS8Q5iHZZJLvU/z1oLm5KsteyW/5W6mwc3p/2x7qUVn
PVx1q7OaAPJ/p/88km2Uan2FEE7jS3Za9Vq7dj6LQOe9+LKmYUTGXg+TALhdUuWfcenqyBJZeIh0
VI2jbKFQbQDXo9mRwlFx7mmUUpfObizRNVUGed85oDkucJZ5GgHLrracNMsUo+OM048dOAXwlO3u
Vv66rD9aYX04v6jGM2L75S4Rp6DVCbDCSBfAxfSfavqVoeivIOXqd/yW67py+4fSdwuCNu+nd1DT
7r2tGOuDhaouNhbxeo0xhi4PLREn7M6C62VuKQ6zlbRYoXaseEn6+zgR90eue1Z/x5KkHaGMeNBx
W6zjrGMjSQO9E/GsBZqQ4xf3hP4R4PyN6vi0ZgXfCTP4CrISYosQGQ83uET6n3aT8NImcfokDAGD
0TEP0tmf/S19Ec3klbWuuE9iA/1++u44o8ay0DLmzgWXSZKojCCyiAz5JwaxaQruOOyZsi2TY4+z
yyzWzxm9cN1J8pf2CstI7HS4R6bqr6XhhH5H+ojbQ9AeUJVCBrxNNgrtDJ6cqZSJ8anBLRrRkiWV
aa9c1XI+vrkMeLWW84UA8mc9mmMZuzkBj48E9F9F11e2Z9LdBzRkvdG2JiODTy0GQtMpffRm8utD
oZacD/HTbmuoEvupn5Tit4myYX5VZOvkknZ6liow5MOLTyoSP9n0vKFY6hmfZf+wAkg7FzC6aSy2
PU1ejZb+h99E5RbBDL7NXMj8EnWqLRScdf3IXEpxUJcgHFWfH6HJvwu3zuL6KnPfUWPY87uC8Zzh
Zs8vLQS51sAUKppCtKQ8S4ID1a6OrM4lklCG8fLm4CFj05anb/FkXyzpAdgx+vJKqxoRcq3+gE5e
gX2q7dcqdkqHLIuJmc9oxPiMqakPaTB47ZPvtMVrGnYp7X9hNbVCDeRWp2GxvTmPrsWzcAslzMk0
MDlkfckA+zAMfVwlVrxB+yuRSnWJU5CaQ99cB9BLSEyJrp78LsuBsv0Akw6LrXNU+LPkYj849qky
629PQKN6r/JfOJWvJElz4WJZ4XHZ8zTMpSofQWISPI2q9c7yiq2qRLhfarUu35uBBZX/6JPPyStj
V3fdwBv9P444fhUKwg49w8p77GEJ48LAM3OAtfjQ7MCg13H168UoNmf6pBvRXCD9tJvn2kDyWBcr
ab640K1fJX/TM30Z7SM+dHAvJ00TfwociOXatcC0jcLNyGwFb4HcSCxYrWMqtKt7sEVUIC6ce/h0
vzouJWpH4V3RBSgSBboasuV+jx1BrJpp5hxPrfTvMRPfZKoaOT1R3bHX+Fi0JJlaYyu/pbWc5tJG
kpSz7DIWLuDLFFa2FETVjUm4poX7T3mlkKc4DqzXdlSgbt8xytCd1wZoV35bVPhApGhpasDcTcsy
g+VmPS25MciSTL6m0tktWYY1cW9o8Jj8YXUtCoQnqAdyzlDu9dXhAhBQmY1Tvs3pzfm9tRP9nPXg
zzRMUZ9zDdTEys6+PFwf06wa/OGTFGs3HMnXtBVlx7UwCWMe2cx0PcZvZH9wHEX3TQ8MjJcJKvLT
WaqQ4oW3x1EEA1CxeTO2XZpxqJdoQWXbOu8lY6o/5TlaseduysiECiv59U8wokdGdPgmmgOWUaSE
0kWxnkqlKDkg0Q3ucVdWZ1Y/XsBxf4qjl3w1D8JznQyaeUdBhTHLuBMTkA2r3ltkABLwa9jIIQxw
1N0WCCM+k9Dtao8NXlcBAZ0R3zIBhfq7YGKYXD4Dxf1ilq5Emt+TXVPHvvMPhVlQIczHOZsYVMjd
fMSqThXAbZO2zlcZhh3K2Ch04XvT7yxCsBUmmTzh7b6tc+ISD9wwFDjHl1hPB82H8IWOtwDEia2a
mELoOEyhGVeA5ZgmUCE9UeisgTbExeFutXRvfpL+ts2jPLvgkyoT83wNFNB3etQnfUxtUbkSu4Xp
BrtPO+aNBOeB9y+TDLQWmfmdB4vNzQOB4dc+0nFZkgBTWDX5n6pypL10eS/Pg+Vxy/Plsi7gOWtR
/rhLFcfyMnjWTyqt6Nc8/wK32kr6pl0AR6vdUq9oiSu4RVQb7YtGoyE0abbbM5CLcDIIhBHEQ+6q
0YdSTufGUdislZxb+lzkcrfFYncNPfpnc65OOp+V/d/SnkkbRHeW/8gnuAbrJ83QvqaElwEkOuEI
kNDqg7GMI8IsOwjBY54v2v1GWOPM+Zg9DQPR2y8/p9fp4sSe6NvPP85nbCtgV3WZnvv4etZcsELa
ts371jHP9kDmc0iFEgqo6tNNsLwfzp6YWc5/qT6Utkl3B5wOg4ezH32nDuX+IHJ6fyfFnlmME6nS
+V0YhxT/NkYdE6d49/uF0os2XD9z/bZ7FTrmsiAIxRVBAhSltqG9vNSz+lwpqrgwaDjZ6QVyv+PC
GM05B52HCUYrkZHB1gdj4gU2VAmpfpCs5KnSsEMZGQbydSmt5UG10z/qOgJvs/+i8hQj3FkrRT8/
H2CrPLO1XFuVPugxd96ntV2TXekjkrGrVuaWu/9RV9yBJcUxsTByAcQ8KkCYdFWYx20dB1q9Lyyd
+YYGn3s1wbeW540S+iGhPvbnkH1OCoPcyR0y9fXSK4kNOoXYUAqwXuVgcos2awLGUU1Mlhgt2zXC
wMG1bKD0UroYupLefuuzQ9pufktgtnVcBmKexZwBF75yOJC88zFVQ3eyVcJHmJYF8ItuOl+GHat0
U/b2jInFfyinxQ2gsRMtKDAinZFZlNqo71DP5pN+Fl7lAgl5XGMau+TOW344yJs1+JwT5woeyNIa
tdyYGfC+3UrSI6Mod2XMtKkDkHBGalHS0r56jJjtha3D0pQeuen+5QposVdf9JgeOQAjwJ3jXp79
43oVulyONVmEhhaKXrZcMcbx08Mq/K7W1gV+GmYXlwPTT1ZJOhf1nJFnrZ0K6hYsnTHkOsR6BBQf
vEtoEoRMuDpvoEciGnI+FBr8goOJ7EAkV4zdgAGSHF5wlkn+jA/vDkowo8M2Os03xrUF2Bx1RGp/
Vtjt1RMRgvCDT7JvEs/89TBZdFkkMyyfB2cyAXGSnJpGTxOBhKQ9BJzswF73PoDKhTKb4PAQgMoI
p5w6h5NdwMkWx93cezaHidgj2h1epOfNPyekw8AZTECoOCXV4BBv0VJbmynAzo6WT7cBMQE7NyvN
X/1Xwbi92TapvoWVKGshCnHGoy281Td5HhbEGPtGdYuzIs9uj4GlvAhD6dEIiJl/aoBIbray+6oA
0ilQ3WBKYrlB0OjHZRmrRErs5sG5AXHg93y9CoqfoKz14ASeqJ/MfXjI7ROlOUL9yqp94YQeb/Ux
Gv1okIkVTHLGyYniWAP6+jXARbbA9TgQBssKnljQjm0jLE7d3ecDQaAmWCWsVJMi1em7VDCmEqB8
TEuFY4zkoJCYyGR4CwK6BiH4slEl+VNDUqe4pDI9dy+xCEv5MFrmOv5xx7R3eC/oUw8FGAe9TfUJ
Mok66TzLbWmSHU1K34rb4/gRXBpXWsJWiua/WybI1pTvuwz8Yh1MSz0qcK+6GI3sW4gRjW7PVLeo
tdM0PkrCxHft9FWrvcuAzaWxdrjVSpeIHFewIwJA5Baj89Cj8R0Nj02cWp7q5z81sx5PklMIbxfi
GZVdc5dk2eGuBzQDYDawXZWpa+C7r6QiUWjTAjFRF/CkWHsEDmdeXPuRsKUafaCrZ6qzabECLbzh
lFlreQXB9qaZ2rdOBrGXf9U8n5JcdcTyXhantNYC55OyGn7JUpxZ7WR1Qneae0tTMKj9ZmleIjkz
2wFmpX92O7ytLZNtS4remraYv5nWo8925QR/6FJC+kFKvaKy3lrCgUd73s4EdhE0VuFjpQR5aEXt
BKv0LQkODS8ZaAqf0IHBF9zijJxM/MEHkUJAKM+a70pTRY3K7lkXXzjpmlCZu/kWO3zc/SFQW2wB
pk2VAv6JSlD7rUjwcKUJCochYnoY8vlMlUGlwfbycBxps0YkIDPbETFB9mTMsbf/6u8v17dQdqyx
/QhbrsCqJTqxBEVdIJDZbwkE4ns9Z3bltT+7embOwUziH0s+Q24Os7wtpkxbORJvIT33fbK3WVjb
Uc5Wyhfi0lPrryip/D5cKqb12a4b7n8l0x8raLLueycgVpr7ww5yINtc0tOH1DhdgAwCDjTDLAYb
4BoyHrO/17i88wR5Q3xH/Gr0ptRvaVUfG5or+owVTNk8sTPH8ABt/q91bjEIvTUV9bZd4cKPSC0g
XfyiCqNM9Po88I23ePKAwvgkAi0Dc/8dx2dkNxh1sUEK+F2UdlmM5J7FTsy0Xd/yHimaAX0/rSSI
xnSYrP0w2BixcSHBTLW8V6zsMjbPWAJWd9FbsZoQixMzxXxlAs726YMPR1bPdM5/BVCzEyASZeOx
PFtV/kkBWnikVCWf5R8pvzds1eLLUW/7/v4cXTZ1lP2khWuNit4xb5BL6N4WBxy073WdEZK0epwN
P4Jr1HL8PNAblepQFL7rykGqAXhm+rO3Ja+vqEcU9NJD2bBe77IIkjKMuGfWnVBN6/4QbPfcHPy3
n5p5EnPUXetnG+PYGylnwjZRCNke7NjLBtJ06sa6NNobiUwXmt/ZOdFN/jTPwNtgFGlcIBkZgDpq
D8FRyTebil2LsdUEFj29Lf1ZVpdIbSD8YSemkEDl2ii9sGQr9qgUKKEWvvWR+au+JAlhh4aRMnBS
gZTtpQYDx91ioDLxRR2H3ykh1fQFho3iqH0yoxnIIvEHifcR3RGb/oZXo569hHAONgMdzip1dk5+
5knmyob3L0irBm2BazZUTx3iEgXu9M/vS/wahB9zVpMxyPc8JRk5SJZ8MHfFll1WdgH3Z2354Zy+
5oADZquGN+X73oi/ivnC2A0KnpNW1efV4IlGwFDvouHPaRyprCg3KicCPp9l0nDvIh4OrTqxaCxH
dfJ/3vZqrfRORYGJoc7NGp6cUA8M2m32WILpRqkAAJQAnUmQfy5FDc2iO0ywnsrYYDjKH5y++FAG
2Ff6UbpjsNlZuOI5yxmQzB6YSADl+WgxoRjx2nlWrgqh+XI9ZfuYXcwbZeIsQv7HtbTEEyVG+8mf
5azAP9nLGcrbyqlE/yfbXg32DoXcBXlp1MPMuN360WLcTSYFe4aPcnKWYY4yPxuuKnnUvAwFEV6l
U3yKjcm1Wx+SomWp7KriMgVCxtDsVBJ5JAinECFUcCYqkJddZaOQIUfz2UlK0RjiZr74f3S0oA07
R2cwFZXyVq+ybUF1s706TZUT6N5porjx5pdaz/eRFAOhmeTkqQmfwhKMxAfVPBAP23gnH/OSCnYY
SeC7ZtlIbcGBJowN/nYVYz7FLi50lemnzVmqVbSvwRWxlFifGi7omp/dA0GsDgGUeCVCTzQj3ur5
MXGNU9vdmRIhiE8+gNfR7EvSxgENmL8YbblCT0SDvfdNv0nGO+1iWotkFUdocyZV3zKh33IUH4yL
1KTto5DE1WMDqhhGjNHlwzrcslQpgI2kfXDsi8jAymhpoJdhniW1VPZpwPafv2XtAa2CgvXsnhqe
JoOF9I4gievJQGEd9AmlvnZv2VAShDLGkddunBo/7K73fnIl3eD3Cdox9yysj/7LUcwzb3HZkTHk
gefAu45qKDPpZrJrzPxdvgqzMb/8g90PndRjvpW/jCHwcELVu5EuExDhC0xOT9WO/KHxt9XQNkBd
E3KXxens01lReBPJHsWpvqOAeVQ6j9GCFJ886ScLlQNhwbGj51xyLJCS2ZRkbo4ETOxyv/x2tx/b
1fW3XJoafVfv7rO16sntQ7438gImoW8VKMMMasyRD3rC5I80CT9BN7YyIz1ReUePyxMrLbMHyqSe
UgYMCx/BwpAOL0DevN/ejHo+LuUIFN8g8nz44etDO/IDbJak2gIIhvDv+lHWIcdPnWWh/MYw4EHG
AzDkO2uPwu1teM2SKgcVdd/C/AGsWzvKMg5L/0aCCkXiWBH/EuRtrmKNz0VLGkH69QuDwql/PDNO
FkMrprS/mz/S+6ZHuSpkYbbSFuHFJQ0vxLjVu4fHkMeeQZdl+CgtP8J3rrhc8+NM89m+idBCEtTR
363RE75vdr6GupSyvD4Nn7RkqSwJpRKoreB+FxO7Rm9kWcfkExEvmiMuBNpYRAtfsSkZt1eJswOb
AYO/g7yvyU0T/1Y5ZpopJPpo5tDIW+VVO11P1D7S+WEv/01YdQGBMIAc87dT6VfLI0qi7KWFUYM5
JgSRWDQfLmsSfrS3o13Gw6gekRBNSK4TRyY3pwvYdtl1XMxdPHWKgjwvUcUGqO0iXhXnVVrMqG95
AG4JGSygQUpgsbxfW4udp0KooqtLngNDbsE1yp82Vj2lGBJfwBQwkPl+ATk/kI34YMtjypRhUw9C
41H7fGNSA8Xdf2Uczf45fwawQj45MEjjRWESQGbSsvCU9uUhQEYLpaHcYa+uIVugDEuYLoUwPShp
4lKDSdH+Y6W1mw/xnCwITyJL7aN+UHtDN4G4ntbK4Rv4cOgQczHFzHXk3tT3FTS8M140vQSa36fG
Rzb41zwawR46XAYQhnfWoXEcNELZZzmh+/raVORPHsu+tTnT4hqFutGpoA94Vgtw4kAU+qhyU8an
MM10vHeIh1WwWdhede+JbZjO9iyvFljm4cQxH6s2hHAyjIGSYxqgVNYvgCAtSs5bc+ik1pe5QjIK
MhMRpsJIuVgwh1iEC4VUjvUgFPPZ92DULKL8vQZS6Af7CxcZHt0RXGzK7sAe9PVZWZlUfEPkPJvZ
u4g09XGR3o0zCPUcNzRrGSjgrLY0rWNIst/pamwaZCmUiJzCzzHJyxGhU1KoxBNMbSLsQcGKUHbU
0tAQEZkO9RMdIcMQIAZFFBmuAxtf1z8Tk2Q366wo5eDv1M8dTplxX74ryDcZo3K59oUOg4A8pOFw
V4htAyhIykPcte7eS8GJ0ZDQlooSQeWruGwNfUhOi/Ev1o+iIAn4MplBjiCoj4pXkNb41i1qiPPJ
t0qTJArcQKjam1ct/XGlLWrQzDhq1xJkheUSTOvydkweH8zj58nWbntGRchtjMMRZ7VQ+YEZF4Ie
y6nGJ0iuijPkL13FSZ/BGMgMWaJDFsw/b4R1irW/jvHADYDoCG7zNI5occVhIOIwsYyChWQoGRhH
li0o2nD/Lf4MhUhb99kidY5L6vBHtoLaBfDel6Mbg0DAdarpMaW4uSSLBgtpoAH6VM/1agVFecf3
gsVz2CguD+2q57kgr4zPV5K7pcAwajQ+1vMbokolZ2H8dqbN9xMRgl2DteD/vogvIm0u/ZxN8cje
R6ni9FZH8RtbRx+LMewM2jxOW96hnRI7ri4oKfXbUlRd4CJDEJCegai6GRXrhRXEBiwi6Dh/t70s
chMaSLti0K16ZSoP4n8hBgR2wdfOesNJqWKCuS8gqlEpUr0QmmC6s09cM0Nb3+bAd+I29Ata8kH9
cv+sWvgPaOBiPvg0yfxqMj8qzRZpbIJL0DqsszzxMY2ifWTSeEE0zanbLY9fblYm9Kcm1R8Jlbek
Qd5azARrYw61chTu0ChblaOVkh7JciS1uu7+poUsvjnZX6AMN6Yy/fitM68pxFj7rNW9yw9JNBOG
jX//y/XfuqWisx8LnVDLz/MChVoJyWE8ASDjKMK3wRobHM5l7Q8UdJkIR9GNrN4QKlZc++LgWgIZ
Taq386tS9MDIZLncutvqxV78UISNThPx1g5rCUCtRsTt1QfJgXdzZptlZC1DGawzUaO3ebI/lzeU
SgmXqRX0P88A9QFrHweGsTVgaouxL4miPuOKw4NKVmjSjGDmVSnXt7zOB9OqxN+rGfSN5V6vOZoP
Rj5mDI4CXXm0XhjfZ1khr89HaYhgSUnW7BrSgxVVUoVeKmFAFvHEksljSGm4tZ+78ZfK7KapfOiO
xofkdki7/7HJJ/97gJFUn1NvRJSTqrSGAIQS74q5S3uJgcRImqD+FJw4JJfEodlYTJzGO3eKLnlG
4Tcsx5vd6U0eG2tlEgJD5q8IOgDJFk7ynCSFi3q5YPujxaBgvui3jEZEoUSmnrL5PMQI25oSqkM7
dy3EON7mt9NZmoeYacfTkPVGOcKHZlWpXbKWbXKDeCLdr/5dN0GBmFtsji7qrRjaG3zwcFdVfjVe
Svbrlldl6zb549L/zKrHIbVQRrV2BYw3RrdjZPdJR/2LQjEIK88UOtG7iWDyqxMcvN7BWR9Ad9ob
kIO1K89rJTCdYsxvDFOhWN//Y0eQ9Rd13Xf89S0U5Dbj5ba0QdKIVCMDRCXhCAdaLj1FXTcTgE0Y
T3jsqLBQE5/8OK60LhjJ16rbBQmEzO+PXpGoOG9SLgSP/jlhb4pTBTMdVMNqThnhY5D0zPrWT8eR
kDQazTMG5V8o4q9/Mq3TTibUOwo+YjZiV8jAEoJtKNHtQ/VLUcIFA9TdAggzCqXGvqjm+Cx9s6kz
sInd9bohBtXgZrOxwsNfLddVsmMqgUjluFnhcdVnmA/2l02pQnUsptBAUIbnT4B8sFOteZ2yE+aC
KPz86PmA6kCoUP/pMqwIAP3CQX+IhH2Vp4xBN+bWUab+cOEpqctpCjb/VKI5DM4zE6sIxVEygF01
e5hNuZy70ZuftTQTibK/B1SGL4kQR6GEkhXOrsMQlkNdOSzTcflhZiv6DN5uKQhBt3V9xD1CZEyT
prh8IT7OO+EPPzJvGyOYpwYPcfblFd/Wy9pn5FGj5cwE7M44eQMCB0LFaVUj01Lni7ZAuI+XzRfv
AkjsyUy94MypRLhSImbB3npA368tMYWywm/e8uAQhypjgEAH1aXbs/85TOQfu9Nsa10dua1Rts1J
OFLKJU5dp2/8nWFvgqXGi7rH7xakmn+AxCuaM62UZw6RVt1FTs79i5+G26E8LZkrwh1BQQFdKJtx
OdOxQchdhhp22QJwCNeXQV2DmysYzSqc7OYhO286smeAfJRVa4+YLsJ7yhK4HolCG4StDeL+5WUe
/yMfrDHf/g5guBht7bKTuXNuWFwJlW3ZpvXOiFWOMPVmNb6OAyrDlOkprE99WkcTQbXW9506H2QO
DusNXARLILxskCgWR7VwUOgsgboF5YBf5S0uPU8JLOmozCMrmpacZdC9dpiLwrT7LB0hTZ3upubG
jWA/bur3YLA6yW5d6oSM7LCOHntSzg7JSwyxrwfP9VGbN8fAOdbz1fsB2wuhQ8qxyP8olfd0nfhK
L/mUZ7+7LeuL7T4At+HWqwL3m1IzL6np5B+ppU5vPeyM3/n16NKhewqfP2ha1PdfBSxypPA2k/Aa
dD4GQXtfZnfe5UmMR6bsHx7ReEfm2zUZAWSahuyIPFXWzF4wwMtCaBrho2xOF5a6lLa7pd+LoTw3
zwQ48PtMSrLJxVkU5mP8f6sZfH4ZXG+xefa0XUxWAAKYf7id8Qv1Oi/6UJT3sJWQNyB1hfhJUghb
tUrV/AtK5D6uHEV2AGsnC0Eww9tiY1w8IpnNSBmWYX9VsDEEKCze025mFtfwisXMrXZHLkwCQDtc
41mWT4RmBQerYB5pK88R5BAZotfzDzY4Ue6euj2S3aESqtA0H4wcTwVJHE819Mwc/U3J9sYmNHlA
eL6qWOn+J+0WP48NzwgbY3yD2gZ3UobrUjpN5hvg2LcotQzEbpwQjs38z6octVabeQ8VYCUwFU3m
bU2yC1u8cwY2Ifbw9zjUT84/qKe+08e0FiIF0H0Qoe4M2BsR42L3QpDvxxV3eb7C4F8pKCFMfLt8
/mTUDIOIpwjuItMdB7HYX/bHe63euq2YtZwVX9/aEpCNyqXWtfAfRIhTwm4UoqdHRmsUhViHZ7Fl
uW/dB8ymRW+5XcTRk9TzbIUyRq5sk6GnRxyeXG14qkYrRGpbSiC8amDQCQTz9XD2qcftJwrqXyxy
oke2k/lPXwMb7bxq38xJOntUGWhAkJQtEiTmJhzgESvvvp/OooGV0NIzDA8ohprzivOwTWkbwlOj
ZmUIzNhM+3vPL/0hY5iU6VrYhGvaQKH6jsQeoZ2tZEMlsGj4YWgrPqBWMC3p/Q4M/D2Z36v/lEME
AMGISUCPLad8pbzNX+qyCx4u1g1NFHQR8vpb0JsGLNY3HSO+1dywWsctFDtHtEF56v3GpfvDlPJs
cJ4r11Z8wbNwm8wIwsaHyzYUrYPZacz3ddF/2tuwPL71awQ54z0n0iDDNze8RPS/T6gs+Zws2Vgq
l+McNgkz+oyabjOOsDwVrrhOyBPpk/t8fxiWutE0KFMZlPqYX2UlHePO0wb3uk+y+RaC4W8SJctv
w38F0niMArEhIOGpoIgiByKugAYNowUkQB+nCzXQt8bG/IwbOndoWJsg32j2PrtbYRlweS1ygUwS
vaX37G1pcsBephzHuH5gJLb4H7WPmWxhRBPvLJiTyhSsHhnOOUPls0eXys4JJKcbrONXajxzd3pH
DBdi6MxP4Z0p4XCKfNrX5h/yXcvRJBHl7HEshGZxnelYHvp7bFgzYHH+gh2oLm9+j8vNxOFG7kxO
b7jCUcNCGBppyLeEsTFtm3WPRAqs+H3DULqGAT1uyE0JgBja7kRZWL4QhU6VD8APG6hK0FFwCZ9D
WACU8rEMbN9cexluoc/KPO/Rxle1lkb9iO/YC7PxsQrl+f80B960gPUhP+NlvJMJsOCO5+2lcvpe
V7pg38oNEfyl7U6YWDoV8TRmrQoPMoSJ762vKBEH4rQNpavFXJTtcjz+T/1iKsm55BkwYU1loRyl
vBIBQMg+TsbXwvggE2PkwLpzUj95d92y0sVC7w1tI0H/tWHS0peIwn9DPryjSyDdzJpfKOYGIqM9
uAeBJRAWlVc3aRCSNAievq/jtVCkRq6y9Kjmd/L+GVdDZCTmTGx/FDqRQl3C6e5/6uw6b3FhF60Y
eY7E230yUgrjkMUrnCe1f8OShxKl0A4Vhgh9EvcwO/cr99DxnqqFVsBdBn29UWYDqr1jz7QrXwxV
P3P+xnC8Q0Ayw7GQDaKKzJZaw4xtFTj4enW7ICSFe91X7y+uJ5xuPbNa7+fM6zhRjhIE5eZNYjBA
LBCvNzLjwGGLmvFUr2gwITAjv74x3VYg+eHTu00Hgq3DcGsje4vWTyR/h0gzUJQ5BbHJ6x118yr+
BZyzKXU/YLZz9XlX7MopliZz51E1bisUKO4JjlRTgH7yJbc4GWbUwyLog8yToSYvIzvVLptM2QM0
mPH8+UYj45qq/dIASUrIfAs/YO18qt34i0xpaXQN+lfuI4/Fxiv0Mq9hgQbE9sA/EOFJNIOIOjDT
NzgSDJRoNkKlSglFsYmlByr4o/FRFfbdhPvnLpJP/Lf4TszA4BQpfr/jmJmrBt/SQFweQ3l+z6Fu
qo/7zbAZEYtQ0SSKTuidfcvyQyz2XWo2vCNM661wBt2cEBBJgaWp5WSUg8xbYAQyT4IK2DEM2qyQ
f/bgUphI4KoPtfet2e0XOMk+eSMPbF+b33yE8XrOeux/TbItktpoJQPI8wNqGTxn9lIyCzn6xe7M
87yWks0WaEULPGUBGFcOCxBGtONTq6SsW45bUWLOqeHKQiWIc7mWRVZsHsHyqPU4JAtXApmv0hj3
IKnWBvDGzAQ8rZtWTAfMVlMJUJO8UVdjegcA59rAWxvIBXsQ1hVfYKfX9S9j1x9jqt12ShJIzqOR
47Y4x/AoXsUd1bnIw4PsYlB+eoHSDM0S9nccsvbu76lj4WBYIJ/WsAYZe9VGH+HVUbqCb25dq5NW
U+VHZEYoA441Kk0oAk0pBuLU2JUyhqcDNQCxTU/ApHKWx/4DJ3R0U4BB8vLRMgfKtJu3xlYI3z1S
UcdFKGI/Gzqf6BQqAM60CvA82UdTeNA5ncitiq9bQ9KeYMHHQQ2RUak/xqpx9gYycBwTlRXbsDWh
g5SNa6XikqbHnp9XRx0PBby9cuW8UBvzbBnEzFZuOwm3zXqU5QYXBrlUm9liAE25fYkEgOTe8KTT
T5EubWWw3FbD/lamrSJAY0nmf96+O97pcwzgUxmCfrAJXYbJMXIcCkxptJH4S6biqGyePPxHGP/L
PI9//f/gnfFEYNWZiT/04MpE741s/FZW0GTulirC/TTyS//9BCpAz7AuFW3F4DynT8eBCo+ndOlo
yWMLOQlnd/RnPWUWVfeopnq7DIoRcdePsQWfVIR242DxQu7zUzEg42MHD+vjsig1+kzjmgNqBzzf
w02FHglxOpPlj79lwtxwMnCWYEAE9Pd8AZghInB9KyZaGYbunEiQHj+QK9fPKJetEACE6EKU/UGA
JuZDzUq7hMjxiafLXH/m+iDoDehQGjEBqGMp5uYaUTxi3X1k+s6Td5DVUV/v+ahEcB0Bu/6Rbg2u
LJ7QFPQb1gPIwMJQXo8NyRJ8TRBXeD696xu8S352nRdPGGfrlHk3VvolzFLDk2oDzEjH1oUFwdw7
VPpbBTdvD2TQBmhlR8oxqwfSMOD8Y4kCEH2mbSEmLA3OGtYoFryJpv6E427TZAcn18/FkFoVYjiW
fwmW812WNiwMtAKP+RVPoFfsg/uSuzeKlxpHGuLW9RGA3K2q1ZcoyLfKON55zs+b+VHbR45kaeZJ
w61KDpDYu+CuO95EW/q6LvpjbP/7zlM3mFHpamGa5pQYf4Sd816JckNsySbzw7JHHT69vjn+SWUz
MuhDdcwCfkI01qk0EDlvLpYK6B8GL8R9DCnbt3Mo5bG5RsSyMFxC7uLz/ahrRh3ka3GbpaCruhHM
jL4kNT+uF7VxEi0MZW3Hy7piQqIpQfWtBDKv0M+zvg5kSVRroKUULgBvv5hZDzB93JtcLhKr/Lx+
yNtGdzu1M4tVq6DEACbBTvUFqmMcQNzfV9zMzZIXxmbkEJxLoVDgZ01+d5sp8ZeZXcSnR81D+ErJ
FjWHzXCWxHuDpMJwE/pBcTsKPGHeyam2KVnNIxyxludR9FFHEElAO338nZW3mdasLdhzCYBdOgh9
BlHMrtR7ipbV2y40woJzboRv96voUSpel69GDekW37SE2XjCPS+s8leuT4zgTWfgJwKch/tUNTny
v7BLliHo1Vj8qVNokHfOYNk5+xHIL5/JBslW6m9sWgVvh7ZJh65xStbndL8ouedZeWh3mGcOhlES
aZmCvIutHLi/bLahJRv/575T7SYpVDieL1wzBN+fE4UMGeIVRxl1y4/HvgeXh5RCRntEAX1UYxwF
XRX/HYcM3XD46Dbp9jRiVvzfaqiNlA1Cq+druxxcEg7i2lFbhxq6ZLBzUxGRWCLRObZl4249J4RN
YLIcmkFaoHwC4KHX07yQKkHxbMMqGcwkUFJ9Tirt0OMcdm1tfTUqcq2P5OaZjDKqrktn6ZtbbA6g
n25I3Cuh61Iq9GnETzbORx7BF9tj4RLvAS313KJVtaauevFTru70YutpwjdyIhLeo/LOv4t7i5lE
Db1gXD6FuW7zVD5maLe115UGJEuAlXC4E4xp64DeiRbezxl8c+xCSwlq+3QJUwZB4Ls/PaGkhqE9
FppgRv0jXS+d+JKbpDspDP+OMh4DriNBu3aYVa8r6rCSsjCYAEJR1R6aj33vH+RyNRIpcEcc56Yj
fXA0nonZ22Y003Af8TMFXH5KLvWjsz2rzuFgHhBE6lsyMwDkZGoG59crlBmWyjyCxvS8RmYRHBS/
jNL/NCUKem1ilmMd6lq971IbnsWRLbpUIZlD9q7Y+cI2t1JC5BJT9nCfr7vVINeBgi/my4cap6yh
shgkCwbslXSt+4TjwRcPYnJB+lbZHSt9mO6LlqOcAQ4lY01ltIZ3lWWsUxG5Mtk05D+JHiXvpmZi
Zny83zsHJzDv3MOXxGIK+oRiWZ2Dr8QzzZsp56tBPiv4V2L/xF1sIzs3W7yMB1WpEF9Xml7EOHsO
PPGVSz9bPhiPqc+8RqYofZBNOYzsheziXMeDGNyqeWqja2BPqB5LV/MlgMWoh8h36QaYXlEyJVbf
J0VuJT3lDSaz8wwoWTH/hSGmmYNDBAvTPly5A4psBpvi4zcIdOo40QLxeMD6xhleXGZc7U4+ia5s
ApKmF54ut5F2RGXj43L9GMz3GFW8CcB4D+GmLzL2AikuIrfkQsF02v7Yj1SRXdOcKS7PHC4lEvWg
VammFSApVGsdbgCysQA/pmlXyUIqDHyC9+yVAFUDRWMaq26twCO1ORxDOxMud8HF92PLVxShK+1S
bzt2M6pDBMYL4Pd50Kk5XzHRj4Wgy0jwI/r3ph0aAlQf+PwOwu6Mb0blzl3KSNmwrkyhI/Sw/uIj
HXDImNm2oFoqbUQSl3nTZA4N9E99uDrkGakCNnNuODWEUzgCPyFcOWO+ewDBiz4cFDq5FCAtVtdM
BTn/yxYBS86UGgIQrH4nUxgno0RY1HDNo4L9Fkli2UtXR2Wymx4X4JAyY26P5VbLYyYWZA6bk0lo
ntFTL3l4+rnDS8Y153Er7DIxzJia/FtRlIyGHeYYkT14tEiLBuFsBEEcfZw/6781a8RKRcBAFIjS
mDfDQ2sVI3ru42K4p4RCN2bQ64a4CBRcOzoRTAowX+jnFE0noHZ79ctrYKyLjyhZHya2moTGlzEo
aYB/RrvzI9WEY8M+VquYFcPUASKHsIoG1WwD0QonaLGXqJgX5HobaAZnkpPG5xtz6wIXO6aYD+KB
bQtLdySBYZEank3VoOjxliyYBG70kjc1poRFcG3Ciptk/eiJU7yPzuLXNPF6WvD2MLCdMrBEzeN3
aDguCqZG8+MG+EFU3EmVEC0uoZSBoMDDtWTLE1w59FsfYXSr8Ai+v8Mk+c1W16m2tz2u+8YdxNih
G+3Rk6ASts1IDEtR+hoBBhC1lOoY5DTpc7rnfWxh+C/380htT3cPEbdp8G1tRnOjMFOz8dJ+e30M
5T26rZxnxX2hL9vuV4SMtYXDDzIRAITPbC26UlbYFNz/K8IA84vp3so9h5cfdIHTE+HgBqv1Z2jr
NRMy9Swqz5St1WCaptDRSkX+jx/SbLqDVuHUQJqhnpz2VZFg1BZuIqBGjl5B4+l2BW0S98NIrc1X
pDefc+hZzN4gXsBTSXXv4rutSkIiajmnBGbOlqFnNfbQEGO9ZEqDXZBrBrmxawQ707l/KLDG+lPm
nf0XKLbudbzyJ6jo9FABope2YImQO5h9GwPbdKdwyC+z4lF3/QB84XrlAWv58tZU/zP/aGKHOtmx
YTyA9PRs/QD35VA2f9ylnaoqMk93YsrmRBjAfOv2lEh1hl3GXvdFNvt1DG3eAQep8Rs5dxIL5ej4
q74GXiaJwTc+7gdYYiXQBJnc/tlVbzH52Ksn1t0CiWqXFIKGe0kA5NkNx3CKxuuzPF5hiwAKLb2C
ng81jdMyXco119TyDDKFiCqS5hd+Dua0qWSMNbc3aMuqoYpWKj314a7Kc2Q2JgxiTq1D2MiAIutD
bxhMKb8uO+lz6PkDpSzWWmMdHZ2XaU+QS7w4ByGb/ThBeGJf1d5FYMCzZxEA6IHktjjRopG7inh6
oJtMMfIfntwQAQtqmKbwWgypwi11TPuYNu3K57Ct2uiRvqB1RLy90ADhTGo6DZpYIMZ5zUaiGFO0
F+D9lFYgniKzshfDM4rvubFOOTrVScGQ+wYoQNcmFAEfDM9xsbfAEaPhhLpuE4hFyv2kQQYc/F4i
igGMJGxSV/EVhf7yZtc2rgdGJjt//DS4iZ8otCazraRSuiAfMERXDy2qLIRfQrvizv0XoidSL0hT
khUOdTiWh3N9RcmV8sTEQm5bc09ouZgUHb0Ji/4YJNqwNEZqF1O0epXAl/gz6CMhFTOJEPBVZ2MO
6vplI1gdXcU23peA8Io9tGIDGMMI74cuWe0rtEunecobVDSawjmjmLN4q6ELnYCT4VBzZX4CR0+f
OnjlefJgfFYvgKoMwAO8NOMjyd/i4+fCmtDRY1P/1w3Yf8LbEBsLs5ArFpcnPIDBJjIufTQPIPkg
LRjeoSrz7YkV2ZrSlvDIEa+BWNBFphcr+d+OLpAacAfLnkrhgJu8qEMNZQooZDhw+XFlKpduNJEc
v+hX8Q6sH+2pbusHU2ZNLVOBLvB3DXM6fRP2+cPe/TO2d60m/CUJFvMfy/TNtRsEFwoBw/IIO1ep
VRi3fl1ZVg12Ep73aShhiAADFU1hL3LBAUX0uOXyiU3znVa7i5APmPh/LIFAZTMOMhQ1ZKRdSOt2
EXA0YIDENNQLrCwNIeAwdVVlhsX24gAEk1t00kzAvdGJ2TBs0lo8RhlVrvddP6wJ/xCDKJBgUMgl
cAiRTMehvAngOK3HFe/lC6Y3oaMQJ+ly5v3SifGZHalQF+BQIRF+AdIEoLLVsz9q5g5T1cq0fQ9u
zApesJ0KuLDtOoap2hpF08AwPa21t6PNyNk+Z07dGEde4L/oEbVGvuZODp9LtHepSl0zstnH70CF
Y/A98kX0g0j8Dxt3px2an3VUJcJnTGgjWz9XVqpzZBYSnepdI2ph8jNYsqHaZz922Npzw8MmR5jM
Zgr/4hbJ9+HvVVoVGzZr07gGUHebi/dUMLjGrPquas7Ct/qL13UzkvnvWNhhiheNDXu7fEYb8UJF
YxgCTdn79/cA7G5RyMpMIZm8zg72uJPUPpbyqd+E5Fx4P+cIGI4/zfyuGTx15WJu4v2S5uW+W/bm
NfiipVHIOEMUh5cwPs58dSKjbqkmDGIYY9/rAAr79aFI1k9NWH3k6nCgSBsUlz198SYnHf1X8+Jb
3TgcPZBthHz+PtY98Iu9lcsgTCsyfklBBP38WcryXylzZH+sfF+VHSIQhm7q4kKuUI0BD7KTv6Uv
6SjYO6cBFNdYtzkwRr9wjGNuNnoRYeZqabvRWpnVcoAnndEXVaMk/RKa85x55j/k6YvqPJUQ6AuP
1dOUGigD3kp5u7Z6jXhzmYGHc+hts/8YztEma4BX9HU5HeMYo22XTNhc2fefYweUwyJD3Ftx5KAp
wcY3qnn4ut3GtHc+jKELtMAqimgCYenFO1g90LE6zijiE3Mcytc0LKPqjoa+PRGmwlRHLPbAHQ7X
Uun7zuwuxmdlw/R+9G6MVTzapZbKnLQv+pVa780MRYvmhFLGaIEEFP6Q1VltejHERTA1nCU/DlS4
dnUwG8/VS9Nl7a168KaMooYY9l89ZTA9AAOfsoM4kw1e9wGmdRe286O/CW0+d5eJsdvHKaAfP/zn
U9YCGpHwpeMQupCUYqNQtu5S8P3Z2l3iPnOJjYLc1BdHkISEPDXqPmJopimRuU+kgK4mIZrrYWaH
NurapVgihb/d+H+XhgnFQFyVwUcL3JL6uyYgapHJ+7FjDTAmoNyGk2+RG6bsTqYayZD77usLKFip
Y4PSINybKM2s7qYlpfkC3Rw6mlcdRGfqHNylLswVPWDG4mfDZyvYNhi2SVjEI3wlzoUwUhehe3LX
FyGr47mEbLApr/qaeUKcmZmZgs/wPOawA3MnHtYQtmh7ihl7K/KAHarVHZg/cFh1/PSnBr9cFJKf
JBKignoDQ6moJ6Rqd6znAeXwHIGnhOW14JnEVKlLrkQ7Fl1j3o7f9teY4MWlYTEdekx0gR3Yd1c+
P+FKaK4syASKOKKVkoHJdyMXgtSvICddo8sx5qESUcmv7pBt/sVfujO/hTlSNkyrKRKr/HtRVYMA
+wlWWTj4Bb6cQzckRQ9M/18YU3Y+8YqchIcgFaWSkOMWZkPgN1JIJWXX1ZV+CmFrfzVRpLEOqMuN
etcYtmyRy7ZR5p12zbpBecgyxra7qSb4H+Y+v8WlhJTeW8B1ATAY6x+QoF5eZLfPvdHWTcbPxkI1
zZyREh5T46QTlnmO8gxIfCu+hp7yMaOF3eCsuE4Yv2YajlKa/g8QTKLXV4NOSoTe/4hlNKiY1KGF
ZFfPgxp1HE2v7UWxffBe9cjw4BIZfiPuMQFsGkCUfBuf+hu4pECtove8H1UO+fRu+dmjtEKBlsRR
vnpdjlMAhgxrD6ljc+fWEIo2GQZGTGDaQGSgBZyR34c+H6Nz4BvB+FN44MOXVQD19Omd1go9kbe7
8eSst2kl/+n2ZMVtv0Xee5LUWbdO5GHRr0StvPERdI73CJGvZ5YYdOx9zq7wpHURFvwoN/mph4l4
C7ZWG9sx/g0KnExa9uxl4I4Rnld+dmX+YLMTc7eBMs1MCinupAl9jYECBOkBAG9nWsZXHWJOCITA
Q5X09mjR/zMBAQ+76992aIQ/Wx/W0ZSeJHnVgn2GHY/PkxcRvoIbOeTxS+HtbexeJLLpxg/DCRFU
rXBNVIkPF3Oz2va2lYZoNxlQPi/D9+DbXvsIEPZ2ioRQKy3i0nIfKmBoRY7wDG3hzuymjkANY6Ho
gHl7Z03co/kXKbQFo/BhB01QF1vB+zrgGppkXLJvBsaWgTqiBNUNmNp5k/BLGZIcGntO69ilcaZl
6URQ6evfBMeeTJkIYIiA/Vg/aY20/IUzEPlpG7x6HtFOHMa/D9XwM2X9Jey/MnfHLvWlZMXni5RB
2ipWtyMhHoxjh83EPj1Je/xY7u6xAtjjb7N6idgqyBh3LFP2jATFGXw4O1BZvR72lInyJ95C3zhi
pSofp+QYl21LunA7KlSgb14WE2xI11i3eQQ9jtWIBwRFWmCqDpXQNez/NXi88LPy1XHowWSiwMxb
3ba8rs0wXTz0qqGsEg333foHw75HGwMqoNXrzegZJnvVW55/fdIm5KOc5SXoLFM4Me5Dx0wek3No
fo3+w9mxGncMvEMRZoRLQR3HfI0SJABZA2C3waw381Rno4QOryGztGKuEiNLK9YzpNoK6815IbI9
IfXmHQKr6y6pPdLZBBTdL/W2LR3aarKYIh3QAK4Sp4lwps0aHA6AKnC2jaPUYhPz0N7SOoc7fESU
lQTXlfkYDx0bA9WkIqzpfchpvdxBgllYUTAw/3putJOW0ox2246uX61SYvPsUmyyfK++R3spxWqm
I65lScjvQHeO4jijXQqm3wCnNAqvqLVbevXlVtBErJDJerVALBgpD7k9JruP5dYmwxa7T1jIfVNW
7b0gteHgA78QyO4w+5Lt1dgnwP3zVgFNzc/y7rrw7LKu3n8PSvwmHQQSkDRZ7I8UCT8RA8/4zJM7
a0+pVzThgAyPHV0XS/4Z18cI6CjohzQNfPNNl6smJVWCvbuvO/NGZXuLHTq+jPFtGnC6gUVVxFVG
sjAl2kHNRwWiEebgqJYEgV04ybU0eoJz355YHKU3jKJSxx2WwTl0weykMYnyYOUqJpS4onWqk2Zz
VI6ldNXcqqWGGpf7JlbOqLdhpEBn5uUJGala92DYh9RKvl3bFpeqPgb7h3EtComB96lxWtAtIorS
JaKAtDYH8As4VgCAdrglNAElV3BQ2CJfjjFt6DCLisve1D9L+6zVa7IvajyzVNhKlc8Nd/eQtQ+P
OJXTkT82PQKvIWABp13YmQLn+dV+7tkwccB6lLPlQXs1livvQIbLjmgYSqhN57beXY5r/E0mV2oV
3O9ApFWpV/vUmB8opY1t9OPdv50mYVkoKoMgwbL4ozoHAqz1q4OobSKFhW1m8sp7Kx6wYHZTLaZH
rrwaRXAel5Uyk6goKXQgOBOLDSqWjzrB0oorbknjJLcDfofNhyCJJSnsjH18oxbw/ZoUEdZz7+Au
vRbnYt1YzXjPAxmhwMjv/1d49qzrh2a37zDBek3KwpITSJKHIptEC9IxqAqmyAfTcDRHJpOdP1dL
DuVJ1jAc29NIZ2+KnhaqUxiMG3d3rsOoGa+TQVrNc/R3ezo6zBkktO0GiamgMP6uWESO2OHdLhRS
wQwxFN6zoMWE7/qG2J6CBuvqjuusrGEjaWPESuea5XYyLK7RGGoU8ojYpiKO1gthQcQqRB0c6A5j
wh+PZVgggmVtkE8rk0qKnuV7xaa2rW6nRChuQsJpENcs5chWb7wCkXPvPrax8tBm8NPra+fDjP+j
jaVCuHoC4VccfkLQv5sJl+Yhoh5sU7fffPC8UKd0AeM1e/coS5MSIRp6vDwFXbz06reY5DIjgPTd
bgU+ZZrKl2bSUPBBUa+Q6VNDK25kp9E4jtDcdt+J2Zsgf4ZYJm0q5x+1zFPq5dDSfASE9aukThtq
meZkPijLiyJJkYm93WiaR2i/qWh1P40ZNLsfkU+XACxfRIFiXSR7yhvsWHXw5JSNFLMt2y6Chsji
3auGCrYmmpFH+V09wcAoxXNzBEUhEomyT+K8qv4Z8KtYkezQmMjq5MrZIjnzk4A/nP2XavfPtqXN
UfhJF/AZfvmRS1zkyTb2qA/41kXQdfCueKpDwwvN1CSvWtzOSstXUSRm7YNJuy+Pbz3G1FFV7dOa
Govg7Db3LmSgJ2lzD31GIc2oNHnFaAiNtp5n98ZGj69z5ckqFneEDLmlGXUXosk1KYq4thKkBTEj
XlZFaHZ6bw7qUZiFxLM9EABbvMeIyEW0Ke5H/yt7vYCY2HjXfQuQCEwwvWy9nABbLIMjr3uGAqdA
yVxazhpwWFG2HuaVSfvHcIqAeG0zwO30FKk/jX2T5j1H28hgDyZFMQNhczqzbJQq7cwk38ovRS7z
v57+zhliHuv2ixiJpOrumGEi7dOS86blFi0RwbNNdDbQPcEsujVhL9n4sAes2diWqgpSuVlN5Hdl
v6fGfNgbGGykO+mWwsWKKl5MSrkNCnPbL62FDGFI8mKQuWom3ZnRCsS0opoft5JMZtHhhnstLDW1
5YqpSvi78Ie11vv/9R5sUphu3QB+ySaso4PAFgg9iSw+nWTaoL0vyZTzCotxQ8H6y91TdzRDFjgs
ZvPtxcCJk6Rk8fcpw6SiSeCXct45GAzyfjoJGWbMwgdKzW5zBbLHMFoKv2x3S69PljYaoZd/+It3
cxzh6eEqwZ1B/xe4DFwtZDQYCZPZbW+EF9qaeL51AYUmJv56zW1tsiuSeJp+tcnZ5ADs0Fzbomrx
8zMAXpyrFeW+nvoFkjgPkEUK6a0cBoq4nLuxirXGZW/D07PcknASEw99IQrRPOP2fVo8E4rOfMkL
+dU7DagOACxf+MWpWTcTpdcaEn4RloXOGFOBCmHb3O5eosfIUM8WzLZTh5rKac+KM1LLJCzMRn9e
Q4W6mvfNSnyGFuD+G8ZKX/sNQYDmDZhT/1WSAYDw86aPiYu2arpSHOrxrfL7+JMZZPbWLIDsLGnF
1KK3PekvM1ysxh7lapzPKYDABfEryAhU/ZxnPuFOkP8McJp/cmrq+umDB9a57aBkJ31G4Pc0S7qc
Jw4yIHaoV/eMvPHaZzpbwg/r+RvG//+V7vGcdfCJl8GYn4dczVjLqVIqiHd26MK5FH30SNHMSYgz
b9qIcrQRwJh2kZSUbXlClpJkmS4TbO+fwKe1/lhX7MCW6uqQi0zuZRF+pHrW+QGKTR10yIKWXW6Q
nm4toAZHv1i7IAKu4SXsAoHIYUFG9NfIvXkYxekZAnbDbUB7KBbxuw8BgN0/pHKPATcA69BTUL+A
d8JNMVkyPd1gJhjsTYD73ktZaOL7k9WXNp5ptzet+cRY5+Z6cAlfZyVw40hOmKACDBFA6eVrVj4n
mEx+nstqKQm24XIZ6h9/52uopdBDAjeY/S3SMhxCXdTROOF+2zeYhBVmT2uL7rgEbOCDNul77lq8
93PPTTIIw4/SsoCpsnB78fC0JR6I0XDkPRKmxfA8ZtsGi54ciJd1UUsDJRnirYF4ZzmPVgfr8wit
v4PbDowIYdXWgPWGa8yD2iERgWmkgYPJBld86eBOf5phmfTELFzifvrj3qoRpatS/JWQD7tRvK6d
/iCVtV7SSdZ0lNKFcs9VjPrRr80a3gEFSMvRRCAWdksTsHz3yV3SW+Z3+Q1rRGF9MKg0/gaTveDq
i4c39lP4CLcdp98NLsLb7iIMGaKrOt2Y6fQG7gII4T7qtLWRcNOG1J7R2xHk4dJhx/CaNoGHnSaO
xO8PDxOH3YuqRMmraRRDu5OyDSMcwkQ3lMQMiuu6dGGkDLLFA6SOszQxNKwCnk/D+XMtNcElHbee
RYLFCHkPgvu2vZ2sje4ohRX5HtCk4jjXN2SZafPzgKbW3L6bZ/5DwqrmFS6uVnC4ScZ0AmiPYqIf
9wpU0ZV17lVdtcK233ukIIklmzFnOz8Cw/ccpgqpc+EJ9SMszYwiMRgCBrrLzMtK7a0DvUuIIKX7
rtq4fwlZ7FPkaoSxMfd9LkknEG9ntKXpAYry1527zAl2FMZ7i963nMNGZXeBkstReJyzpEaye9TJ
+jL99qGWXjFXrxFwv6MW89bYTlcL7FZqyqrbzHErv0DUlKt9G4FbwpieU8hhN5FkzQqTYS9d4SC9
q8dyWr/Kr7+TaRd7HH+6S8KKm6EsZDLKoGtlqDKRKvdq34U44Iab3P9aEZdY6k74Oauvp1FaXBt9
UnoeCS3hvDEfXq9wwhDUlokSz3nfF5dut+oKWMJFd+14lnm/DhpPiBESHcEsbMxipx90PrOMAfmu
IVCTNxQYRSjcJhxwK+ZK+jINt+qLljFUQPEA+t44SCzu7/98qDo/vbsTlNWTU30PM96BnhhyR52S
NMypqayTHLpjnllK0k6mONAonkHwPjGZx51o7Pwabc5j3xIlLHhpce/SRL0v0U3wvXCSOJrgfMCe
okun6+9Sn57wTOF2JVhhvz+gZDh2S5iMlqm1I3tsWr0kwS4oobKjGfAWvio05xnTzZjsC+HSWzrH
reeYCTy81Z05IayWxggLymLmCAB00CLW4goLcMb3IyLJDZ4xpDJJWLkZKmEwZPj5DSi6ET04J2+W
teoT1xQkp8j8vwOYKNTSpgXftyYUzFmib7JO2J2mGkz5maTZj+d8SeF1NW9kBLUPkCs32P6hXyft
PYkRlynY6u/snWWbPR83vfdL+QFEH/qZoGHtyGOTNrD68JB+Q9su2N/oLd8anzopJ4VUW4oEQcz/
xEWCE3xEOXVxVgNVEEIVprIewFYRlU71P/AAbCQgDeGXt8rur0nPVp/1tWqWnweDiQ/9cNil5a3u
EHMCBsLAhn4p1mRpUSwvorOb6nXNjuwIfdFHwLu/xwE7m+SfLsbIuP38LeGWnHD1W8YwSbqQtSoO
B1fdjdlfjedvwyFBeJuG9k0k/auThugTjX/8RP8Wphqw5/OYlgOLK6PcEyeLIacAM3eIHTpmSgSy
hbBgdCwuL32+lcJxWxalKkV715l6c5HgISbdK1SpJo1UwXUuBCADyXmjmdD4PyhWGFxbzLQvY98U
7I8wCvdcTFaMsI1duJxqbXyD+KZ6LI42nUAkWX4m8+O22FegYqCJs+8kGOBncLnHeV+6mPHrpEtA
VJ6VZlnKzdq6+zxRz3tfEkCx/SVlFfK494dmR1UG3yXZiZEojewrliuMdXxes7L5wQS3G9rF1HVt
T6Qc8P2u9HImoJHI2goVqXDGQ2Db66Ydj8fDugCuZLdBgi5n2P5FSoWU+vVf1st9WNP9C7R4Rqby
PV31JCTgDRASvxZGf489q0A9tUNgtbchJ8W7kuU7TPZmh4bXHq6NTVorvTjCWhzOfD3wc/QaxMxd
D4/pwtEgrgdctYp6dP01zIXDOY87xFjPykpooQ+oijSaBzzRArxG+K+zzC2fjFICLcYEENXCBI4u
xW0Tv69E6t3peK6t1v01RMpXzt+2Mz7szksRFby7oUPxhDlr7xWnQdvI9YVkQQkkX7Xfkg7pfiKH
Quk3Sv2M2tAhS6zzXrTK6wDATMA6RgYoCUHM+yZyffcIpdCLPrdKXjur0+UWa+DaBvgCvzK5NOIX
wRPp6sTc1FmM2G+TZ5V6vcTERAAwImD6Y0ajXy02y+2lydZacSI2Bke/Qoz2KYiIw9yt+CH9G6Re
dL42YhUnoigCbZoph4ccLLFdA/V15pdXo5qeNQOqpIBWfbH4DZdMwPYsFriNaviEhUlCVvJclG2k
TkSUeXORDxSv0pkQeXGvDqmg1C0XJWlw1tOiTat2l2ULp7N4EZz5fcCJlXysRN/9FFfO+r7vWQfs
iujmQKyVQsAAPhKbPEYQMIzRhmodIqUrHMomeuC4kx+qC1/r9qAKzM/GcdA5dGV3ix3djGJKMDrj
gvSEqrzMnlFutdwDQch6c5m/rTu9fuNUYxbdoWlTmbnhY9KEIoZrufGuZ1lszoyw2dc+J+SphIyW
w2pox5Lc5AOMSOsSfnrWUCl6Ihd1+Jpepo0YqeYkoTOipDahfCrg7wO/LgN0V+jKg6uQA9KvnQpc
8Gd/ow6kh8etszRYpf7wE79pUTl/OLbxr1mWJ0XGDsoloP+rCV7XVMymJAp/stLo+iBZyPOtANhF
Fj+wUE5Pad+W5bhxv5w03VPIydmzYBov/wJ7mb11keOYlr7umV/r4+IwDQCn4gi3DOxVf8opajvu
YvCYNBBKEkIFCA+v9YavURT3/XG7IaAHhe7cWWypKYqnkQU1t+oF2uob+/633Up46nbK/FmiRwGa
mJWAhqHiJcrpBSIYrNQNi9XsC5udVGrKtcFQ03txX+kEk/NMcG6vDRuQ/qhIZ+GjiX/1rCFiZX7O
0kXM8u7FpSaq2DtzrUMO/QkbXPTlutUUwT2cHyN/JXq8BJmeRNZ8xlYbYSoFtcgijkj61ZtZxC+g
mQmZLcXCpkALW3OK3Fq0V18Vxulaibu45UnuOvMy8KPrPmVIBzzCy/CICU4cnVec8JqgCAGbMWOe
ZthRxzHcCgCAAjS3CSUYHRJ6YmRMizIKBJxAYwWNAJFuDPeGdyBIvyjvfAdiBigegI75CdD8W4l2
cU2z4hOdeQF8NNud/XGII9OwzDWkalKffpFFRpnEoNV0dwKrEasL0zBGMftk5c87xzfxfFFLyKBy
NeESzLFUHcN3L/eELnXabKpi7b8RySGvv/89sc1H6lpNQ27bPNsd5aAz2N2QcULSNkB76BVyO4Ke
ZIhEB1Qz0nZf0fjFLMfmQOTjNDlHGPS9S1UTmFCpNoDPfpdcoTCv/vfoaAhR7ZmknRErPxGBhFo1
Q011/PPjIYoIN9OJqBWyj0381P7PsA6LL0BVuMNnF38z9p8yjB6CKTLD4oSP7tmWHTf3f4ubWJlZ
U65lnakg8HRnhRfO0Bd6FrHTUfi2RAjU+fA12J3rzA7mwfDIjLRvfB0pRXIOkIAiqOZ9lxbn2o/m
UvUq0VyOx1LTLwRbQP+sUjpRgSBKLbJNiKSnFMKOavS/CeySyOoSmxsy38uoAo5rn6Qq89hOLI77
ShoMVXf657FgiVgqAfHy95eKDrwiXT70nwXOEvj2LL2eOcB/rJ0ArUIj5msg9VK1GVcXOYNtuCOj
Y8FinnC39C4AcVwNW4qyVQ3shCvFYNVlR3HRkZ4Hdy+WgyEPPbVy6GbY5QHaY81EN0Ei/rYOxpKP
O8OGJd49UCYwlQ3nNCOTCKiBQ+P4i9w9HhfSvhi+gj+FRCTWbH8UeTWx/I9MsvbT9xnsY0Cy0sWf
AsM/pvLnoW2Sb8LJ333J+M3vMHGOLADe8pOn1xyMKqLgGTAle48uDPD1wywEl0ousbJTywD2QxnN
26jMQX8SJ/4fKxAEQCr1tKdkrY02FMwWY5ElOZGnNmR601xg9ZSgWG/vdw19etZT5p2XUsAvqMz5
gGXWc6vUWf2XqVrxhVGZs7tXskphEkV+YJsajNE9NKUmPCOhtQCw7T1MKHL9IZgewv65ECVyclkm
tnnYcAuT7czH61rYAHR7AlzlZ/nRZoTQFX6N6MNzLZebNXr4/2+o50cD7l/X1zH6T8J/Xgb2jB/O
zAA+C5YVAym/vL50JglqrwrZzRiBlDevFqgupW4zxONonlFxRC22l87b0WSoraiakB5E+LdSaS66
sakYA1cFTXKO8Wy3YnEpiICd5RMCsiTXdfL5LvagoJeLc4uDzUfkeieeMSsm0RgloNeHhyojYBH7
OhOHSDIYjxldBg8vSzaUqDyGUaRpUl3DejDkYCE3qu6czdoXCAflEmDUItw6kfyPxL2+FWY8xZ+R
JbzfLbvaAvCx6jsmedhTFjzMitQmXbOTFyP5+FRIfO2frehm+Ksq3ItpZsH3szg92g+pbIds6wQx
5Feovgrx+dJnrPaJmJCFSNyjdDzDoWQeBXOUEJJJuvVABqhjB1JQNUzelR07EZeomtQJKgYjX55/
aeq7+H/oeM8FK+4gXqYbts+DwNrxbzKnqWsEdO/DD9Bj6jwFMvdAosyb2hdRrQxdiuw972lqD2FR
++w1l20gnfMh5vyjb+xq90K/WPypayy3ZDtI3lnlKsxg0pWGcx/PLWr/OrKxfoxuCh73zdGO9Xfm
s8Yi0PemuNpIU9HpkLi1P67xPpFeSENBNsfjmDmPgK/wfVARC3vII+i4LFncrPp5iCleSxfW+MSJ
2hdkh4S7ijl6e54bPclx5CW986xrTtCPw9AUyQISiCM5CJlanOvITD+eDewGGAmDIKkwqXtug+MV
ObGGFL1OQwA30u0t7QDqlRLTLKE2aCGhY/Enh9hmaebcsmW1B7FSXGqArUN4Yv4EfXwzUSVfCzhX
UZfs8S599S6o6yUdT8GO9yE63Kwcxp5bSaJCN7iTt1axiT31h6I7DVcCj794YhzEQTlZxgV6Ig8I
Wj1X5vmqEBPQcmjx0d2i6qmLuzx8o83/FAxpHFxYy5zht/zOmsLgK0Y7AwkqR7pwX9W+p2Q6q+mj
f6393HM97gK98xn9fKwgM6OPB1aHHXLGNr2GbSTRzxFYSOhliyildk+99jksael0bCQ4buO/NK4H
kw2PBV1Z8btSXhTiMb02EES+XufPxwaKdXD803xkq5F+Zrm+WleL9w4Hv3PgIvRr/Jxhu3rr76XK
39ge0j6sQsUTlJfqvuBqCB8T2p6iRvK3lh1FjJirIhu9LUiD119zslkwLLw0XbUDH3NXmyaIiKDO
xo/YwqMePOymqtwVzuU6gb8D0XXrsnvh4H0D9KgMla8UydqaEOr8kyiQI08Pdn/LYeiSJOcSiHiM
I3V/xvTavNY8K+XK5H8/VQxekYcEyDc3JnhvneO2ICRpnHT35ZczwqWVuZTqFJnJR3OOJeeZAQ0o
9rMewc5x7WASqAMSC94S6owBcgGYnMXITG4YQSSAhjpKp2rZeexfmFhKCRRwX5wXuQpb+ORW/u1C
frUshqH35fBnzhbDeKDJzae99aa2cA+8vRzTql2hs/CCrXahNd5aMZ65K+0BwUqNoIiMDXBft9zm
LMYpH/tMj5OfAeMPF4brywH6qxTGE3z+N3uCgp1AIt8by4ELjOOhcJybRLm2ffykJVxf/WmLii2Y
WAS7oV4094m2ReSXa/VUEbKa4P9mh8QwHLKxvvSCC91DBhLFxbCuU6ThfyNT9ouwd5haBlfc71z9
41kU70/KnzcT107KoLD+wtsPsZ4EJkc/ezb4n4RhqL+Y8xWnjRtwA2LWmzcOJpf1FCr5qBW/96Ya
hMeehPOyYm0BKzG9INxYLqPyMnm3p33EbsQc3D8frtY17uRU1EiF4q1NECCEmtXmoQz7oQVJCXE9
UzAqzzRVg0W7jZ4GbCKqOgkdj7mImu3ci1PAeUZF+NJkSLJ1YcNrW+vTWJYmGp3zUEwHISr1alhD
ghesdWZuOSiam/QWfIXhkH7rfDX6j5IGuo5xMajMDPkOkEbxbnCokKmOsXfzmPSP5nvKtDoCF7Ph
dNMvjBqzVx9vNWwoNTa4pcs+f4raX/MVceLSUJiI78K83RP6Y3gLk+GrpEOftB30ODuyrqGboZjt
ZqPidxc3dWGzmA4oCHtLiDy7emym5wYgOyLOsub27j9HgLO2nlBC5FK9uOXsepxS/YB+fPr73tBm
ZwOdNrJBBhoBp0+irx98kZ0GnPVLmMP2bLZ+fp3vvn//4QEr3aTqoGuTuR2VSozKmDcnCX2OH0wt
+NWew/2ePg3qucVoRd790CKbeloXMoS4mfQpLV2cY/ixpZnea1cSHO4b2XUuwv8Jlohvxadn1AST
3G3C6aZmVsWpYP+IXLVbRS/t5mmG2n45s1XvVewI6+j3cwiFvGkszFUOKhXvHytHqqmA13BM8AWd
uuUEWSOmK5lU+lVdTFXzLeye87WAytxRMrzFxHrnA7czbZKu+/WgzTCGxZIlqoIC/8cl0jWl0k4I
hlDZzMjaWiRJO0p33IsNYffgETvanHMVJPngdFnESUlszWaBggpY+yzwSWrj6OLhUz8HS3hvj3vJ
5gNrA1mceXxfLySWTZ6zcIPMys8mb9zGnTrp/Vuj+PKrqjoI24bgVMbGmI3Nj53qlhOyHTv/NdK4
EHJ+56v8z3MdrsAtto04RMPjEp72auUkcaEWon/+JOHHiOA6vt7Jwit0wq2KC/h3SzZ1VLlWz4Vj
p7SJdJc9QECwc4HWoeml9DNN4snyAwC1JyKoVWNJHYNIsLk4BgfgNZmsaTPq74x0hU+JoA4TUpf0
cFUz/oqObnGv6hdL0bFCHhfKCLeb3X4/8l7cn2HEPpaSvtmxUcwPokvH0wn3lFsbpLqlKgoUbQV6
y9Gq5xw6EZOO1xNMm15c8NEn/JqvV5akaJ47s8kkTKDJlp0IKV8l0TlVCjBTuNu0Sh8lbg0Cf8Qs
RLAt5bFRQbNnlhAJOOE+PYpLepbwZFfRlVXS89f5jrOglRo+S7u9gWnqKG6lVxqDNOpzb6H1LLXv
XxV4xhmVJOQ/y9dZZ/dTXWvtPTZb1/FpC+DOp1oHMnw9C91BgnPrjOi4yAPsXPsI+i2qdUygqPgp
g1JGT6rgPQAHF/eq9hRdjNuFRat5c2xrs9Pj6WCZddmbAydjEb1F3gAfch2V4cxlBjiXNC9Ri+jj
sIeoBEWIXfr6GS4ZLCDJYUWojS484cv4nxcH+wfMY2W12jsABH4vBxGAWH0f4VpZSzHl7/QASMeI
rdfaSIyPxHbdO94+Vsd8ais+WFJ6gUlU/IJboP8JJKP6S2JU2HwoUyuPPZ6VRd5zVRuHeeLdS+cB
GIlgozirGkMoOiL71LUSWAdP+aedF5GXoWEOhtFNEhPS5oweknHOxXzHHlJPHfHsaUojr09Y8twe
022M2MNM/0wjZsiVfe5/6dmwONiN1KgKIG6avhV7w1ODiNlIE+ey5I3Cf+/mAxLtVBUrCb0MsNqm
NU0zO6pEIpYhTUEMpNqJ0ExGr9W3qD2+1DzPvVbCOzhXvwS5gA5JSphs6S9V3z0Tk76xQdWswu96
09MhH/VBpEbRCoUbaOc8UuHRSzi2NMZGf8rMSJPEoc8Vi5bVT+uM1Jnc6HPAesro0VUu9TlS0Xwi
+tZtPwoBoRWKygkDqYbe+4m+Rl8RGswm/04hbE/cOwfu3U5dWXWgGW6+hLngKGFE5UJ2AbSQdxUB
5AMmvAp5YJ5VDKHB61fA8BfhWJmkFLi+VVVXksyLmkiN5gxF/cf0CXSh1PueyZWVt6yugXMj5nSr
ZzPDXocaG06nwSUE3bthuH0/3WbC2fFQAW8trA9mgIqmjLzZECph4oW/s+WW0YtDDXoRWRY58hw8
ZlI/MVmGdZr/WuRxzWYl3LQS9s0sY1cbUVzAP0fL3CdhM2cfTYwSTg0SndYYhlhEbOGBmJ4jKJom
WpejAwlMyco6NkYtVIYfaBKm6MSmjYg1dAmn1GPOxbKFIi4uDuxnV4qQVvSXjTLIkScvB9NWwZSx
b8XiardSDM47EYKFOidF1k8Q9ba/8C+o80xuFRBfGQGauBsRsKvmmDyJJKmVmLXuH04UAE4upneH
vP6Z9khijVs20AYc+XZmPs6N5MI5xdZuSqbXMpCsdLtz3IZE6hl3fGa2VSOyCVLa6l2IHzOL8XOd
hI4KEw085vjuE26pAeDcEz3J2KQE60hHiUu3+XQntRWIYxDKg3ucXcJ0zwgY9oR/PzaBGDHx9o5D
zjrcK7uaUHRbKtw9BjmcYaeJFotmN2H3Bcdrrt4K310Iq25woGLrv//GMYwenXTfRt0YDq8/ZO7E
9Jof8aZkN51tWqxI+kQZLJT/UJwGowv1JTy5fWmV1lRpq0iFLWOUXPQhNGNtwzzbGYo77iF5I1hH
ynUwRB6JtEXNedvwGflj/g5xM0925qENxVMDy3TIOMe2arZZ7lWdRV8a2QnjSfTitjlYkDeqYqUQ
JimvtEKOzIZmJUbusu2Vig0DQ03ioJ7WXjmoSJy15HFbSK/kZIpwHGAHFX0OtuJRHWQnmfehncZE
n4fQ9MfA4sHpJxkxAYzeCUGCWIWQTlesTTrjLibmIMVPjL4JfxBZQqi4HmKH7M/4GYJbcL1Gg8p9
aSgv5PcNzE6Ilq9zZih+eXKATOIFiIju78M8hVX1IgBI1cNQhbmL7PF59TnSQsbFmLPuszKU76Rq
Rzssah+tCoW1ZPHPyyohFA+N+i4ctYPPfdtqKBHsDgGq+rvSrh5X1D4fMNDolDsYKcbNpYktCiDy
dlIQfK/4Ns6Dxcu1Bddm851cUdXj1F1TNyA1eiRnoCpRyS/R7I07XpFFo4Mp7cy1sw1BmHqmYspQ
9YzD0Zav4ObldWZkQU69W8U0B3JsvpH7rInk6M/XJ8QamuGsC9Xykp3Dyj380TO9E4tqlZQeaOd7
0q/BeO0X+t0K56Q3OHDd6rKG6q6pNVUfVBE7zoc4/Qv2dwO3/9266DHkUniHrwdofgj8kECRd+qs
ED27S/waNXH0vuHT6jLfVzDveazmV88fbqo2XgGmsYS0r7PutOiENdj7cRNSdw6vcGnruDSGEqm7
reL8z4AyUoRM4wmi4AMibQCFb3j7b/bJCm3pfPkTFNfNipuxjzNYsPABzmVcxsblAi5JkOo72+eL
xNbuorp6JTnMVkeHgsYQi0abWOuB3Xmem3/ZksCFNqykySVatwIU5Otr11vWh89VqDqd/X3EbVj0
jya03FT6za47dMgk3VOF8Mo4dBOWVki8Mw/y2sdzpOkyt7HodjEdKw0R5b6aVSgKJrIc7XOB2GrV
28olpjvrdcudDzX6+XR2e8lDYOuKR5l3PddyE+L+xoTe3xuIqiubKHaqhB+t7PQIRYRN2/7MFwZG
GDNKGxO7uV8d40K5o+z+cKeNn6drGqctuHaOYVn4ofXJDL9ClnGX+TU3oJIEMhpoIoGcq9evnIhb
46IoMtNNv4duVi5oAjVvTbuOE1ponWJoC5oO+8mNoy5FZe+68VO+2NzP9Kwnrfr6R40breNWO7bB
e6hmUCimgAvYeSAc1s9pmxdMlhaASfjyFKhDS0PdGi2OIrDvkwgu/Q0GaAAsXTHdHWLYDm9Wkick
/Fa5KQbDY70Y0CmXt+3JH3kkZsCta0IpCKYHO4SFoelqeciQVJq9yjXGDVYl8EAZ498+XppKGnWp
tGd2xkNEbTjzvDZ2bVz7EoKgjm9Y2xpXSxzN+R25bZuSUv1u+yLv8d7b0uqaWyyStEYEGmPdpcc/
HfHItWN3pznDzcj8rK2asH2MCDcuYXs2Z6j+O6a8a1hBDcmr0chJbTk95teQr/AL2o81DulL5Kss
SkVnkBCND9L4sD7Gtk9rY6zWjz/DEEfYtFlR9xF86hxyqdhE1tqy3VL4rT69Z0N0tsfBJtwzhKcl
86njY21knBgGke6dz3BLWVpYhCtPvt6FDiwpLuXSinYLoyH/JmOVZjp8y+SMspA70dxIlJZcGUlN
rpcbMfLt1GkXBh3EQueNMIa/I5AhXLqdsBi3JaBg+zlWqvvXhZtowX5V7YZzYqwseeYwYeoeDPaK
diJ56JDyiq6nA/4Ecs4B3BOgpw6xjLPmUb70oDZawzggQ+NK1tn5LjeG9TpZUsPGO+oEJAwkmFgR
Zfy1WIYTrlqioKjiYcJs6y2sI6PCqrcoFWUI1w9GUFuYTHChk4o/78IE1Z1dW78zZU9QNItOg0O/
yIu9lDkMlxGV3vo2QNbiwlT3OdCc3SMo9ktA0naWMqaeK2wvsUHEMAeVJsdY8dG8x81HCWNbP9Hi
ftCNfWAQC42waU7q6TtVTL4sZQg7O+5AOtntMBIumwXqkx3Gs267pnqp56DWMI+ACWWY90F3pm2t
uh+6AXh1eFc4pBhZEmhgeIgJCM3lKF8KXBZCAQRjMbwcKkvFGL5tRNWOkCf5MYjrRlV+WNUfXjN6
hN+QbcJbDbSbyZTiJRO9XK8GXHjohs3x38LfFZBohDlODocZ74v6c7yRaf5VleZ1HTeyZf7KMRcZ
lCJ4pJ5psOr1gGsVHMGRQETAXUT9g6du+AoLXZJ8R+/MmXIFhctgZGlAqF+gJ8SzX8gfhIG9kCh+
UUK7LHXff2zzwTJbrKWXNbrHy81y9B7TQEG6+X7QsPL7UQ0mEtnGAPlWrzpvruqqnwHq/QKNGkPv
D+yaUrWYo4K3+Yiceae6SoaAJRkSAOA6kCDaaIKXr1/YPhN9c7/RbrZt4vwkH1OEgsISv2Ie3xxD
de0caC6gfwVmpTSbRBPCONrcwTS1iVA4Oih8xfKak/91wEtBh+QMaLE2mMWKEsebG4muEl3nq2q2
yNPU8N+QlsnnGbKu4autgD5C2M/Z1MAJxoJ67FS9mB4hVkcX507KKomX+BQBYDRHTeG455PR+NY1
WQSuAaVuIClMOMOiB1nL+8PfldkZzq59J1980+ZTEtKOw3E+gbySdM6qwOlygleYpqQ/6tNHUejX
FE7lGI5w+JDXC7cJpOO96jr4DITeXXTgaLkBtlxYU/AoJUOHaTqONZT5+XCna7BRr2oOWmtB/d9O
2xVHBlx+cRBKVTHQ1YaHNeRvOvxVUFGqgcrSFv8giGJARdQqUjXnELUNWQJcfbEgJlfbC9Y57xJm
d5Yf8kdLnMHFPwXw+oUalbfUtiPTyQtKBEmOMkDcHoGDNz9G006I5mx47qhTbSLp6It3XgpvUpsA
RkCEwr/a7Q2iQaQKloVoAA7A+8+O3+YGw/sCs1iEYZKlI0aHaO4j45dYFCPAZQw/NDwmzPSDHBv2
fUY4vCCDuBMlT2rPNRlMmnFkTzRb/mSup0cQknKNTwMJTXv1k9TkhtWtOyUG09n4Ftb85pKBZEeS
kKDIiVJvy23aNA5jOiuzoPzpubn3g646s4QbQflR5pctt1u4EZngLGa0ENYWdvpbohcAde6VZy9v
1bc6H2pfmzHqw+fUH07/QMv0SUICUsHGHHR1WOE/7WraVcM6s1oIr4x46vyptkFiTYdAA/4bPCgk
qwTqMvo15MEBUfkf4dypjNPjtKYlsSh9SZ/G3s1y6Ck1M6FLFp8IOXri4TzUaJshXQ6ihd62Mkzb
KxDjJQFgUMh8cgDlpHhFfyvSvPEzi/k/YjmxcP/PGL8lVUAXjV8r4JD9XtUoaueji7cj5HkHDS8U
o5JXRUXgBmN6H/KNYJA4whPxEisNbd8XvQT8QnhYWNm3NZuiOi3CGIvmxxqjPOJCHzxcuQKkPcdF
qJsq+ponHONY1swUS2ga7d/f3TzCTPnNMgbPbWGY+LLSygMwQPiI6gcFOQJlOCcY1ocoaE4dwtQ7
GwSFocAeXcpyTkTvxpWCtSzRuHhP6E70/FzDXvS9uVb3ViCOl88ha2rK73Jtci7ETgR37xXs2wlz
JW9rUEjfqP9ZGG5jYO6La37UZB2XhtDjhbfNie4qMsGAg6oS4kJA4Yp8oSMnsLlRcXkzdWqKna/8
NVSRqUYn72M/96BALBulmx/R+KfGfiv9p2BIBP6r5i7/kqjV+ZZeCF+HgHr+ulJpXkb8L52GFrb/
fATE3Zqve+3t2+2dpS1RsMi8Wi17Frt5llmrYDd8GRUyJhCPrTdJdy3yHFnEx19ClucPcBoJlRCa
ipfbdxdkwVhgLnM0FI6Z44rEwdgpZ5qWqm3EM8/DB9aTecngbHw1xKoNdL6Zb0E5qdMg7BjpIsev
vPe9RZzsaSvogca97cLkK61WmnQUnnzBgvbnd4DpjDHAPuiFnOC10LHOOyqoBWi7NoymdlJPVWHm
ZrDa/JBaJoZsBfQSdpm7aXXyeqpdmV60PRYwTKVBKlorS7TNFJTbKGgwk9c0ssPSoZ8cvzbf533k
D/VKlWAjY3Y/SlU0y8z6Yc2DMUgVE3Cjkwuwo1YtY/fvKMD3qONr78MQlDX4fgBgfOXSlz2rNw3R
qJlLeTx5anwyQIUwyUfnUe4yG9/RJJSnjZJiN3pIdhL4e7h8UD0CycQfakE7ZnlYKbqUgVI+p+DO
HHzkUsiKFdED/TgP3CZ5gHRiHeQ8bceWiKLAhjmJY+EevMb7M/07IvirF6OLVx6e+Y3bf476GlHQ
EfxQDumvAwlLqSyfoBcNfuyEiimnMckBOzR+Ba4B+yp28CnUlPsJaRIU5hAG4tOZ5SXT6HRjtplr
nSiYPYNzzaH5hxyiyjn1WtxhK33wSNkHd0AncXORUmI1YlNOAPPCJY9CBDlMoK/den0cXpfYGBpN
4j7BCqSa4KEiPD2PbRMnqmNomrCbqMl1XzjLWLYEnRAXnksd7tJ9fS32niAeOdqFlumJQJiXIPGH
DTCFofjIMseu1/EwgabXQtJYpOpVVo8mYa7QWwZUuniyu0HpkegzyJkponp5pmNmqOPqrJlp47/x
0aJDMdbHndIs/Sv4rRKGr+yRb3Y3V+iKUGFkNuUTLtyoyUF7zCrAO6w5oG9EVzjVH3khK/SJqdt+
klc7heGK/Lgv5VtijYsvVmct4XwOhaG9C6qpF+gSBy2eAcJV4c3xyOgBi6iTn7CX4Ttcdv9reu3i
bWdl1/sUKw3lbK2BRsTNXmIiSfy+Nca0LGDbKJ4RDZNjEalN5RsF+DXPsFEgKGixyRbl07wihrc7
p9r9W2N67KHdZLYLhCUZapMXlvJF4JW7aw26XpKd4EHvQDotDbC+yprNppa3wKSo3OL7B+XlUbo6
ufKl91oyQH+w3pi9OMtWCMX9mn+5bx6ZUGlAPGNdgTXuQHldVyg5MpapBs+OTVVjUgXNCcunoIDb
bz78OJgXl1sGDLZheixRBS+SZEuFdr4FMas0hILVEh2VDV8tuExoWJ+YyKpggj/oUNeOplTg8kR3
aNUXNcouYY1QGTus3cReHJvVZhgRUc9ytVCSYkfh9u3y+E9PO6rR5OAhWe68m1wc3Kq+avcdlPjW
Ej3NYq+O3lnfhhVVgyI6WKvjURz9bSmUQTklPqPtYFkBfX2gZy4Tn1lUW1I6BdPEOQXOfKNN4msH
A6qjBbrqDyBQzZo2+zs3Bz+HhyntEe9O2Aw1PmrunvCQ0u4rjEb/0jBIRY913FJvUwpflWUCLJPK
4fkokbOlc+MjSmQbjnVcLU0/IwxRANKAaEpEsCm7JhWqn+TTOCfdDqpGjn6rWBL0IqA4cgoN9QH8
nehysCNgovFoajWDUfQoBQ3lledGLLoFmOyerJpIRfqOkwiyzEm9phk75jRpEparRKe3NrZaXyYV
Qiwtsk57tsaNdX8zgeHX+gBsjWtcNTDpX6/0WCOS4jUtx8DXKH7JM8V7L5xTZzkBq5tWPbErIy0U
HkMojg/iiZzWNt+K1IAuofGrnmgC5xIVDc9kycSW+NMBB+0YZXTVICtBggMvj5krL97iFTHc9Taq
z1kV1CJZcKswq+K7M+usyip7GBkg5iCqPkYIcLW1iB+4Zv642MofXnelY6QyEZ5o7casvvd9iYPi
MgseHbBrLFPxrOwiFzTuRlsL0ag3GQ8rNaaxqnQx9AZGXdX0x6GWxMF7AuAbfadxxi6Cb9ypLPBz
6OC4VxGRfTtfveanuRcZqgspRJawU9PMqHYsgRb0zn2+Ok5DngznmgJaf8vJKCmmLKf6DIo8viKn
jdg3Y9661FsL7d1z0kAeTOcKCdty8bu/c4VpU6lrKv2jBwZ1X9zoisLleLLxJ18KQ1ji4+DzD0vz
3nfjXG/orV1E2xnSFQ9P29PTtK9LltP4Shv2sukzpVyN2PUXmHsQGLAcS8rf8cyabu13dscjKXZu
uN523a6C5nAmnr+NkitA9ab0DgdRWKFMHOVlbD0m+L2oAhm8NrRZb4ZzuBQl7QKfJDUWtX/0c28l
yPbTjgg7nxPvveLrKb8p8lO1uL04RDKEjK4n0eMKYtDeFoNv5W7MDaKb3mr0SSlkDASl7Knng8RR
tKGVIGDtZwTgutzIpGznWzv7twBvP5DpSACOq3NsInKwbQUBCVPoXXL039v4CZDJ0F2E4RnuLJgj
JsHLJFAdknxVTV/wDJIusLiftyMfhe4gIdsxaiCTKcrb8BQdZLX0u07xDcbtatkresF+4QK1Y+XC
ABa8hvQgSBcWRgUNj1Mz0126C/uvjrV4y03uenKqVf/zXUYfJhiiKoU90spxChaxw3umo0AJPLLw
e0qJNMmAsX909OD7Ns2oJ54MQNaNcOd4C3n6SDDAbofNCLOJaH0L9SGVEbcEDCIWekn9KozmBcuK
jfgKQ6kSpJiRBJwOGFxP6XvoI1tTaDoVoX70waIeSqIYLM8eNWT1pjaJPlCl5sP25I3rxAsdoncf
+WWY5sUxrE9h3kraw5u+8p17GyN30UaxdV/41F/Xc0otRUkIhODOv4lPbjbHAHzx7duCX67aGLPT
wq001d8bJdx5VTuC6OIFhPheEDwvt56iU8gmho5yy/dhUBkA5h1jRe9JamABhOVxMJ5EzGQmfk8Q
aCHGxUHCAs1huEMp1N8dfpb27CPErtfjIZVB/QT+JwOoiVrzW5a8IFamrb9zXew/3IfNS5JWH2Jv
tK6y0BzQjurv3QtLGxC3dM0Gxa9T8HjVYev4j5r9+7vtLK9juNxKX+cES58ahz15FhfZ/baGWouG
DCrxqCoVkcOFQfeORsmM0qVP+eET0gsMNbkhL07zb0bToKqEE9LywOVO/Ac1sE3S51mZxjv2lQdL
vwTYT2XMc7YFgAgHpLj+4OWSD8qnDoAvVunxJL5Zgu44OfdQqW9Ox8n5Nt44tDnYdvD2a7Au9af9
jpS1x5oc6Iv1mvZWrL+o2bJ5TP22dVQbLsVRDfBg3jDyeCf2u5/2XqxHZDBmIXbPDKkx8F1mta95
pcA4lQSaGpsPgFOSO+R5z0ccUBHaBW2L/gG2OusZYdBwi6FJdjsSGVjp5ajD/NPqRylSB7M+/69r
EEGj3fcsOEaQlbQs5Fm62XTU7oRi/wZKSkjMqXlAJ6hY1M1itEcgAZ6XrLZezXgokfDRFIkJfle/
vrwk2+8MNJGpyckQ/vX1CHkv66mLRD44hZtYwVnDUwYlBoToW/BBMjm2lIhtd+c5RE0mZOArlJAr
zquUzyEDnZ3YkvxAP1dExLZQl+J1WkEfOc+iXRWMHOyYjWxQJ0wrF05KosnJDE3+vZdiRjSNH18D
skqix2z0bUscxF3FACQAtslG8A0Db/THUfOUN00Yb419gV0Q5WcUlSVJt+KmQeI3ZTS8vqIefyPL
5PhozY5fEJXrBSpJqHHTASbbVtefTgIDgNEmaMuFcMgroEIiV/PbQmKBY0wIk4pcHoLzaoZG6SP3
mB6RaaEhH4Ah4lUPfyX7GxyamzUtXzXPh3+68EM/eb/sp4leRnL1FC4+ZAdFAaDQM7Qiqv4FV1/t
oprUGq5lChZS/R3HSgLKF7Iarpkl9NliE+PtD3QFKd9RMClJ/6JZ1RiXc3YlXOPYH/0R3JHtaN1y
UNjf1lPGUf2N7VbBj2Nf6kD4CaGWDXUTCn6bpxP2w9MnB7KKnk81P9/Dhv9hwfuOp22DJm0lmA9U
2wePjo3QdZKwT+odJ8TuIdi9SQx+Z9fRRczI1fPhS2VLO6H8E5j7Wns7BPzS2vKsQUdtL76THhK6
ml7snbxLYXdVF/hjcqMscu0NAYYYAG05qK3gAIO1iNdBSmidoH6fZ95VZFnwdbNb9mkMfTQ2zpEb
5fJURabbf2I703gjhv9coA3hWqPtMrJoxzS4wN5T9uLCUo9aMkO1e+IMzaN/HwSJrl63zirqdKNA
Zc3lBwWVNES3KtwK6QqYwKdg4fbEa2uuj6ogQ8pMiGAlRb8BI11CMq5szPJ89jfWeVe8hwLLWPL8
TWBW1ZHT9r4Iyy9slYslbeaM216HCVrc46WJ2lNqxf8mMvNNaSqRr07PjhrQRLNv19VadLWfNYSG
JZimjJC7g/f9GpZ0v5hI13uKxfxyS0W0JAahDUaqwqplBgtF+fP/VJmUfxWIXfMhYLbbfcevNycQ
pQ3jmTy+Bx/PcYxxTMQsp7LfWjYnE9Tev7ch+L86h37dtD5lS9uPVTt/R5Zz6GuwngdLOxMb+lVg
CluxAjgJlTx2Q9U4yEOYf/fN7YfnClUtu4X5rLKGVSYbKJW3nGkTe55nY4mEwShpljbooYAOZasG
COjhSbQxRrLYPjv/gJLuyI2xcnsqjO7wsq+mP1pt9d/eRl/CK7cGKvg5NyWVwD10M2teNNaMWmMx
pz4d+nPnYF2iZaUQJxuXGYy3WnfSffId4QGObCxeJ2C+KeyKNja1ZR+honGbaaZXrmy57jbZnxdz
erV9jWMu/Bc2zhCVebkuifJA5nXO0HW+Hb8uZce/hhzmP8kEYLKYiC0tW8A+BhTeskzgYy1u7Js5
cZCQ49lEITiSfIja9ZuDIRQEnpt38wzy66/beBRziet5XednFhC4DfWlz/+KYhpQqo1KUiTQK8/9
a2w2nSWurQtvGQxOH8xE4FIKcXoSh+mw0xjRJfDp1j0/B4cqFdDcnczljBm7jqLDPMm8/hnkOkpe
SCrIzxzOBFligd3TS6C19zu+6Sex8T7Cmy4Doeci8Tc80op+EYu5MzNeqwTtCaam4ESLgZeo78Gj
gAOaytmuFXdOpBj16Id965Pb8iLeMHtuaCrsWYqLYJjTdWX68C1gI/aQRqHg0vMRQidr7RmhECjS
EC9/lJNxbG+tgPA+N43ooTTWg5h0m+pqo6msEPaW7AuzagTfCdpJOW5Nh6Zf0w8xKoSRmop+dkcY
msjDxuiHUPsuuKXGWjO/EeJVAiW/nY/TeiMP12OMO3CIgvlFCxbXBwswXLXGYf7oPxIAqgzCBlZz
+qJIJDZTcC4I0us90u8illGuyMLdGCIBEOltrsDm5LwfDorD8FlF+sFNqPX4Rvtvk/k6xl/18Ocp
qpL5lN15w1OlxNOxXXjhKt2d/iWzMf3wU5yMPgR6GoXlSarEgCXzTPdrMu4VA3xBrqGHhjh88lwn
aA/0WBLYiSQTKsH/PFOWMpWEo/1F7trqCuimZbze2pxBDr9ta2lKVlobaEpv/tH/cW36XmG/RnMW
YFtvp01EbRV2bHPqlPOYLYfAg1u4JPe+6nHfZTToE7kXdnVU0T7WupE4Xe/ayAdViyaz9rbBi2wG
9F9lB259ea3o5mGM2rSRVthMJU/VZSuTAN0/HolmvixjqKWbDN8+uFCu9JLeQIxakAlcSZSA87gB
o4SFIlbrBER04zpApB/Gv+Bq78DUvBhrYE3CEbLBgXbLTgNPiWsRWf1ITuSGp/aVSBDxkYDnYOoi
9H8wLZv0Z1SFdpFzcrFFyHva0JV5kWo5xAnRZ5L0CHCdmUMI8/lNRj0Qk4OzAMpfjUIurM+x/DRo
XwGtpJITpLwgXaTw/d0DESNmje9us2b5s8lQKRXuVtB0sggYh45SI1wXjiFQIkpUChjZDqFs9o3c
8qRRcIfojJS4c9bJzadXwvSaLK4DbqxXfuJWtrdJpASqUrb97XKnSYvU7mvRSrpV2IilhWkIckp2
AWYn5NyvWkCBSvryoKvvjhqxeZDc3jp2LddhOf3z9oARuKbthpUdRE2291PaAyKqPza4YFsrySic
WS1DKaPN8HphzpNqQuYUUKVuEA/pmjIcutw5K2e7LMrWyTI1mQaNfe7oBlCr7nNuPmbF4GEG2+Sh
+/8sczJaZ9heLHWCiwwR4Oa03B8l/m3g+YZoYCoFKovNAD3AM9RAEZgYx/rD1d+GMi9Gc/hgFU4Q
5Mnn4F1fYmOmCTi94pQcGr5132att2scT3cuRdDQ9dJJAEHPUrFVAHHEDx3Z8WF/9rlKwsdKrvRt
Jm7LJQcidSTEyT2UyxG80PotxL1TKeOhcyky6NCMz2vNNmRTfoKaehmMSs3d7KUTHp+ks+sm/ZsL
TQu87BntbRNtSrYiYfs+cFrpqKTzs8BMriBV6mqR+ntDEKH8BD94GmiDB0BYrZXz4cFm47R/Eti5
raaMdyfmqEvmCjprU67jnxR6rELJHjQKhGe8c3+3LDdl/Ztd1o1t8JagFISzZIfZfCFgSnNxFoFx
vi24Ta1xEQVRcuiCj5PnuwE9TyEJvaRR4ega2ytJ9tUlcIKUDPj4MzUTvy4y84pW7XeznwULUIpG
nVP0FyR1tOqqRO9QKY/yh4uuQ7twv6B8ydVbhhaVXCMNV94+2m4QE2BwvKqEUvxBtU9Ul2Y5Sy4A
EvSQq6qJfpwlTDZjaDoqgZyBnxXuFWxBEsBNyXyfmswJowuzvvR2+dzy9T1v/bRae60ofZUGUO2N
fDplmLX29NWhHDN5WzJy3l1yAsW2z/6NYeSKpGD+CWEChR/L0fWebik8OPhvH6k5KGdovVVpXvVc
MPIjx1I1Rs6d11Sggra0fXjACu2BNWH/552hyem8GWCQtM4YxKL5qCCvXYtjBgUEmsIhYCk4Aaft
5pfGzbuqPVKejqlOBapYI+/eYlrwx28AZIdD11EEk8qn0N0edRnssYpDmOmfrHerPfJF2IBMTEPB
SpP9N1W2EQPWaLlzHFrWj3No6/jFPdDxshsyVYHbFknI3YK6WjHOnJS4HpHl7MQb+EcHDbPq9c7O
PmLjvi7Xi7BHJd/V/m0EtswTVYEoz79R51mWZReRbhdp9gG/WyJ0ee3qDdp0aWxx6nv7Rgm67oUF
/DgJNRseF+h5VNpZ3ZVtbot19J8nsEEUnRJH4AVzRvEgYdq21Vkfd8X9kDUsw29KEc6h/AS2+H1T
XP+jsxkm1gdZ1zCUFemBJsvezyFNVVxwBxKAybFaLQeJC8LnwYWotvOUwlyIAceq+9+FjxZDOjj1
dc/Aojx/bmM6v6pa7TuYgeazZPctG0d1vaNenV83E9UoCPXmFtS+CZrepPFmViJrr3m4VxnvA9yQ
bTRR2EQv57ltXJbCbozT3Zl9X56XL6PnnSwmvNs5ylEZnCqXySYawEG3dAyIUTGjtyDDhO12mmBF
j0Tuf56vgBp+LexPJXNL27ft+ta4Cg79TD1xJ8aWycsgj/RUw3eZQGib3f2DriR7LVdfzQsiZRhn
7BNlNSSNNHZ2mQq0A2qwVLQ0R/aWlCsX2BjW/wKhExNGuORhdLljHtFB93wu0XcIr31JtS9HtbkN
BkrTtOXLeHwqA9cndO5lOyXmczUJMlqODC9zzq7dMXR6FQBgLVtzvBxJ7kktyJFASY/+AeBfSB3o
G+s0ZLcwcIDF6nZWh5Bm6jDR18iQso5b07fhfCYw7hCy3/NOZe6sVcXalmtUgFToH1OFY0hllH1Q
Nso4rBLxY8Tj2X+CCbV5vZ/ewazENU3xdt2lhE4sTf9r2XIPoF1HsQLZzBhpcvX5c0kzmoZeDa+B
HsibmAskj1wqbUP4cQqSrZis6Ujgagn7uRTrxCMymbISqYLDLTECfVPf2rhTCSCG7pOhYhq0MhyS
+Oot1SHdpkIQxWaWfD3Q0szGphzE7RG4c2cmVig5RRiMbCxPE3c/P32X09KlMrwje6iZ3QCHICJo
CKoUD7esGAJA+RYd+x0v0wU58Szg3h7fh0kxUBD1fKCioD5yxNKoXuDLx31iR4qULLqlnLu6S2Pf
zFJQA/2rqPCqxZ7aHexB8S88lod8Yd+z58ve8ampfmC6AHr8/v+jee15dzNVyXM5/BHDMaQxNCb0
WRSD9lobe5ivWM19zF2njCe3FsFQmm0PTi/8gvsYThJqRs0XenHD34sVqma3F+Me7sOoMu1yQn+R
Vf8omPAh9BUt4wZPCI6J3xdzxMdLYIEqkun87ClBxUUEzSwcy3EY+R4igrJQDV+6S7ZuvBbzTz+u
I3XTfWyRIqKSYd94Vsqa7fvIOdwlEuNC7i+hWlRXevQb/HYEccnqFFwQkFNyHjLlPjK14gCdT2po
ImnNluZ1xSkKWLTaBADGd2vJ1VzETqsjnUDKk6oSucm6ToAS5PpA8lvZrSTf0Ci8B5/4TVXrNnXl
amxcUgljNeZDMmAsyft6YxtQmxJRMrjmz9QYazV71AZot136i5/aBIZuYDXl+W2mXOw+LVQrapX9
gnnXXWfBcveB0ziFqwV2QrMkcxWwsK23BQGRlN5/RF++ItOZiPP9CNRNfXBA7SigmOkO0z8LbmEZ
/aM28RODDv124+XuTRzbtvHubBjacE7O1qXtBXfKYbVH38wOxHJJmaZvFl3w93El2A1t/WVbQWji
94EL7f2fOHnXCdE4zXAA12SbnjBR15pVXEjfKdSaxKuikLjgHXM6zL0RwhPbhbS13HR1VZ/h5qi0
5bKfBp12A0KYy3Qh9QRrfyj3ecm0VBfaaphdxRdpUzQJ0/pLGKXVkaoIO48JpnASOoovHxn1BZbp
KFzQRKjWp0dKMk7Ia1rKUihxBdRFAJ6XD5Aw8b/wyPbyqPIO3neV7MaJ19YDsRM+XJy/EYzzhS1o
C1gnXC2ubBADqjGgutoKzHMq+3NI1xTHDJpBHFYkKkZYNRhkd/LKcRNzkyt6mTtGEwwhYjywo6gy
9AX2Ncioz3NDU1Fs3T+AUck7mjx2Bk+lKnCuMkhAUUJZu5pj8l2txlUs06zJmzwHcn4WLHOoID/r
bYakPTdCBEzMuzyRgoyLnmpD1FTPvWzufIjc69sZpQil+8UBHTdhfkWiLxJfpf9F5EbsrrE0CNB0
ohrKjR0pJ7uOENY9c3grWg9Rf3rdIRmF9xHCo+vxbMmjc0CExO4wMNmi3NcAO2BFJMjXFSMDNqU7
Egijd5JOyL9zeOYToyKXSeERcBW1izWxSbAW2Co43vD1aRMLEeipfJ7iUuhcGF/bcIFVwfczlzjh
bo4RS1EEheytsyh5RDfIroUkNyR8AZ4K06XEqeGfN/stFdXdMUiDMK30aJoJwb/hvXlMh6WpvXIw
1ynsqmN3vabDc4P31rZRTix85VnKYgJAAaej390g3MdVQ2zpMqkxkLASSA9qcPi3mfVFE2r/xmEQ
cdJM0TRATQGhnbGx2CbZ+hWX4jQQgn/NJT0TMNHuDK3IP5iH6P6y0NWBP8533hs70sCP2wUU09Pe
8sgTpRgS/DeigIr6xWlK4Qoh0pWxFTG57MfBRSTIeNN4ylaNklMynmnhSbSbbTrVbR8YuyY6Veg3
o0zbZTre4NKm9yPRTrkgep8R9ZJtRUS1s7PL4e5MIV1V6SGdrb1c/eUAu1p9AclQidFn7J5Yy+sF
cA2J9K2lipJoVG2T0NvtJyX1iRvX13daHy3L4G0JcBh2yzWvx6qdP61AHUgvwL2PMs8SzFYlCwHW
GLchVvymCPa9VZRAUAwMYKcyzDcKJdf5diY1FUJwqM7NgoSA89ODsPgM8csLcvDMX/OaOZ7gR97l
9y9FIzUq8598hOcCuInHUiuwFLKwjo9LScJ9KskQDVvUyP5QTqOw8aUWgcmXFfFWV2JoSNqktktf
vU3cvCHh2dGDemg5OmCZ162g1oiGWbtMAA17qnK+vsIlZr3S4YInp7aVhRVyFfKsIo2vugn3Bd8C
sdh4XraBnrj2XwmiSGNBsVbmBL+tK+RQ/fanIgZcyOJG/7AqHl03GSZ4MQZsE95jxrix3Ea389SS
KrTmRqVjWlHYkzhkpW9DCph+aAY/1AkbVw8Jay8+yTJqz9Z9g6Otdm8IJDNCMCUcY3Cm5TmKt7Wh
0o5x2xXKA3rrtKi77m2alAnNry0tB7TsiMLRKrJsjkR4TjtwMfBT2N7vfRM3hNMX52Eb/Ftu1ihY
dFmZQOmcRo3AeIKX6/4MISyOGl9iTw9/iAiTqt9uG/kDTGe2YGwRZ9GmdNep8ypKi98UycvPLkuR
itiT87G9sCKgTWztasiHVhD3o2kyf1ViNDZ3QKx6tx2Tzv8f9T8Y+DPTIZX6v4qnzh71Ywz7FmZA
63zrtlxIBxRXqY7zAQVKiIOre7+rErLbtEUzJwahQ4U7D/A9qc7i/bwqVzkPOi4ezpZ2tlKCKTu2
C7677Hq1rRh1kmQNd9yG6hvV/N6loXOjU5qvEq2pGtEXi5QM3LqFk+PoYyIEkojgqWp7Of25QM7G
+dqGcixT1iwz1u9ekZKa2XCQLO/gfFZayaBl93nJcw47zzLOJq3BEy4fHW5beoaUp46ZEnUxyVan
n541rAUz9nJLdfBqIDlJcEBX+AQxeqvSXT5sLoulyNWqGQerQLXwM0F+HPgmbDKoKVjfxQmeqhXp
bt1EGvTQhUjYlDI7FQhOXU/5o/dKgnOIvxNRwhrcX5KaEi852cZ0RVLFZoinXBSJKs8fZxSweGzo
0t8z1Tmhj8g2CC02TwN08N5YSDSncfTWLp1ozfJD7bbYLPFTjpv0tG+edwtwUVJO7F26j72HuuNy
Q7xxlXTdx0F6a6fW8nRDl2PPCXdf6Fxf97CmnBTeO/8ZM1EMENvF3MA9mH+JNxMAeeFOlSTEgjnn
oDQs5hZxY763REj8d80wclWvrGEozEbmyTGhYJs7pKHogPn+2w/Bf2/H2ni0MWmhP3gPm5eotNpR
anwKxeFrrZ+M6NETKM1JKX7yN/kdvzyYmNz7Tbf34AYxgBt9NfcWnkEW/3v3GIJea+/7forrj8e0
fBhuBSXVaUwKsS+2WWm4hlvJMJbsfbwMFJUaj6iWyAf1qs3kS0UbCo5myWorliIDxIGyM6ZxGVui
WppZDa8O5mEY/SJyR6HsWEGWjXrr6HHX18DY3h37AhBhJKCSFyvdxsEBiYI8dTfwBkvtEiEVyy1b
/EhBkOGUxZcD61Wss8OyOXhJZEwkOrWhHE9apdmGeJCphmUf37EYQrzhe0SzgnV292RspV2v6BMH
Jyx9WApDcY1hJOU2sQ4b/WWv+ZQ+EyFmk4le9Dtv8E5GmaOpULksVsaafd0JtvXXjVgIhpzuqcgM
o53IEMPFsbNJlmWHEj1/kKtZ2e0bd5/HEc47vx+KW0tUj/3nSEd3zPhGcfgpPWy4LtqsaepObD22
95SgWTyCW8cNggsAbTQw3UcntdSfsEZ8XSexCUmpSWch6Ch+WpmekM4etJWPHxyMTCJxGtV+8UmC
emUwoJNj5kz9fnHwa83tHDZsNf3ZDMoEhge2FzcQLjiMnmHHvL6XR7YIbAAAeq98WE4wo7J89baL
IQbfSAsrktPJktaTFZT2YCXDcpAlb5jCpO6uB6iPCywqYYO8nRSetQQsdnFQ5xZjVFx78NwGnV+u
v6gAhnn7AEKUY+dhRFOx86SsTuipC9jEK+Z2/Vyhi3U9jtumslduoZPkcIHwCYbyiVxgKfKnVaKJ
7f0GGsoTNd7UNlMFoe0EBKzp35duAh4THViX6FIaXTWmugXyzc4Vcu575YS/Fno7NBN7HaPaEXY3
NqWb4KV7wQt5T7pC5a+gWgToNhiYGdxut31wuqdVK2wnSr0m9VP7I6IdoZ/GPsZ2Mau7i8c0yISz
Nnxm2IudAjW3v1TTZb1bIPaiKaLOdDSn5D1YHXmCsOBwVQ10XwWtcXTYF9qk8rKGMS127GEUDzYu
sDRan04fxIrS05rc+1t6gBwLn0Lp851krl3d7OTcrZ4OeacnTU2iYqETUsA9Oy2xXlbRF9XHiWC5
CFjvIoqdVIj7MHHN66JCagMtq2AQfiMBT5q9J+F8GHiDmmqevcSGk2ROBY8fev5n05ByGY0At6zP
auTK+SgbEaxaZ41PxnarSZytsOtquHyeK3U97XElp4b3spn/BDvIRub6KGNZjn/ki/Kln2v3TjfC
B6440xUf7tV3UMWHFYSjiojNbdmtE7CRB6NuFFXhw6P0FW/3CNQaMceD+kZDPKSjyEyDYOv9+ZrV
9TkB1G/h8Vfb4RUDueh5Kl2AmPz7g4oHxomg5SGkansaz7xp1WD7McceqNPNEfBe16//xutHUk5h
bxc1VWEhjsHuTuLZc80TwGA/A+Uf7EWC2h3T2N1dX1QIME4+vBdLsuJi8PhSs0kPR4/PYVqUvcDB
fSfdRHbFLg7PsOpB5WrMU6rUnSosM2FSBdU0PSwNSvm/wY3uWzNYIXfI+pui1gRLCbYlXdrhfRH1
CgD5iy5eP/+YegBleiPqXshriMh8m6wSR36ps9Xig/XvUQsswSF0GDX1IHCDf46yNqu2PpSLZFCP
67NXBB7B5KXCvNKtjTxV55EpJWWudZgQ9q1rFhGDLdmNExKJWfDCJneIqn0jPurzpPSTY1j7FN7y
oo5b4YfuHguilxFKfzNZwPPNCq39vnm9TUtRw1imavBGELYhzkP4jku3G3YqOwXWM3xDgv+Dgpxz
dmfjY+0zR73ZXS+J+TeJ0Yyf5UKkCbApzhZOhLgpZjdbRi7KpbeAgrid9DA7PgX470pL5Jj2UC2j
90wvGACtO8woH1ReAlBbLH9xap+fz8rallLnUyF8/8BI5Cw5RBEa4Ni+7f0NkJXqK09+4KydDU3s
7DK3GFD1biYe8kniorNk0a4Uuyz2ejKachMQJevutnrFAX6CA/MHdd/gDg+jTOJXqPU8Lzwt7KX0
ZEImAVovvrg7jqpCtn5LN6qU61aP2+fhQJIoO594QDU/K2y4ULhh3x37ExRP1EQjt3tpb1RgBgg1
C09iS3DKQnQqDG2Ph1xlZ3G1ZzyHSuPCdvTR+Haq+aAlx4er0zyKBi1n7A83lX20BOBrCFHTeUkL
BLkp97OwdNiZUVkIPXZguKAtFinhpvLOTWfoh0BmK+UDrWfZI4k0isKBnWnN/qkZj46/F2GvCT7Q
O08BaU363pKNH8WF9udLD8dGq/EanETPfdqv75qy37e3Y20pdzwGownJbXsDT1pbLB9WOGC5ifGw
hUInIYCDfCQaOChBenmdTdW+V331ZlUHgeyCdJQko4XhFjNDrlOfChtRQD5L0GN2Ue+rbQ/UUuYQ
ZJ8YdLPZRCZvEVRQENkY0b53VCULQljpI28BI5WIHtaBavb9cOuks4nLematH/b+9v6obU9EhEkR
PP85idXsLgFOI4F8G/ojHtHgW8kwUcc2t6a0KcTpKjzNlsvj7AgyK+X4l8Qikmi812L45Xmr17yz
vz/Demd/9RaSR/Jis3G72wUO2YN6BejKgHSeqNBcpigSUc84vRgn3ZWnLIZiGK6H7brIHpluluYB
+Qo9sB2VO2C1y1pUmeSwkxIQ1RLf/3P9be941QOd2c5NdbM8HO5GpA2Xg1KRKK8lF6IK1mbj30X1
g0Rwa3/3tEOK0zwb73k71Vmm1nHerly5KWHKvLApVgOXBetpzDrxYyAAue8hUVhXECNW9m8Skw79
DUeIhPuqXaV7unEZe/WKLZHWDrHJqWP5Dfs7ISxr6YMZZ4z1O+Fbe104ISI3sCd8pyiUZg27RmpT
IthxXYTDNdri7dVVwHbC6GivfGIeF3v8Om2QwB09+oIxJ5ZcI+80l+oFGmOUaW6qRjgcQwl+HbKJ
z/NKMioI6JkPfFqo+QOZBFu1fpTIxunOvISyMShvscFm5yLFy05+7XyvCUqS29FFbVOyVDvIPufa
w2NdebCeJYp3IxbnMO72TZYE8tO7kVwXGMUe2TpMwGcUwSpZlup0s4knUWeOBCARr1DPHvAIMME6
g8dRnVST9tIS+L7fxsImEwjPzseisV2V596yMtI5QGjOn/z7Hm7ChJn6L/LtrqM//4DYFf3HGfrA
SPggkbfS2uA4BJiFUMGqzkza3DCE2gwAJJpRXOSf7jZYK1WRbYm1B9HRLwRX3EbDGP8glDY+USoD
iNAYw3zN5zgplx4EQuqZXJLYy3arcTDAQIE4QUTM+40Jhlu/v6ypdrgvMEabl6L2HpbIr97KQCgH
RGq5lWI7bXLtQCqJ/G6g/3OE5XSEvlhfN2omTpTPxFCf9ILv6PiFS7Ek+TUxP1iCBBKnD354vNcA
jgwx2eXiSDWHdFuJdsqXmj7D6ui6UsWEbUHqiSKdz2znfPXTAdveCrNmBCttyzK6m0f/s4zC/yUw
bIoo/283qnCraSS8KXNHWWRZpa8Jg8E9eKfuE+OH91yxaBvHSrY6SeJeYABmnjInlPL6prkfF/jT
WbyKs/kbq0m+4pT7QLJC7gwfH1F4d3CXS5a8dfKDY3MFh1spEqEcJT6mQTOmkMoe/J3nMLT5cLf9
PsC9A7wB6mEes+/FFOEKEW4apUXAfXPkajjCwTQ6YxqAyDS4QMMA3vKBLUTuHEGCiFs/ggR3YUvB
rTfdnnyB0m4sEFFIdCF3DKQxAl4FaIcBGPB0AzfSvfA57rmo8wf0aSGSlPAOdNLzYYYQpX1KGnzv
y4avFdWS0wEMHU7bVPW1fTPA/oHzSFm+b87kuyibqGeCToEO9bFG7tlk2cG0zIrKl9rkTmReHcbX
OmVbR2RZfGrpk8AOhfYcQ2v2inqSgicxAZ5rXbtVazLzOYfr/DEmyuYuXGHzvNxHEh9xJ7yUu0a0
fR6ygknlpvgXGK0Y0whxE08TUBp/H7TYVPzEasWqrPsf0MgYNPidpnzige9gzy931Iq3sk0l0tje
SjyU+WQFh61FsftJkIYK7aZQasPlhRwGCD6uuMr6eXPADsiauAGRHngHnTQvPfqlkv2WxPatXCo4
AHmKiF/836kGzd1MY9COif/fMxwi+7fg+vX1KCEDgyC7mnnvMZboMR8KnhLoqmGu9IkLMr+sQwKO
OaGQVqsXaDiA7BWo/UtHe0GkRJLMjEUxnnMwS8Xu+4qSBEOCLU9+yAwtrcUhaP4KqzKxM30Omr8l
2fGdqoSckFuQ6q1IZEtO8TXo6f1EOkqEM/sw8hjEZn0dzDJIgfwAIeQwKx/segTD+mZ15VUQYwE1
fnrIRHWMQOiLormzuWdgoIy0hpvKj7sV9F1HjfFnNkY1Pxb/Qow8KuYbVFZ+Rd845pp5fPooDBFX
u9I9AednTMZZoz1qWSImbUimaBqXkES4vF1lHiShjBd36Kn29WBQlO1ZOvptRe2Vt0rc1j5zHZ6Z
3heV2xV9UrGufFeGlGP/yOSrN7h4VGJ3kdCcqLJgGCUiEk77gTYkbt/yvw+cOoZiLrgNCD/HO8Qw
WPZ9qFR8/4DYzWRapP+8Dt/x0JUM0X2Gwq9mK9I+Re+r+YC/jvW3/j9vMD5TyCKXpuAUBlPeMvAU
5Swtls/hsiObJzGIxylVLM1uQ9OyQJcAuTd2gjPbZWznRk/8nMEIQcA8s/lk3v4n01YSWvSLSbgi
38jsATQ4HG576f5JRacDDkgY98TiAInpPKVJJdpYUbYaEzwi8/qEKUyoqwliC0COWWnrcn5pdyA7
xAZkUJ7lE7678B/BsiGYpEoM8mBdBJWk2CMZuRIbvePudHMHPORwDMy4ct4ZJIL6x5+AkJHxeFgQ
RcMzrWAHxI/4BA2BCrcG3jFskIl/AWEsDSGs5YJ28/rtv8/1QMu1h+gk7tWTw3n/hz8rUILeJRfi
z9E94wa3oCQLkXq09AM3pHSpMe6qIeF9sc89IFu+D4TKrAM74yHVK7FAMl3KsSg/SUwJzCzoyH+z
oSUXMaIDkwmDMeg8RYucMWgMUs6aXUU5bkrT+hnqcklI1W/FL+hoMkbBuqjThCmbkkSWWoCTF2s1
mGryU3qVz1wzv+IroIJPtfRPowM/Z6ml7j1+V76tJsDj6OSmh22UuO+kg+HcoKXFlYbCcGJCFtDv
rw/xUYWvYYSddG6/x2L0Nx+LLFa6LqINm5prSD+lp27aNxIrNBs4tz3VwTgruBcX3CZOKslHCYnj
zVZ5nnLvb1gIy7sgbrFmnm79LuaTrA7FYVE7/ThdHJLlApcaD435hoQ2l7qSYxEqf/xfnC3Sc6rc
NdWlcxtAjAjyxSaKK5/RLazDmnCILijBd7bNj1jPQffiNOjBR6MMn/PC8uffifR5geirJIm4Ujy/
CgGFcFnSkNurJY2F1Jnkh0LJKvgn7cfAkzLUiN7KOfosFLAfcWiQJf4cJ+pAKcQmuTCsI/w0hi1M
0Ldr1rSJ5G+C3YP4j2vcd5HwkaJQIIJwloMklOoBnEpfChnwg5UjiGponEjYk12NYtRJ2boDwJKL
tcnxbgymgyAYXzDvVJ9Rzf1r1cRj1tPTf7tX5sqq73cKFxKfehZPZOM6gh8SAYPTk6eGKDmCqsUX
tSYzJ6DJSnrHMQnF7JDLSccR8cHor2JE6QGjvojyq13v2ZlEq5guMAXZQb5E9MuNb7ONw50mQjTq
vHiFkJhhunFUGd+vcZp2oASFqhkChJDz7e3ff3cHljrGCxlh1bI6z5RTUx1btowr6tn5+O7YbeNY
Yc1+SiljwSBgS9HfCLmwehPomZVW9yhB0wComcJJz//Pjz3F0w8blCVW3DD+YRqHpkX5VKFwPrc9
JkQrqhMlwYcg5G7xKtJedR2WYFpQD9zRdq9Xuls7UXLB5HDXDz8UY/SbbO6iHtHxdFbhm2R5d5Ch
a5quDyDbP15Kq3FkCNFnlVo5EV4zXsyWOJELefETrb8tKvQSlY5IWAFhsnagpSrlt91YvdkKK5yf
ze/i06t+mgjc2uh1C26EhzVZ4mEztQxT05q3k3jJYXjbeyMTDDMTndYaAo/VWJpk9V9ZMT2KgypU
CNTDJSg1jn2CVPnpC7k3WtAuwWLSqRTu5UOkZdHQgUA+d0fq+a5CmYDyLUxTr3egGuUwQFop0SD8
FhsNtLR7L5cAYIr5gQnyq13vStpRhICArrfLpwyxJjacDVfM5fhn09fS4g2HBz3bc0WuhThtTEkS
iCEXFOM7yxEkXl4PqXMQjTJqsS4hYllUn8LyPp4ClguQuhLTugHLTUUEFvY6Y6655WMwd4fibR9Y
JRDzncgOdpNCpakx39QH+BJTXOCs/XgSRlyOwlLCY+1Q8Ds0UGGXfJ0Qen/8SgHg8gYXvRf70y0C
tg03v+085MIr4wosbjpRkTQvR06B6nJG9CsSh+TVm+Kp+YRYmU31sbkM6Aov24dVdhwBIqoH3A76
Yt+x++vergDqxxv6vHh3EdpDPVbVb2VZrSX00nTcSBHXxCFIo4sJEfVr2ZkXokwkH8tdDwz5Sdn6
kaXDmpqY5fbx4EUefE1wuwkU0oqCSWOPmV+Vry5x796sy8MgkTtVWC9FA58IfEir8W+DgzCqh3ah
UcqNu8Lr1ayxh+TbK30TmR9qwM2Ja4VB7LqpQWA2pWZU1ewBfjsC5n2rkC7diXJsVyGQttCQ6Mo3
UjPEnUs44orsTyKK77gBNs3quO6E4Fmh0cf3LfsL0LXy3kFcLu+k+ahgAQyrH0OvcOQuG0xarx+2
a3uDhk1NCX6v4/YK8EaKOTx+aYhFWw2pND4UEKhxNq9n2X5MMeUQJdy91R5+xOQCsB65KLiTqYlb
b1zk3YH8O07MjKI62b4kV/qF4zt3KMH6iVFchnULw0yKXVV/4fnBA9DThgSUegeblo7PeFonXTMl
/v0pJa19j8jomGyq/WALTSOmEluu24pNY8vW2aL/Pdk4lp+S14xO/6nVddLHI0SQDD9C46XyIjh9
WZusjd5c5IfYSGe9JX3+98QfAvgIszKNdED3xhQbrW+AwYDOmUKezYXOvHNxDXa8df2UJH/O8Y1K
L6WSTuMX89Pp5RH1Cty4k2zwWsVYWd3fLmJbCbis3t3uTDK8PwY4LsYEoHe9HJrA19PW6owc7VPP
gS5jM40tiasOoa8APcpsF4mn0OyAW7OZ+vVtuFYgxmOyqnghSy8MUA9fFf1/cXGlOJfS6defOx55
hcqIW33ebhJ0m82Z6MATBwzrwn1XIuKZYtV20DxK90JjQsnR+0dYP37Us5MN7OUhoBNaIrocLSnu
M7ID9GxGrw6UOxgUsB80Rk3QK+2LkrA8pJMc66E3P5ovga6VyE3Q0J/ZoXl1c7rDw+bRCq5bjhge
uXdreBObp6dYib9pvBrDyLlM4QJDdOAb36CtL+0juE1UGF0p8O4BddvXznUX31qtdAl36VNAmZzX
LDZQdMREJ5OqiW4MaB68RBeaxvyopIjUlsC5HGkZgJdHQDj90v4u6SdvQRZD0SKHcVrU7ii5lXqm
ixeYT07uqhnDsPG/OpRi5jmvBwoR13PXpqtEQVGcyScmw3g6PFc9cFMGeFj9JLOhzfUiq3+C8n5V
kDvIrpgk1k39t9BI2SeM3u3eJtDX3qqmsZsGkt2vbmOXvKFDGJiDg45pVVNXVwscy9Pcl9IPGLRQ
fmsJXwioPx6/t18t7Y1IUNMoFgMhC5PphYOxRihVZBmv+lLJ5HRmZYFgNfO7yy+Ub8P6emknSCqg
la0Z0dbGbMFK4qyAx93psdvrcDL0qoPwQQYgzLeMzyAmMaepnpBFcwoNc/GHlvlzQdk9nBowC+0l
5+SGKdKjKayFAXgVC7rRCaJBADty3nQ2QfvYfALOSjIxN3CaJxgQg90AT0f1+o1i4oa+4wAxk+d8
5bZFDlExZ2HUJnZjbm16cswFh2oLvKYtgi7x8RqHKGb85XVm7r6As35CEcMCLwrNkXdq1n2D5TTk
lOPRvuX/EqxQTg3kLyJMT0XBN/Fx1kuqWwlXrdVSqhiItXKj7FerW//HZb/Ucpg9PDFq6g+DZx+W
hvy99aMsFpm0gIPlljWOFF5+aoTk6JHzOY2OpbF9SR2mlbH/teKjL39mRFKnmWjUmRERoziYE+by
JQFwYEKnqaI6HlBwDmQOEIOffUDfxyE+4t5QTPHo0QYRGELhDHkXisRQtWicOFZ7BiWC3Mo2Acjs
vNd95LfDmklNY9YUgbSWMXXN0sz0F1hY6YOv7/3vXcjQIyzjY8NBSQkbiLg0oRW9lkwCQRp3lJg2
WgIHHuiE+tM5e0W/xKXipAZml/MXBI4S9T/NC7tFnP2xYkPhAOMCckSwFSXeueq5j8u8Ey818ZKY
DqoqvjZ3C0xxYThO0AZcA+ca1Xgp0hZeUc3xqeDfoYxXX5KwTce09iVLBeptoZGlYw7JbomcFkB6
qriGWckQs7p1PlVUSta55/BeUD9+f72AtXNIbdMzuNxo9PvuXQwRzlfzOahW9tOuISXB6kk6hOcU
NAgIi1k3F9gMCWJEPDzDNuaOBhhAR3LQWlKvt1BgXNwkRHdHrqpKjfjgRCejgxLqir1XY8kZwpGz
IoAC8RLP6fKYieZrfL0Fj1z+LPeStrLlKtg7rMUbd3M0piRagPNDNeug4mdWdBw6lH4vwG7eXY8Z
7jBILPCfJ9Xbn41YbYmGV24+Ya5VHosC6mDn6b5oT2AWA2SyXtVsFwKsHAb3eJYnPfRohtxB6LQO
QdRpuMHIq2dxPqNA1pd8sZwuK+c2PBestYHyqbkLBuxWMEXTmwIPLVe2MXEATBRLMMnSHXpz25mT
sJFizNnAVOqr/HNVIN1m+VOI3W89ULMea0ulFcnAgo1TCTS0+3gdlq4JgjSzZ3l+Szp03M0XEpMh
T3FHwXd5yueUaMIjqBiznRfCXCue6gO9p89ds+ctnS02u3oXcq/6bZqXLUXFEXfUWJuYIkZwUHdO
BDcKxMyhkR3q6X+15xpgKLL2SqEbHpkGOBzDKgdffxJN987e9qnz5FM683Iad/16CZCzT3RXm9ld
g78onyTM/qYZDq8Mxb8yKMB4tQfSobFpziepeLW9aJGsymBrx7ayp2vcG/+7bDpaMr4WdN0akRG2
iLzp8o5430wUME8dJ8FF6KY33sc/a2x1qBItAzlmyd/7dPJn3n6RgmtlefrQTCiremGig9oGRVGc
qhOMucnbXHs6piln6HpbzEepyUoiGiGd1Ve/jyVyWmZriGy6w4BZrFZeUdPlP/0THQ4xZEJdW2xN
4GdeQ8dHl+fxykDue3ltdwJNNxxEFolfMJM6FznnDcC6FkLrGqTMuA9RMidscgDt046zil1usrOa
GyScP2BixzZD3Zsx75mgliMChJDCniRS9AkXVsAcS+rpCA2hYFbt48a00xceVW7pAuJo7OkSpiWP
QpCX5WOTwTBMZse1veTVZag9dOzVLscFnk6s6a0K3u6s+cT66J86yayRHs4mLBFVoLcrl78odGiY
GnDnWZlkhPjTzFHloi5Uv9Grdzx4xlFvkX6xCidb4tn428Zon4m/rB7FA8rhTym6/boYxW0153qh
p61baihS4p8HmeIcdVp96o1x4EOcoB2Rap3geMfzngwXNk1DKTHlw9Vfw094OoJ8IbfGm0Xfm2/1
ngoeDWS+CIr262awwHx2TIaiXo2CM/3UmAiqHYtAA/Ceb9cO+9ilfsRmx/V9xw8ji33G51iEI9Wl
Ei6BmO9xtJ0taA3KZjYy9ZQH32WlrwB1MQ8+QXXzdZKYAf4SsoIJUw2FfiBlBGzAS1hSGQcDN+Mn
UcNnHpxBbjOzPCfy8+pi+F+oLSCQxxN5VriFv3On/jfrKHkKrawgWCsW5y5mjFKNiADNBgfD2Sit
t8jwropev+3VNQhVOM8yoD+AiuHMvj6CdZ/y0T4UW++HE7Czx1WVrAnHI/Q6cGb5KdoiITFNf1vl
T/yCN1wxrHX0s2JTwRUh/YUxldxjAJhz5+IQeFCfHd4y27imHLjuCDWhVM9eQ1Ma5V0Geya6U4C3
ZIA26TkZwDEuVGiZHppvJT5k59Xev5frK12waBdNFjzMSyQVWazAow/5PU1IDvDg7XkXi+IjHpUc
yqvjjTkxfICj2T09oOk9b3K78kpWhdNJLzd9DFl4MSXs6uBQKyX/MQXNV0KII0/arPzkysWSzwz3
AjClOUu2eMO6z+GVT7vWiwGGZgVkQlj/964SGWCXSpigFjTV41jEBGQ8VAOGvl/mlQ73j6yecme/
yQChJafy7wrE1GAiwmimychFDj9Bs3GQfrop4M8/3dk3SROP4KD+OcJYY+xuL5WrebxSt/bcAvLp
/qxJxHvzB9zGmQ4lb94dCnCIOKguCvGKG9PupdiGOLfFEtCK0CqzbBxFYpyBqRhRrVYNSginKkXU
PyFzVroGP1AbDBgs+5hqre7TN+ZKfQ1eiS2I27/V27aTdIKOxQDvhZ/wrR16t6NI2/lDd1oiUMw4
BAeKjbGeWzMmEASy8t7MD/HPZWFzuD+Q1zsG9Q9heVkXeiOPgaDh+d6Xd5E7uzaqO6m7FAdEDcgd
LNHThqIHJp+unuMGzflUYR5rA+xp5t5eN++HtxpB48S02rbt3c2TmvBVOJ6tcDoX4CB0c5ehQWhP
aGGxF+xGcDqC+q7WTtfLKWmzIl0jPLaUsXub2WbXimduFSzD1SJ5sfECGIAtE2eVhKjjtRgKWjA4
u2FuOBjZ3cptIe3AwBIIIqCl65r2UrreDc9+rRfbIhRWBK6RGSHrrpEBPUiTOH/EZFga8LOhnl3F
HgOfNssFaaKh6ueWd1orfmEhlU/6tU3mYR1MlGMeIzQ3ylwjsv9JzfRermBAIGzXCwyblPnplaeB
eiQZ/mi0oMgn+bo41iEckY63VUKcZ/w7zG6HTxAZ/zvG0G8oUttZdQTEMT4INGYY8fzBoYWwLhsp
8YPuPi5YZPxR/9Lp/fXSgSGjS3kOjlIbvsCwi4a+MFli1m4a2EZMzfM4GcZGl00X4ZIEEjPe/Dhp
52bA1+iLVv67+YnljN7+zIq/b87rvv0CGtlrfKoY5hPWGqZcNt7LONzcCs6qd+OFm71ohxMzCe38
quO+EdAl1cs3QixafsH5yCkKWfVkBXzoVz8knYnZpC5hQ34jCbqa+mrQCctv9S8e7MM9iFxigBkT
shq31jB10OSiPxGtIIXIhe01kpwVnRZlORluZM+Ijp5T1h+GlKmIXwOGJjX9fNHvbfbiqf2Zqe3D
xTvFbbn4nBOScR/l6nps4EOY3dYd1cBgiH+oxEyPQJ4TtT1Wa68q80X32VlTwn0/qpGBJARS5h7K
impI/2/MbvSz5NvnkjrXnS5vnDrlxSDj/fucPOK/KNZjRUMVi1PxeoVkjJvl7CqkAjXqRZS/Kohs
v7r+4Y63+UDHhHZk4takS2u62TUcLDsQo6OeOPgdBL1wugRmrEHSqYvj3U4IfyWjCAel/IyS3NVb
ZHURsTxGItaNmbsCkP6wzpLXvrYxWzw1Yoo7gRfuTJXWyeOvtei7JJ64lZoV0VN2jnwzKzW3TE1y
aHtMARScy0DUoAddpmEQfWbBnytwBCM6RXzACR1yTG/dwbt8kYPtLx2zDLuKoj86EbLN8kAmlFDF
p7HtxUjmPDWYv1/8DkLnSg2YQjuSYfMFYmRBkh0+IgsK9cOfuYSGC4uszVGq8PMzt/AXBS9u/sPg
OJT615lGWp4VTZHseBQd2BU4bGNKk1fEKtwShDAIg4Iai5GpySlgZyU4rPfFqTQdfJhqc0WMzppL
yz51IAl1IAHuD4AzOBR02Lq8k1u8Q9MQQnXIdfUwltqJyBZ1MOp76I9OV+4BVMK3Wn2THfawvDDT
kqRmvb2ERMuj2zW1zk34qE7E/WgnlkmpTDuJElCB0lRBmrdXzUrNsVi+bHO75h/pitivXnklSiEG
kWSbUvmDR8zYJcYioUw1opNtezT0wYMbf2LVrYrt8wPZTIk8cu3F/ZnxNeYSDd3LQrdTaZnBxlqf
L8mibS9BZsSChCcoS3yk2SwVdqqMvPoMaksH7OZaQhAvri3Rl3ipl4x0s+3H4+Yt/E1VVw4QdoPf
7QWtN/me9aNTeYrR/GC8OEAg2NvO/ow9FxCCSNH/4kXz8QuKhYGmyjlL2vIAotZFdRacEFiWC8U3
caXraLV170XDNPo3fX/b7kVjaAO6897kOB5MdOIyrpjOKVXi+/wIoyWXBs1U++lVEPKlPa45VDGM
v1z2w/15AtzOzEvCK7kUDdNGjrdl3/k+gOeqYXRouhFdeyv8Kv9FrOolgPc0uaMLG71HeITx7mRi
iNjSdI4A2CGtdFn3T2CkWIqgxcyof/WG7k2pf/Lwnv62EGaa1fT6bQNhtkdH7T5jpbG512xBUbB2
+GqiYTEFe37y82Yvzc8X6vAH+K3J/EG4udGJjbY2diRs4+053Rf94Z8swkKOIeiskuw1vHFeNByX
WEetDdHnvoYRt7kunIik6kxr5BVPuPetD86ugAS2YPso+jdhIvqLNgprlKY2KTcWxh3eqeq447ef
icnmT+Y0VMExrlhS4HbpJ6gjFwNhiU9LeBqd/wQNZ6XzIcygH0wdiHDckOlolXmIwEbtLY5+f87i
9X/7DjB0XWja2/3Wi+UYhTItoy8uTZF1b7+hdrlpy8Q9Ca3X4HfM2c8ztXYqM3hLBx2ZSWppOf/+
YerZUL27hHLDb3bDkFkl1uB5O6O3rsy8ey6YVgHRRTil2nRwaVtuarO51/Uye88D/IssSJfFOFIm
kK1/295YI5A0mbhfKU2AC6wheyNECjji/4OgOJ7mtA5yxd0gYXlRhNebsUW/DJxfI15juVR59fZW
wEZcbznAn5Jx/EgO33mvTGBKpVu9DeVmUh1Qde3KacWHZFRLsjAELwoLm+iy9UaFutx+K1x4hYcy
7LL4mKbd1yKBAS1TYN/MNu8mYk7f1iV5PAqZCJxuTDacp17GZ2CO942ZcAVt8KFy0yZAPTlahUum
ZLeUSphM22G212dl9iAqI6YU7qwpKqbVmY5M/esVmWRJMI6ocJIrSNsF/w+PZUOVEjr8PHPl4/CM
IH76ZtgdeTT7aBuLzHstj+mFTqXFPgkINBpJEdTdun7b/jBBWdA9DAgPCcy17dtyu/s1K1detkAX
LrwYkCUKqPuYovNfhVPX0HFwwJ8saDo3cHeMftnZWjoyXwzDcP+YlaE3tx2zFxx22bRO9QA4K4Lc
q5SqfJR6zFs8M62kBAhjQ4L1lUDJVlABlU88j5p+08Q6Sz19WPcG+gj283RbDbSh0igljHtt1SI7
Dx25fij2ft7Wsmvr1iEHSvNRNQMVQxNndvhTsLVx/QkMeY8s9Zhd0iB4RwmLNaDyYipYNZpb3Bvu
WRdSI4irhw9NaO13H2s3/VX9wyGvprz18alyqu1gIqQHFx15hBUvPJTfJuEirJguD5Vrgdhdi9bY
yXjn0+Rdj2Ue2V3hItykq7ree+P40gnggGYUDgPWZed0/bmIDGjbJmZQeiwf/Qld2H0TP/JEyJbP
cIODFwt3EaB/BFeQlWzbQmHKr1iqdR7V9Skq7KnDSIipR3akX7Z8078/C/p6Uk6wXqnszp3kMyWt
+C67T52uRTZ/y70IYmS4ZWuZ+XB2IB/Q3AQeS7O6kgPI6m/OkWTx54CMMAWdNC7E53l+x1H7tXwX
huK7kXk7FjHdNOkKDb8EzkuHW9Fv5zy0Yop/8HxqVyom1MCs7W/QKk6WK1jlWvRF916uWVGztY6N
CskGQD0it+v4NtySfYwbEq0pT4eMTNgG6UUjqPw17o6kgnhiuX+e4dfSwx9/mEnzZQPJQQD7k3au
HliBHWVv7q4z1Kq4K4d9rvR69g9pfgNbCGefvUxH6+3nWf6DQDRee6LT/gh7YPB0J1djISFntQ9U
+PBJ7pxEvqJQ0Yrjc5N8v4LSs+NIkr/4iim/RnMG4/8dJhi3c4VbrFat7dBT1dNw05nRc28zZZFq
y0sG/E5h5xGaI89e2XcqGgJ0XrsjkPAaMSgCuuorU5gqGk/OviT3VLpyPwYPgBIEXVNwQC9XwW6K
J4jTp+I72AmrlLqsGw3m6j7v4hd/yD1oRuNfASAkbhwMTgjXEuwstEGPfedZOze0HT2oU7FcbiUA
7g9V9z3bOcWh/+nRxDyYvpboy2yWatXJu+/uuLV0rHlOqd1cmNpGGk8UuP3puzFR+Kl8ZNc631Uu
NziAi0ntS8I2xLn6cwumOZhIpuwZkOwkMIWoKtR3oYLGCIDHKw2BsQA+QdDHaMYKpZi8RNp3Qf3l
nvljhmoE7402PUYg3zYGCLOGlJnWJbtFPPQFvvGpUJ44QRrIrvKdcd3Ze1D58TiJsR+nS5+Qd7fR
AfXC0tqA7DxlkWGDq+rYddQf/KK07uixiansL9qQbb3FQhGelAwrepJWEoadRBbSrw5FMHlF/k0T
sTwTNOaMdJWWkiIwRPr39UASkOXjQvlkGp0LGjdRESs3CoKlXzSrFTBFYTitssCeb15sXoSOZKVH
MU8Zkqbbt7tiWCqoJmph0fN2wucboudH9LGeL7f8xq4NGmUO5qYHA1GQV6LoHFtO0nkyYLadScfM
UAkpj1BkhKsPHwHnMPQ6t3vIkh2hOutJO4+ozZJ06JWe0jPScQ2tIQZ30To8skl/laK9Wmck6GWP
Pn3xKUG4mH6kFVdSpVak5o9tUoak7vvmDUu7teFI3HzuX7TIPzopmktZ/pq4JlI0NORDVUhnWFY6
JPSwtdHA6snTOYmsY2JTrDdm8BmAMlUL0t/pzbitZWUPx4i8LU57wZOrj4DyTGZ233j3f/QjUWjy
YjdC0yJiFeNwTRnN7+IfHsS/tzIqSLviZXwDu6un8YqsgAoB7OIovYGjyw463Xs1vhOP8SDkCB8/
sJQLfsbNMozZ/kA4pToT5n4KRUBARy8VZImegxKMM5ErqfUARnKaQk/+YBreckgbQ4PcCMYPCA8K
aqOPQNXdR3z9e2s0nCH3ICoXsMXxgME7umo/BFTh3Q46QNW8oeO/6whEcg8h90U8M+EOj/zuEDz9
vl+PPhodsIWoMSGUESyudu+OrEDPXJRFC4FUK+up4v3HE5VaFF1rTZYQUVbRGuJGUx/R0LPpTy5+
AuQc0kJL33y4w2FO9bgx6I6uxD8rghzaNolPywyxIjYWzqr3Z4URm6FX5iHCWDk1UXZkfkq8kNoW
g/sC6TJ1WzuOnN/YsI6j+3dvonErfiBYybavotcoCB+0TopYeUso8GNWu3H9joOn8CNa2BlxW0O2
djvZdEFAb7qDEoaz5P9GCNxKiwMFGHr7EvxPagkOMPP6GJQJpHyKmtrIzKjBljEvHPjh0Ktipi44
E/L+9JnvDVwBFI0QGWAC9hBkcJWKR1D0s1CclHYVS2CdCxO2DFqhsHceKFBFMnveLL72ARryg9Uv
g9PHtVjSPTK7XX/0k+hF3QqGeYs+cmrOlHjMXF4fEfRov4tvTI/Vu7+4CgEkLD7A509Z7fPsa4GS
Y71z1dAGv51GB+NW6a4SBxXSOlic7721A/HfE9F8xCmjpG5xZc1nIK343lLwqkZ25YVE7RojKdj3
SlgMWahWIKMUIyuQF02tFy9jJEbA1j+xfwb6r6hzkVRMkenJdbLCkciLkAEpHoxxqRx8wCFNzxSm
MGtgBjtDbHvaxLfGJubKSdBu0rqG6O6rAyMokRjepJOnSdAFXG95G64BSvGkGV2ls4IOUJx14E69
a7zNInPpDTch1+m4l7fIsW/iFk69nraC5bjosU0PHi5e17A6Aoe9fhaDQ8nJVEKu1hlQIv0pPHCB
Mx4+guZ7NWCk5RyDlqGM9ocmlyN9NViT8FwKAcHctegexc1b/kcnf07/KkixKtneuog65o5T19zl
fu9ENgObXYRpxAMrveERfRWUwBY9gc0NXHQToi6TgXgIGy4o7lVjChZTV1dJGIrz3OHKDkKOO6eC
nD1bmJnC5BL1VnyHglw7elb4k+iiOsD49lh85dXsDFpHExgINko5To5ccaWzO4Hg+8vpb5TTI6h9
X+dXO8cwcwmuHxNPJGDQY8yE37nLh43B5VcTuJdUb+B/JS+EnK2c3bFfHy8OXktaaap3Dm+zQjx9
9ycFJJ985AlDJz6qVdazohvwMCLHhw4I7ABQmuX9z/P3LONJHgxKkGdBGObxm3OIUGcVTRrK0p8i
mQn/tfr0f7WKL2En3AH4r/CMihpsLrv1gOrb0y/v8yoAfSLZCGOnGw6Tvosa84WHfIbp5WdpPFWc
DT6j8uxfpG1yQErZVpp1Gw2ArIXzWGc6v9tn29Fte9/WPmT9xWT3xIwzv7AI4YhipT+yJeW9jcPB
pzOlmZdIbwO5Ocmz3tP6/IgIq5bxe2wEsqTJL8etujIUHmkKzQzkW/WRzUf4TTB5rLgLoOrUrv/F
xwYWdfqP9uMdHt8+fa/IXCw+MJ+WaFLiAGvMohvoAmLcZ23mgNSqBGWCksGe3UgZlkRODkAFcjMa
7ohQJ7t6lDyyLsHMedUmsOFf7hsmnO/TRyGFRIjP6cjiUbC2mB3E8mWrUHIY/24EuLJYAMljTru8
knAorxEPQlNOH9Hg0wxnzqH3x80JbYb5V87EsgJ9e6IUBuDLJOqZeTVyPjHRIpgD08E6FqtG88Ei
4hCpTLRBqvcsCw9sdfp5Q4nV9UOsDADui7yVdyjaLTP+U+5obx1qTUs/JVw6hgS790ZWxgNSdPU3
yeRWcpTPo1XyToH0LfS3aVn0Wrkd+VrQs/hxMv5f/+MSjNSKdx0gMx0ExJj8vyyB+P3JqohvzSoK
g3Z8NX+h0Vs1J1+oX1/DJ43iFwttJIOwU4FfBE1d+TNz5/jhis4hHeGsB648whHDMkPg4BU9WUHJ
B6KVn4wXgodtg288PuVAAeSuAj9l+JoLnnQvqzYPAJ7BO1hS8Ps3E4cqfuhnn0ysMd36uSJHTZb0
/yk9zZITInotaqOoaDJX6cQHo2xTqeYuJyhNYK/n8puVIUTZEfo6NzC3bYyOK+FFil8YiqoHDr/v
90ZCKcAYtwTdR+/mkob42k8Yg1tEGqBh+VaVSV7aBNuMyNjjSjgU4qOXsFfUiGYBsuVkRjCPNJzd
SRoxY2QJb0K5Tfo8zBDbrqpF1Q6dMHxMRQPi5QdvCAEYf8tdrwTblGm9uqFRvOgixDf8v0NJFWGi
lAiBnDtTJgA5Z8nRWz7pOWV3+dhm8NmZAwqF2X/SZPJCVv0PB2BHTBr9rZmhv4x2qvs5HZuGlS9X
aPHLZi0tNluFT5MOHcYrur0gFYkQ1Nt9SK4gy4tTc0aACPrUTJbwLFt4nlWMMO/ZOp53Jh/lv95T
jwg4DRcWB+IAu5j6Bw9x4OsEN1X2jZaK80bNXRunKtwykKYiplPhr2MbN7EqZ1BRQ8UjLvs04NfY
4mSJdvr/hmHA9tnPDsPMs6QhMjtf65IkttxMtox9E8KnVbwAWez8r3RuNXRZ2PADy1+M19SFOrv4
CnRHa2j5EPgG6MUO0w9IeKmykyF990LlHyT3O93xzwxgRlzlVBW2xIH01OV2xoBMO2XwWjw4B3iH
TMq2GIMH96iFzoGCRDR2vOTr49jqbooKWl6HhrOvkV+dyZSn7MfYYJtGp4b3NOyc9vN6FjK4GbTU
Unn8Oq5AKkKtjQzGnUL69N8OvyPl8UpQdaB1xooCVcdBVzIcexnvtdNAgEkHMPK7SdyZhe3XFf/R
lqVX7/pcWJMULzFCpbORxiIzKIUao40enaajgQPY984rLhLxz94OCo82G5uo+G65p8Dd3YUDuIo+
2waKDhsfKUwD7ZsMhgFVgBmf9BkVZAHg+qH+M9fN8p32DoH71JfNyh16+jKgkfqwu4V6LDoS1dPt
/EbPMYQqobthEsTgQEu/+KLlrxz5mmhz11HaqLUfdvkVOzk6htMQ8j89fDs/9KSQeAJ7/wWigVEg
xe/kJx2GayLhNdwNgJQXfVLNnMFGwZVMqMclnJmtmKW1FwKWDhlOC/KCGhjhATHxSsQwlaBv6+wF
8F+1ly9zEeBsaUjW6VY4nusoEhR94CT4hS937XcdBmW49nv82Dy5Jx42q4fAIAv5CsJ9/qUciDpn
3zOjj2IEsUoKClmYsYZumVzyTCg5mC/9O081oBSc+nBoz44UkrSx9b+LtjYSHnD9GvSRPCK4YIpx
demYalPBiLtmK0RtNJFeB4FgGs/nTKeYAgHeCdGKAlPuZclLyyWEuoAvp7yOJWHWsGZvXaleMY+w
lsl+RB5y+r1KI6xGZXbfsy6kWur1UGdIDUOT4ovqAAuTOMee+nPUm7+n0kKoiX/ALZLhhkXLUW8/
RWHpAZ8vGtJbvYeHvI+eO0fO3KE/mGokJD9MVUWbt6mgAdhNQ8MSS1gkREroLUTy7GiyYRBaqM+w
22NITGu8e5rV/KK0HW/X4ln+a51blWAhY6FZJi3GAEgfFsR6i21d4o/xBWJaOYz2cjTJYLm5Kozi
YXuTgR7IdLv5uQe3Fruovt1virDJeVQbkWRPHcpTpOAW8C+yLyhol8oQnwx96RGiHNdxrIomVlDT
DAghTO82M2FNnQgAbz3Rxmrnh3rfR2FGZKDdFGpj/pw0kayw+C75kdsN8hCTDrE1zndOQI/zPMoa
/QiC3BXPJy2+AX7NZ8uoPnF1gTXoIJg3jfOGnGPfHM38p4i+rDFd318IJuV2CCdQgYiMk29OIBDW
Tg0EBuXqtVK0Ugfo+Yuu2I6g9Q2oKjisM6GNgOJ85wHeWCYyLvM8WV23V6e/odgqt0IycPLS+leP
lJj7aFNsVg+0wAm7zaZsi86M9KeSqOmUMp48Gxf+9j6vy4ymSwNkCawhfhCG8v44oevbGzR3qqQH
RhTj8R3mYet6PmS9q7cP0fnGnWMKBDunlyNDNrN3Nv5AFB4khKhOSbBlgmJ7YzfEkPIa/7MfCwI6
YB2GBeB36WYoGRRDb6HjjCV6iOtBeLFYQeo0SrKZ/tdvi9obbahEwgLldUJL0DYUMiIPND95At0T
fjAg4cpDNFBKla1AU54h0dlvKkvufsV2etgtKjTyAsXkECxMWJjJ/OrFxCLMYI8TzbW+NkHE5Awa
VJYFCpsmsUNx9JM0jppSZyL5K0XSrLHOY25a6W7/IR3L/LJ1fewcddsGyhcQgw7GMOIfbjKiDbcY
IMPSB4UBBRsQs+zP8A8/yW9OP9lpu6OpRsAF1L1iBw43qe3pr1oFtWxhXS9Y3lxqgCEvXrFIN92f
IoxuJKt6Z61XSvSQQnmvIw42btSiuxG++88PSZG1/sEkWdPMUptiv/gXXIYW26U8alF96mxnTsB3
9DRT/1s4Gn0r76o/vpCYgE6DH56TJBzqGryzN3QgD1D2L3JsD7pX2ZMp+MZp2cPDLfyEknzNgnZe
Ct83bdu4aNTkxeH6td1gXWAexHt/3YV04pjDUjRvG2jrPp9ijK4+SHhWNpSV4X2AE+55pKLc355l
QEh8OWDBCkEiGOuFsh7LeL+8oq2ZJ38c/BQb2KdSKtA1pwn8ED8l+Qxc/NiZwKfEsJGLdrkRdnpL
NtbN11QbJCu/H1sk1sbYQS4xDHm66jP21irL2okOBFzQ85GCnXJWCCROFrxEG9gCd4G+M4H9f8WN
+0UMTbwPJq8LNom2OV1S4GMKX3Lv7b4JbXacOQ7uMeB6czc6iTZ2FsXxHAL3HKPtRuM0dWnzJvrW
3OaC4uBw16dUB+sID+JCoyzftqvA5F9GncQeGLdiHrEbOMQ6GRLxBtsr1YWGY40eqaO4BbLPmJyX
iwESIT3WFQP2lmUH1rzWX8QS2u7Y0x2JVPatPybeXuIDh3cuXhIsaZB7wJ/GeBPwlbAb738frcOq
GRwO0ezzMaX42YKQGxVdjENCB7KQ8rAhlF+xJoviylBT/jrYHpYpFgBxjQGKlHV8BxGKmHVryzi7
EC7ekIqLQWsI53BoJPYtnVUhJwaSQH0YyOA0PrGyOkvgdtf+42/D9y3oSkJxwa3lzsuLt7Ur9N2f
ryD67GF6FAPVBem1fhQG+j8IVJvoNgWFRhKDrLPAU+eJUvk9MOzL662O90H9gAgMWsq0sUQkyePm
fLNjOWNC3WnM0S6wzFWny+87DjKSon+b5dJKK5Zlm1rK9a6aoWT26Lim5ZQ3+GNiJG/Uyaj781pY
gKeeFB0R8pONu+vla9pJgy1dHcEiCTAc7WhZKwaFPbHjRLAT86ZMO4PZcu1Of/MX466Ae545b2zG
B5kSyA/F3YM6fV8f2UzxIpAMpFvzELZzzrmjhP/zP9WSVn+Y4GtbeMsVb9hTHjIvvXjpF9ms6oBR
aXNX5W01wdfpqhNQOISrpEPJm/c8SHSReLI3QKJihuE8kJ7Tyf+H9/gxo2k0mTPUjMLlhlMC4wap
L2aZGK9GRZJVZyDNA1M58BrjvAwPIkSKr/fG/5HQrJ7edfcwArjmX/X/JuRHnFNbzfkgx4VdY946
oNawq14XGZKIEA1/Qveo7XJnTjWltf8CKXvfs/Sp3M1qJVqxnVDY2Sfo/tbswwf3wdO13vTel/al
ZkmPUuyFzVZAdrYv3JOBYHUCHvxTDnb7X0ExwBenH1k4UAaw3M1krk4WbI7/eDv7QquVjcqu+yzb
huQ0nZheeNew+aLRX2+BCsQEJL9BAQ7/jFgp3BHNiGOFGJcJsdzxRWzUI8xe8d6GBAuGuWOovcV7
H6JF1pIDjiqPINfjM2bP8AemLtojSLRnZp2ZYbZpyRrEzNva6rOGN57JT+D1y7YoU3D0YEL2ZOeA
PLK6/uaAdcGF01ekDuEMklyLOPta/RgNGSWPfPBOvsD5ZRnQh2hS2qYFQgjUomud/KtjXfru8Jk6
GiP7siOmb5x7IUwFWuQhpJGXxDus9c4t+aVF0lkyJT1cllkuBSbHVJk/7wPfVqz+kVLmrOmoPL3I
0visGtNvk01z6RuNdXsoWXaU0cjbJiwSE4V6N8TFI0K434iF88ZWKvglIrmVIkx+IwOIDi2kAndj
oLKL/BImicctk4f/etKUVgEDrhvjkFkk+zS0HVnWUE0UZ5O02Un3OTkrT7jiE5YmUjAlYpdifEuK
My/tdSPvUyuFLVtyNr5zSMfgzKrukNyXdDwjNB5Sio4O21NvgRaYXQHWYmFuOyONhcpbRlKZN1ox
JygOJKHfnSWY4FrDdmscEeBovzFo50gSWZktcn6JJH0AL0xPRCy4+80cQdGeJh/MbUGRBe7dP+qB
hk+idOk+DdOlLy1234s5R9ZBbn1bD4O6rwjSvHQRVVrC9OcnCCw7r2qxv9J368m3T6+AKrvBnKsC
7yzqjV/ek8ed6huD8EPnSUS09knssa6y+pyKfMBMOr6ADVhICQ913deKnbULsnJNhRXlsk1Zts1B
qtFAF9vfaiWl4BZ7GpBOqPSdOWKgtQHqlgd+fge0GMsS4JIx9aXq5Mu9/HLdqC3iHeZcm7oKn3Jo
WyJyn6spvSEzTOrVomDUCt9cS2M0R07/nfRQaiMF4nqQXdD2Niue8ajEw313KV6+GdwZCl3rbDNt
Y2b9h0Zy23INkXT6kHShXvL52tUc/8W09DIGGs4FdmFjfjZCfQnQczHhDgczwQlaTYkrTgA5Ek8g
afYfQdwboTJf0/NwOljdYAxkZ4yVKjQ2zo64gL0zqEYeqhqEOs4N0m4T4+Cmr7PUqFLFokGn6Lu9
KqH/hRCKcXpiz11qZMmxUfjs0DEHj+BfnZ5oV5HKvPU+kL485q83IWAVNuVuKaA1p+higWdx2Bum
+n7hpscuL8OTqne3At54Bk6HCCTKk3UmU6wtf5WzYY+AoCp09mTERICFX+YSVPKgZE530U29wg1K
ghaDrmRR97EqTYDDmHzTFHvaEYbbv6kANDta1PeSVylJcJKXLXPorjocNpkSe7wOCyUasNPaBSCk
lsO0fC1j4Fg//lQa7OikNIKboCt4M1B3hWo/0ZOxxPTI0WaylFbLc7rugCPcIirLNsERKno1A39Z
R1bebgtFZpTBICWjH927wxMG0s3F+FyjCn9m0hdkmSr8gBqUeBK5d1FVlm5y6wbvrBJH0oN5dRDB
EACo31tUcWn57ZnquJEPxYF8nEWLz1QV9m7HWSUvFGQa5IswIoaq0PMmHABEZ16j3gMqhLZWu4WG
xyKVA7pdp7/CoePMKvEbgjkF5dadg7AFbg9DpKCo6ZTnekVvAVwY3bzRmj/R8CXEFPVVXshHE2Pc
A8Rd0JhOyQzba5RuK3uIIbRfnlIOaTpEznrvgq1w+riSScZyPb8iH+TydMnDUUSz5wJCTA4X1/6B
PJlIKFGz49/hMcCk6zRlwIorJHzSjNlrw1ukjWqPwcxDIxEYlldqBZtSXSVMVTMLbAn+c8PREGGX
Uml4vXQPJOfO9DZiXLBdXU7IfvAhweW7TWjUHHFxirnPO0OFpoKixytJQ9Xoj6HyyNXgWnDGXKks
yqa1S99B3SdlqKvg2D3X9qdQIXMw0VkDF9ZYFH5IdIffmIOM7mPou8J9ehMSMns/m48Zp1Ii8hfR
65v06cGOBOU5N/phT6cpE2A51iaMxheUWuu8JVXnCfem/cXOqy0rFCoSGo2DfyiV2pWtGrWb4AFV
lFTAYueaBJiGrfFqGclQadLsNw4E8GtYupH0eLKQthgiBzTyLUj8sUXASLLA+5YzmuOWC4QhTFuV
W8xclzWEbo0/i49PY2ODMo8fjZn45OMtJTHwtF4B0Qg8jPCWkUrQJGz3WJa2huYALLCZ/vssZbOD
4g8YX/LxE2z88mEzIZ9EPpzYyoJJts/P0AxKQTelaA4DI390Au7ctYBYcOUKeroxJPieIaPasJWT
6LY3RTMEVujUbsYpdZUeLalbIZMO5mHaIovTYm/hThhbJmJufhg4nzW+t2j0MNrfMp9WI7wquh2t
s/DQlBY2FBGanIVZH6E6Pb0dDDP6juu7RNAhbPmaKalDVYTtlP50moguKV22M7ENgpHRcF3ERFvH
ju/RVOt8m7SqT56GCzN1hhTkgWdkqmsUxYXvjyG2uFChlvDZm4FG1b5+q7OWPvUGXMRNH/q/wD/c
b8nnWlFsvRg10PlLSHO2kNXuQrFWdWIJpsQsRsfNBl49mwkf9S+6vFAOLIqDjnWng1tGNGL1byeC
TDZKD2o6pvuTk/qrhkeWEt/jnQf0mQxIjXRamXsS0NJVVQDH729ltar01jLwsgBUGO21Z4ugd20f
IAf7VuYyBwBEmDOL9E6gLdOEzOO1fpmeOxs4xorF8WCfWmRuzOQNi9JHqFmCOGXaO2dg8aFwFVib
4bWN7OYEWgKpKmzqDd94aXeNdWV1MDYGpn3OsNUHDtw2JXs42BOqPOBHhQsj1rpIe6wRwI/SEJTo
26FVY1G9NOr7qgQxDaVJK+nYwOda0DdrqhWoo2mlTrS9RXsdyij9L7XnX65IqBQngQ35ZtxPMoDr
fQKyQlsMKVf2PPLh+H/G6Pu06vODvGMYIiMT//2N+0U3dAc7nOlWx9rcJ8cGTWBuQd1A3+89sJsd
CMeO2jtSevUeGfYUAYVY7R3qAOmI3imiFmb7+dZ58w/wdtVEonvet2++Osg1YbXBQgDcTCYkoVG4
uy4eEInnt1YsWsQ1zGrf82zYnF8oaSuxYITho8tjLoMdc/7eWyxhCnFIUN1DkZdsQPB2OkyIsIXZ
JsWknQySMVdqWPIQZGjnUgjXZ1t+e0eZYxi9qM6uQ0BjiA3NmPoA/n1sRMPDqXbTW6rUXUhKEvWM
RgSYrnApaJ6TolMp+kE5lm0FSaCKcdKgVHU0jdUpgRLK6nPs3lnT/3ToXT/J19/DVj2f3gu7dRqm
RyefbkM0xTocxdbI2Gx4KZj5wJJAJFbUzp4ZomqVHySt+1itUnSCzDHGAEKNT3EqogVqjW53zy6z
sqSarFPq4x3lnVjWu2pZWhSujSmA3dSbAXd5mxHfTFOVx788iCiCYjZnzpoSvCg4bJepADLCp49x
oeBgcFjV5XAwsFXVoxj6WIWBawtJk4s2GKe/8GWikWDpuH6bnfQ8wPmxGqqx372wSFegIxPVd8Sw
rhmffdphKH2bbDex7p6II9RR3iXEyw32Vo4j1sn6DRJVXV5J/qxxC+ybWOArvR7lxDbo8MRqsfZN
nmKr2BZLCWJk0cICg6iC7UJT2kY6ucfCaq5dobd9esEoLRkQEttaPeNhQVGGKASbU/J9wP5d+dNR
p7yuoE8afZC3OINKbE4MwAnkUxkOWlZO1oNF3wV383Q+ou1jPtaSviiZ9qI1oFcqLEGjGJ6E6sQn
c+d3kof3hGB9zO5CvNUGcnquYnJMqDSAbia+mWot7lUPO7FHs0nwiNgh2SiBvSuhuHqUVoQiFS0m
ghLIpVdu4rbAwfw3XsWdJSU1BeZBvQ22L1bGTp8crV6ZdkfqLet6O6ZIZcc96iL1n7xBj3ks+YE4
OY1j0nlq9rauMsox2jmUkQAmERf7Zfb9d/zij9kg543nVXEU7SEjDQhxWoq676KZT1n6nUGzP6jl
ZJh7Bd3LugInZYlYGJnRNUvOip6ouNxP0cPbh4oYagZXdsq6vuDUA87ui+IvAKQBQPd09c6gewD2
upHeDW9LZ1FMNZzQrV1qiKdaPDaBLgXsBmkfhYmhk2X4EasKvTKQCXUAQBBh1Rz13A19RsBhQ//B
N3MtPEPRk614pcqtNb/V1C+3IpQRa3pBvmsvKvV9W+IgqrgBBEYF8g/oCrW7PuyEKtGpIkZOQ65z
fr9r1fsRD07vgRYyh5uoCNiE2sWoouAs9/A5fXB9yfAjPp+cHmQArSz8w14/QKl691B7gKr5Q/bi
WzgEktjxU2Oc3t5GvxrQqJlUNXup7mWk6kb5DBwa2YWMhnfwAI5pl6YnROBCzYw3IvhGwhA+BJnf
pFFOV2DcE2shW5zk05tc9GUIEvkLviLpjU58Y/6TBaj7dJSYnY6Uzwj7pBPcDhhZFBTJT0rnBE7L
Q4iYPSeYLeiJceEBrAK9vDGG6b3ePi/x9mafmL6shyU6zxZhkYzA4Ps2iFLjSwAA8oZd1YJHWt3J
ve2fJczUaEVND1cvRPLZPcmgCSyoToVEU6GvBxScZbDblg52Z3YKhgd78w1J2ooZ541IRoa9xjA7
Jl8POJWQjyccI6YSoZ1Ww8edqOrPX6GP2O7eslSQMmY4r7L+OyvArCvcNqOpQwhiiDyKs2A5De7M
6Cf8LX01pp5E2P8hjFMO328aNBkJ+0FGowwKWx40gv1YPQFrJOSuJnolIw/ByPyMJtSBRJX+RtBp
BgYgss72qyzjLvMOJgnfQBCGJZkh3iNZHJ4e3bDtdObSLDipITfIbBiSvIlyprwinEtHshV2U2QY
7h5EyKL2y3zEVhsLqGilOXt0XLmrVqRl7v+4QKlXZu+Z9hROq+EiVKPWeq9gvGTyWxgJ2M4iy+et
H8KvFQ4Xj/shA1NszBW4N8MCxgc+OlniHqJLfTjOOEnUD26y5opqlAHyYyPDE93CTNglLFCg+STc
zN8ShMH+1buSk/akxzzs6dKYGy5B1Nw1XtHK8Xaf9I4TCvTS7NgsE8tTleH1NSaardzgL7OIMQSu
g3iUP/Hs8tjKARpPMbxmoqI/K6XpYgzCkDlpgQ9I14eqoPcQqfZs9rgPpSxljZGwp/Ygebwiomhg
EUNn4qIvbicDj7GkHivJKRSe3tZrdodb2bcyRf7WYD/pxq1LD6Q4CyAtawwvF5FjXrOrgftv6+X8
R3ChbEOicCRzWr89+mlwnH0w002oqqg1SOZLp/5mAyXjoLh9i3a9xztU6rJV+k2D/niSYW0vHX/w
hGAFUDSYOXvEK/WJckbJhe2j0Hg+dWyWB8G/jf9NA64/d7dkOSzeFhFMeSCK4ywURWh1j73wdl2m
RUSLRnHaV6DGdx23jYPlPhAFmHWjv1Q85IrSAyT4nMNIor3gf3pWB+bX70NpNAY2nqfexAeU4KVp
wOXeDxFeuEEe0hvpUjFlvRshgoAx95BcigUQV587Z4abVN4ybv+vl2o1YUU3PqUdfKY2HqHeemoK
XMcGZldfr+NZKLdjW5ruDdpJV5Obtk6PVbJkSxuE4qXrMIJjlolpUVtkG/Dnx33PiInZiuecVBGW
kFssXauXijCc6TGyPSggjT/OA0IdjeN+MXTdw+qcL3VCLYyPKnYZNaqEQ1fdazH2eSdzlhH5e7TI
tq6TXsBFPolnkEABN6QvFj+VUS8cuYcOftVHVWEKz3kt3VIJzTlWhb2Q3yk11pDlCKUnYpoLBSqU
qep4b/Qpi6kxRrdkz2V3zOUEGeAKaNsn9yzmwoXEdX1hoUHM2RVuJkmvcTlctFM4DZ98e4c6vdgL
WkpDBwRiUqdfzfryr+DN8IxQLTc3Dgq1Cn+CU3fxz2sptA3hxscR39K4aLH25sAnFLat/E5by0t/
Whap0ThZjhJelptImrLbVGoJIZMm0yYIsFo39mitcpQinkhni2BM6xTWOXz/pQeLFROvjU0nxqt3
4KuVxF3s9AHSJPpAfIxp92xNw4bBRQtw3tf5YM8xwyt2myCdkY8e7C3jpXOEr/7XIG+3pymhshzN
uAkJTHXiuz8XmGTpZyVyRbKFpeccNeB/33qNdSZkKtV388XIQv4ekCDYKaJ0ipGZRAO8XX/L5Bmc
6WeeDHUYqAwBb8kr+faeoWYzxy5i3IbPnuWEuoZaR6m6zAJ33AFAzW3byHjY3WflKoL87ViKVNRQ
VSGKt4rnbtFUM7mVE9Wj3Y1Sc9N6KaAitWbtryTy7zhP2zoCmjG+Mfn974NStdQL+//g93TNM8Sh
NiMykaOpRwFVoNyviXRNT76aHUzCXYpBFHjlqzZxDdi+bXTodZMf+9yy+fLIEuE+PmQXcppsOFfV
tOE8nxyfauvya1eFYnB729ynAhaL3sHUG+a8qkPdNLBs3ENkhNl7WTKb14vFjpr0FABnbDLTjCci
AKfCYB9SRrK0luupbZOd+wNt8pi981XJCpw2s5rfV8GXjPjviwobhJFSCrUgZc4jY9NdKQL+GSLu
BcukJBhLjsNvAKun1KF1kZEjfN30qiM0LGfkpgn/9lNGaL/cqwMt9OrO1LxfDjBxzWHftTY1brhy
EPtaGmWQncz+mckvsDFQ856gEmGs5X8blCyeQPI91/dQ47nktJ+CPolSzQ6VD0+Ns9oMZhx4v8Q+
bmBIOfrNcUSrDtfO9mb1cMkT5YxkBxmZ+13nD0Ycpa4HsUuAjs84Mls6aKdr7fkx1Vziq+ukwXM5
+EvysaWk5Wa7FwPMjtFQ9Il/r56oWqcBKABX0qNBCKmod49Xh8HAIxWIr+SG0BCs39QZ3xn332F4
qoVcbZEyzDDoYy+bblACAMpAaqsAQrljwDoRENvJyHEQ3WHx1SpLYoD0Dh5tOGrUfpKR/usoN9h+
TpMiUf0YFdR9fZiUO7ax4uUSDPYAjUucxgb3LQMexcvr7AcAqliHNT9IM2o0aYe2MQ6dRl+w5Ip/
+UKYN1n4iGE2UsTb7+fdYNyLt3Evncd3wV+UNvmnJbR87drKOl2wRIOdkRKHSa8vFh4tGLQ1ClWd
zee+tWCzFuoV7yqtNU5uE7XnOymyZuWc/qp5GHZtut+o1bi++BfIdHS4uT+yqQbvvAuIDLv0MmC8
859/bcbf2G9R29Q3pVY6+ubEdxkIVU1sTvGL+nNKBnVnEh2sPkcCm/kVtilcacB8EvP2/F7EibVY
AFHBGwL3gpnO8K/epn5prFiJdAuX/SwEYo7WM+8hPGy+NU9ZDVnHXR8uN7zH4YaU200tBjEE2Flc
Iq+YjI1uzZb2PEWAIO1r6oY3ZlC9qu2rpoNo7d1++voLP7p52Dqnf7J/ESOwBPfqxafkEwLXVXel
kkRYE37f1H2mS+1X4/HU20vfF1AgPA0Z/alzYVSDkvawoLMW9PG53F25LYwfRbGD5tAJ/nzUtR0O
hTZQHmFkxeYd9ZdRkMj55nxzQWqPpOrr/h8WisAldsXgwpsuAFDesGRi84W2NWFkALCF598vMaN8
i1LDWMMVzquvW5bKhEra9OcvjjflSYXc/3SCcJylLJnshXZGECs/8LhNNsloB92I2n6YDwLSo9i1
bCtIPpgMjTKIUgRj/TQ8dD5ZwsKDMxqm0TtgtVHL2ijyCM9rjpFO0Y/6M76MTDz05yP2OwLgbECq
PWrsEDJ57ohG881U32nwjL9FIc0w2PDeVbIkt/DFPSfC4QTn0SjZ8pWXigr4qjJVDcmr1ivSB+lm
V0tibSJ5xB1ga49VmrgUdZYBfeCTbWoP7F9CG5v48hiNwVir5CCOkIF3SPhjYdnwwFpysX8WHfJl
OadRIhScSHhHm/qNhuR0BBk/ddH55WUCmoUiP25sYYXnSKEw8/TuoK8/gegn7iq4W7DLxdTLlRCQ
7xbpEu0ZiQE4TL72l+c+j8wL/Kttl2l/QU1EHVAVD5Le+LUYyiAc+mXbCK0/WBif200x36OV3Xp3
RqV70ciLaQ9BqPCYkHEW7TVmERsIE4nMA2OIpgZiUqA+yk62cAKkltBEbq9Y5n7GE9VwiIVG7gV8
VdyDFQ8lcIQQly8Gs7uEfJWAxIdbzEZA0C6dsUBQ/M7YwS7pDPJm6d73OQSwc2Yu3/4+BdegArzt
/qpHDNo5RsjLCCX59z0m/uWoFXwgrZdiKKsyk0Ps31TOWyTLJUcbMMt+SI5H+CQnTImc/9R+5k4R
0EynfKQvzXik/wwZ8F0Hf4iv+ps3P2c2S7mITtO52Fo5T5k9tVABSXAqTPZw6+5r6Lm53rEaGiMY
YPdaY8hePgl6GTunpW6dEkDjaK36UUrf/vz+qETmIlbuXCh49akKqOgIVzmiCmDfcApj+xWfgVsJ
jzsWWLEeeoWZdHhVxfBbsVpBjXBOHjX22vS7MWLHbN3mYjTTWTvZrdONR4PPeSSbD5XoSv0mZhVD
3nU1H6pFHi7jX4hIZ95K9sy3Zlb9Tvg/Zz788dzMZcwJFXMZ82M/QHdTdoZ3vQCMnUeSPM7I0bcz
50i7coZwluEZ1kcoXRacWAJD4CqgfkrkS7KoUWuhBfCW3I/SOxb1ma46/CzVo4s6eeXNVCYvlDE8
XyUjU2++VhSucsBMUZ78HK54cfAtJAEt/zRQR3Y7CkdOih4wpzce9hLT6PMzytovq4sYA51dJKjK
RNdNksOFnLakxm2+nWqnuGqAONFM8CoNXO0oMjRssGFbNrFViqwM2FgF+EzY6haS1ZjmZyo1XpBN
7pDBjXs3wvTM2XDTXpGU3y6CCwLgCRb1uQXf+OIAWPc01Kt/aXM7eOQgFO+Ly548gnzEFHURBMtK
lDpa9q4lLvo0ULJL8CQnO92SiO64PTxrblHPh7c55WT5+lt2m/8Q1By+tqlnRtA41kWQ0ibgoqf8
V4AAgNYbS132BOtvmFDSAi4rGPi2ozDd1QdRl+jSTyXo9jVGVuIoW09lMlG4vGcMsM6NE+1kwl3n
mvQWz+liUJEoTQ7KdNP20jBiddCSPs0JRlEYc+DL/gniMqZ3iV905TzPSq1LM1IAbqqHvT7U+hn0
Ypbk8pOzap09+yR4wb/VN9u+eF2976JUeq90G2kQtuhXtui5zPWsE4NxlfnpLB9FXRrCanaNG/k3
vJKBLzwsuiY7PhuwFU2k8pFpRPgkCitnIFI/C11FQ2wxlcZ/LwLwPdgwnXK4Y1pz7aBj9DYAwpkJ
CHc/7t90peeTQlB1hIYAaX03h5lsoZnbSG7rgU9JA+ocFltldea5w7+p7o7YhLCHYVPJjJ/brkJ7
4ZRJcs0ip6awgRD/1ixCFIvSxjUTJmWT8jgDJULfnw7hsz/TFGduoIxlfuOuqOZsOpUzf6+ZeieU
h6UCCacO+VBYBlZcdhbxBCY2LztJxVmGq17ueRQnlUMpksdF7ixzb4ZgUQwZ8oAK2hlzEUsMI7Xq
Tphq+4WmrjwhC6RfR4yaKqOPheQ1B40WNcEZ3kcsyMzYBtXeiyrdYO9noEGC5ucolJxQ/flMzhga
KpA7G0Y5Zj6UqJVD4ZwD4ooIlgVi/x4HFLq5vWsaw766GScDbsvfHLPeovKlVcMeuszfu4/H5zCr
FB0FloROB16IcoVGlzedgCmuATG4QRKLwfrO11zxDGbVhaA6o7In6wBmc71rMxTJfkIIt52tYigE
JI0ZYShLDRLVLLYiJ3cXsrmPmbQ1Q3ogMWDLLGWa+kNad0j2k9bklO4OvCifGYkv8jqa8kDt++AL
Zdoo49ueVi55pHW1xmPDvlotQ6sE6DNBiwcQGUmJ8i8xu9DkY3n6PN2CcAiQJDWpeucAAZFN2An5
jSxBf3mIUKCNGYMxk9/zj4Tkg3J8KSn/6RDkw053dNLRH6Ymk1kedKiC0it9NDV57pIWfB11aTrJ
aiQtz6ZDLIPjZ5I1Z366anFuCZSwIzgdJLoXQq3xAjN3qblbIdin0l6xuuF2ovf1rilFnL1vca5M
hLe9C4PvDlt8atxsEQQy2arteI9seLdlZ169UygJ/e3uG5ot0NzZ8rhNVQCEEmGqQwS30798hVVv
cjm6yfcgEIRbIIBwkpwx45CIM9AqPWjAtUyqI+V6qdHMjskdE1XpAUNQDdxtturul6Hxstfhfpo7
jei/zwpOWCBnIW7bQQbaFpvLx/MQ+osSxTW7EM6GN80fte2RKetURRqgmRLOtOQCG23uQs/E8Uaj
PxxAIxwwYyI2gGSDlpv80Ezl9PGnFQHgvL9vYEXIW2O2B3NtEBCFr/imVY8BHKbSkkW7ug0agQMh
vee+7zUOC86l1kQWvXkjcaGj+TC3vVNMxmM9AzBLt6RN/wuBsdtadvdNw/qp5w4pD3zqD688u+To
FNBsDZQ0Dwh+U0Dx2TDVDlRCl18v2c7SVFOkLqWW37c8x7UfSFOSwc3D7Z1hLRgcNG1PfSF72y0L
ThBuVcaKpJgM+x0HA8NugSicIWQemX6Qe0dza6BjSBnTjielu+4o8OZg6Rxy816bDxzcfqiqSyXU
R7dmHKNzg5Moe1a5vw+dSxK34KNJu4xt1kShrCTWRMotCvyv1zIQQbnEND023lWPaoPgm64jRvgD
QXDKFndO8YC0UnI1zi/OZ/9BvC+HzMc/RsD/gCTUEPi/uIAifRRab3nAi0DAwuzs85NwLhdeaktA
IWTyn42vhkYO5r7y+ViEW3X8L9B3IAgDlhpkLEXGZ/+t6k2MWdetpoT//eFhmAroUHp7VE86TBwd
g73s/8vXsbCeVcMi7YJzPN8TEaiiVT2y4tEtWUYER1ADPmVhqKZZTMvpGpzLt9w+GSnKmfw9EeXY
LcWe9MjkDwWi+di4lSHQLb4IfLmywnZqfwpN6OGartnS+TorGF6olgC6YS4uxN/nlre2XJA8ozkG
y8uUzlDy7z8OXeUZ8eW/guvncpVqCBG9vMjE0sVUQcYfnXZwwUHRuNymk39DNrJrCq0+ldyQ68ms
ux8ugcpzd0brPSJXR1MrDhxuQ7vlnUFfOuBCYpTtwRXUkC5YHfXA2d92BbcrMJHtiLondEcV9czK
EuTTyWLqvfksdGZrqFpmwVZnN2uqvR3XD1PxVfWuZQ7uWkmbWNAFEmMWgYHE4f3bCM2SMjJTCJ0b
nbw3kV0VHgu6R9tziVqwriywpKyyb7sMguEMh0KC89E8L4SdOVugzPeJ/T5EoK0bNJu/LTafhBmh
O9ZDLgnlIEvq8dLCsApvnEScoXUKryYdog5XOh/yNrJE8pTgTWgWCCmYj0vsnTKtCxCLgni+DAGG
rc5OB+HX4P9RaXQ1hWMRigrsOI+sod4x4vvzrcMZQHT+W0D/13Mi+s21E7U2AWgOR28e7Cpqc3xW
c8Cqy/Ejv1Z4SVqNUIPV3uA7XWjC8xVWVGl3BOKlOFPD6danMX7ZAFsdtcDW/CKLfoh4sONau7Y5
fMFsbjK98p/Nf2rmp5vuJsTTvrHH7TnA7GPjV/XhFhgDluenSHRBE+hI6GH4ONY+SUULwOVnrJDD
zKezewLkWxTXIfyeilpj5lczWfK3o0Ol8wZeSwFYM7NhDWF2O1Eg2QhNg8hdSuqVWU84Wykiv+aJ
qJHfPhNV0ueTUAy5RJRhOsnbO5JKJyp55oyRq6dRLlSrT3SC4SWNExfQVe7WuvHQ+iiT1XzYkjW0
NcltoGPTGfbTlcULMwQqQuyCbRVa1jG8k/8hfr/gkeBX3+PBR3p0go78arAJFepMAbPVrjSKOxYM
KC/E/ZybSPowXL/OxCnycVS0rX6Gx1TyC/m9Sjjs6lq9mkXVEuaRlkiT6Xgq5aB9P3ix0MlbEaqL
v0LXpgn52bXxI8iVZEJV/bAG3OvwcYBq6KXixSgd1Dw3xqRFF6uLvKMhSB/wxSnz+WlWolpYQ5AY
fqWn3+fN/KyWL7YkrZdLp5EAPglc4PlcqPcdD7pBQRpL+4H7Qv9RX3sDAYkYVK8PK+cPMmkuwQSU
ePF5iOMPHq/NQTfuaGyiWVqHE7B7ErADJx/1fjse0uD3d8cW4CjSkXSWbq/NQFaetNuCZig/8o3B
hE6O6Tm3CA3f2Zyqe6jkRNp4xcQ3HWk552ohu9Dpp99DUU0Fq1vrsJ3pbj7oZeox2T/v7pMz5LLf
e/yOOIZfQlUoOEm9P4MszglJd2JtvHyFKCWCtWt2i9CDrkwQJJYj4orktyO4cFg9EIlqDgjrM5Id
wNvUoPSMikfqZguV0Qq9HrfDmCn1orEXuGjDvZnwRI4eZLHz3PO+EOqi3jZ8dYCCcrgpZ0RAaom3
zOlnwEPFVkEa7fahLfTRjwpELI3pQlKMqG15Vjw4/Le8kgJiBQI89vM/jVJ4tBrEeM3XDImVlmtE
HyJ4mTAHAUOZv9gueg5f2Y/mBfCP9fH/emwu6ryQtHGgj+JuuUpWfGzOee147I8g9Buw2pGv1z9S
6E2745U1um6n9zDJEn05y4i8EiOyVG4a4CTk8WhzZLcE0XnT2XflifqCKbfNeqaYtPjyaYd6HcYM
da+f8m5BS+UX6qPTXztgDOH5BMv1Pu+eXDmLgeuT/AE8G5ja0eHEJfkMGKNHd9T0+jbnRr/Ot19l
mNU1clVdwc1EZs0N3hdgR418/b/k1p9JD3TQnpZF73JD5qNcy93XyHC37l4qRzI3n+2qnsBygk3I
k1oPKY8jPyFDIgOarzCRPBYOs7JLEf6DgGDzj/dNMILJ2sAV8nt0WVkrQ4sJ3NznM/Z40j0RoqH0
LzlpleDpXrQN2QG+cxk5CxS8vAgSAJkc82Lf18GERPI9bwvG4its3fcVh6sDp57TMuft2DSiqgl1
IXXROGltVu+oeTHgJjHerKLMVdd+paMgDbqKIIJ4+tNdr1ZoPPzOX6+6737N9XEMpWv2Sr5ni+Rj
Kmxq2ptBfmEbn18iK6B6IZC2hMvFx9oljkaZHP2/QWOZLWsLooiMMePTMjUb2gZ9wCOFnr042ojj
sWxR7e8JTyFISn8aQDomrLxU1don5GBfCNWOBPfhvGyajwaO+OsCNMYBUuJUj2FDWAcbCr2ZCoQI
orTqMHPDRvi75OmtY0e4nYvEJQ1hIv9sCrWMaezqiCAvS2xh4wsXqYpi6HyDWSsktTvFqvVE8eBD
KcZqvECTGBnExBcRc54VZth27+oDCecgeq1aVl17dyUqzUIlzGanfgshYTeTCLlo63LPnRx7a74t
14TX7IXtgAx3+FxSRvNNT1nCKYUa+lmuUBLXyJ/kdzE59ivj88FFMN9uQ50lVHZNQYX+kNzi44tx
kP0AqnVzscgJDdmvJQBsxQ9XA67st4gCzRE0nitzF4JibKk1EQjTewkM3xbiIBKq60UJ1cr1gGab
XhVOTHIrGaJuYE952iC0zaAdUbp0D/YxrfsF9xKsDdGMdIKgoEY7oEWRI7885Lc9f5VGDvoXaIgy
ZuWz6Lo9SX8c13ZnHoQjG5GTn08J+Pkeimr/6A9X1ng+AVTq/eZYyrbBc+n4XPVDhkzO6hwNwZC6
j6RGfwqTe4ya6s9Lk9ovcjy36tF/DuLagK5rad05i5gUb/8Q5TWUlffpvdS6XEeW/+0g+EojoqYh
31FJU8ciA/b1lc5UGYyKlyETA/M9wjQG248z6Q+BWE8GGE9ZxnT98/QacIciQMz7J8QwScUHk1b6
MnNmZBDRsTGsOWJkYF5Hq00npmWb4o1REdDWBZEj3Lk3AhgsjU13Js8+zH/UrZI6RIv/FMPNulT9
QQ/KtuWAeZ+At4vAI8QCnIKgXOQ5CUayZukgwkTX/thXhi2T4/fVJ1F6oP+HNoalexr0qCFslJtD
ZVv2l6TFeyKS2r7QvbMFWaT4getPCFh+jM8Q5EuTNN77CQj5n0WNI3mfAFr6WimADIAH6nW3dG3v
YSjPX53jaU6qRIV9zIAbcTNJKwua8SkQx2k+dGig83iCJ/ZvDGsa4w2t3Iygag8clRVnq7ebWsWp
Dsosa8eOwEPiyroLBq9lRGLvJUYCYqUo6KKNgj2jYyE6kcgMtxZvr+jlRndYvFQur4+XQDHoR0fA
a9xMZDe/CY/q+2i/VNQL/hIoZNFiO3gZu3lFgetvmO3+JdSC+jvyRvbzKTNeaGrcDiDi8Kq5liNm
zNgxiB/hAkz2JmvF8v6/wUhc51exWXQpR9ab1K9JKJo+/H27VbznMiKsqv0395p9CvI6iTQAwOVV
4boNlPcWNAIkAF5EgVI+prmc0XeCnN3PKxyZ3RQGax1LojBm9QfMmuaG5z3TSXstYW/fQmV5LrQ6
jTdqVKkX33N38JX0/ruFcVUH/HZaHEDoPxRr5EXZcbeWn6WL9SVJi4rLiLseZ4xi/jhRhnceUq2q
vbsq444eZg2eRolqySxl3nz8tcNdW4qa7evZIGUeJvZ4Cuf9YlgIDjdefDEU5Dwz/cf14MXDvwEh
u2ZYVarPJujTuzY+FWoQblyhLm/8w7Lb8xS2Jy1cYjZmRz/7Pr+S8aIqspQyUE0VbRdSjFceVcRc
dJ/gGaoVOo7PtRj9S0aqW3OtnM9MfUqe9stvbNC/wj4/V1wcMUSOdftOiTbH4b8Xd7SwssPE20tl
HU9NRg9Yno70u+NikSVsBEvntrEMpZpYRmoge081Kxfvr++aFB95UYg+pJoIXwmwbnJdM7MwL/4p
UjM19L4s5yDp3Zcn40n/SnTSzbfDHZw0+RS62P7+LMj8NwcIzcMahl2iQzFN4O55Gn3uKmOzoBwU
lcdtcJTZkhLiTwJJ+N87bzi6ySMMWnkcNlNL2RTSUBEXJkgWY9KByXazYlGddEmN115YFejIkKv7
KbFg952TG/lbni1LV1tM5q5qW/2q/adUGrSLXFXXT+D9phbd1/Xi8yMe6TEuKhisbIttbhwQ+njA
UmrglSkQpgZsL1ZYxWqo+g0U0b0SCGGFhzaGRkFOcgiCrq/RIZbUmZ/OBqTxrGVyHxlY7xvLnreI
r5hXmU/rG3Jn+3NmeCv2+63fSH9skwtM4yjiic64y2tVx41+h/2rXvAWrbHix+aYWlfGoioyYelM
NechiADS/iEgTRwjcfIpcO1qL/8YzE1j4ctNfnBgTIIZ3oJs4wv5FlJiMJjFw2uZgD2LcOxykhjO
8rFT4OviYEfhGmprpQQNc+zN0tT5Uj7BjyFwcl3kgRrj+u925jc48t7DPhoJJlyxV9Zj31/0XYZz
AIXf9RHP2hdUCJBTypaQrC9T7AS9yonRnqfamT6dLPXb06B3KWYhJ6dcfY3I1bOLUXbhJ+sfZuTd
MJab2SxlvCJ5g7Uu2sqEtt+Rcx9h0riXgIF2/BrBzBhXtyOWSvS0kU2+vHEZshQVqaxYUe8ZCaOf
D+XpePCJk1Mid9Wz2zAVYl4bA2ThXRRcxFQta9OxOYFXKDzaG3gP4ilD1w8oljZuEQFIS0qQwUeE
VRTEBgjSbNQ0YJ9DylGyfmmcIs1vR6a341BXjkFTMt8iW4gB4jPotnQ5MPdXPFQGHIsoON2yL9fW
3qRLJp4QPsknIr9P9y9ziKX0hG+BlWdE/Bq3mcg5b4w5uZX0nkxXebSlgOQijrEeZhrfbwX+PJkz
c1rT9IFoBLw/4FDlDsbQ5bvCgCstH700//OxRCpKtWYOpZ4+H1gfr03RyapC2lK98I8xzKJp81fE
Yijt2cYNHhfDbhf1qJdgT8ihVW0bPi/uKUuvMLnDzPvfCtVUEwHGxKMzL/Nez88Mm9EpQpJndC5X
CI0op9Ice6/zp6ac65a81TloqNzjoPMe+KxpaAiv8DLqomXyRRESehXvK0Rr0ddpJkX29DVIc4oL
AgaEbq3NyWtzQoADkcj7G80BaizTGIajzWO9BOA3643WHtUUWPhr5NANQPHu4NVom0PgYzbDvT6m
If0/5cEMTmrxrh8wJuLw97tEecru+k9hQKNwHsbHoc0cuE+S5MplVMhCS5XEYA61aePV48fljcbM
Ym24DprK8fLpaDgxN2MppHprOao783T6wKKzg6noUDxneIhWiEoKx56N0yg8hDGiUccEuiSgw5sk
BQUHUs+fUl/EXl/ApveUaTTaK9sDe04HOA/8HT3MCv9yHiM5ZqjT/ugrkXy2+NOeBBVWFywa0zJK
N2ojiObRZOvozX2EoMva/fbBwm3c7dW2/uj1U12LjabaKPe3d1VjHTb4gzRxY333FK1Ff4t2jf6A
gH5Ih4K6dPCrICy7uwYk31eyyGsopz8lYxdkgqMqKd31KKyCTJN9oL+sdOXwy1VzdURiIrrsiawg
PIQX/znt3mzrO1Brmwv08P17zUCEJNkyXPY6fHRA9GsXS5w8hk3IGpHEQ+KH6kMNCWpQwnZbdtmy
kGSzYsZlFFq5SZnWiUCfJWwTm1nwAK+nYjGs4RuuCfTaYGHMpxOcmxEZv39NogjK9IEkbMRqRTZC
pTC68okHVGQFsi6v28xNOzsLkKVOQtQ6QqWjC4cw5/d3KtyjWGl2PZa9cBeWWHmMijKBebUsHpux
rQzlONAK5X4jHuocj1V2KF996U2yHoWbFH/pLNsucfETcbT4UT2f7YNIzBjh83SVStCqqNeVihVE
cbVd1F0SqCTtE+Quwdu0savqDhO2pRXY069r/tTbvOqtO+eU35TkcQWXGxvYEL1jTj1dlIb4Agnz
AL6cmhfQ+Pe4EROVX/+h37e2E+o50Fq9oRFkqKTKg/Egj3THdzfRJMO8AYIQfyxK/z2jb6f0RkUX
9OI/PGNI1qSWCkkaX5Rnwp9INwruyVZZmrwMY8yEjAHSvxmCDZNIs2VFnQPhm6iS8IPgbea3HhfH
e1N1EshCjvN9stFxfahUikO2DRMWgXR/fj9iU9LMIP3X1jjuqr6qlZm9+fb5AUI3XS+EV4DSDzfa
hEGRaOj6P0ZsaZARioOQT7kwnY0TG2M+r3W76irywThKlDQ0kR8UYktu3XDt/EERDqpGg+oGDnZS
v2B+GmTTD9BfYMto6yDKQ1LBiBdROe52XcAWrDTR401I03DsVPt+4Ds1DNaEG9pdJ1yPihDKfOY+
cKSpxavY0dYSES2/Ai/8KlwdZhbNdfkqJ2jhIOU8n8g7P8aG7K2CGdQDsy0w/Jbm0ffSgAXuhX6y
b+RWaWxhnzXO2bMmQSMGkkpEuOKCo2TlWdByJuBtMeY/EX/Ze4PBPL46kk7K28ibf1MAk7+WjBMh
+XMDJnnY5MZvM13WiVE8II7nllqAV6TeapYv4v8EWWqsIJIokMv/G6dFlkDn3WevfpxX5YB1ixd1
zF9WjPvSWcqH4r9S22JLIlgAUildSlSM6KoDfrbmPshtPA7ZYwaGSlwfkIsWGOAclFFlz7uuUZL0
Kjo5nyaYiUVTxqSZqD4TrzbgtjPFDUD7yP9eCLTWdQTHJ1PeYUBRrcgImKX5gHslwHjtn0Ky/45+
4H5FxAeyQ8XyFtM7mTkHeyHnOjmvKB0XcJKkhd1744514sd2SWaJZYFMo7MmQRivJ9oJCAUMIHQc
5JFeh5DsNtC3RIlB3LaQz7ynh8/LVrRuWq4us4MkT9j5+N0S5HttIfOw78CGU1nGpkLWoMNs9pLA
BbaaZZFmBR0ySNmYFGaJPCVgg1rm8TdAqTXAAJP+QfZ8o0fRBviyZp7ougW1r3JZpmnsI/NO+fxM
nSoa4z8Ki0NT+kpZLQPqL9N7dmhaQksCfhi0j06BaB4+ehe4ogZHwyzKNDKxF8FLyHPVitegNCEd
dK457Q2kaVvaOq2U7qDj4sxC4PL9NTFyTBWEc2p21tUZaymSK/R5mY5OYAZVxMd0twU3vsjtN4/H
2dHkZALijjGIbxQsy6q3EoxtnGMjmrQVgatCeBvoDhx1D6AYZQujf1MiNbUyKFaWrmscn2+NO8KX
uTBXx5RHd2JcS3AY0sq3XL2btnJzwEM9pg2S5jo5sP1JogdEQg0VKCI6qOxz0HwQSU3H3j3Z0Nha
Rir5tW7cMt2pQC6o6pQihfdwb8jh7VF6qItzQZknxJElBnUgDIk+RWt7z29u9CILKxywJKX6dY3J
oQqsU2yhwPAIUTXrdoqYjLCA7RgRI0KLfiiTH3Tj6Q5DaqZSaExltR0yFPmitKSt5juafxBfzkJ5
1atdn1bMlkrjOAORIs1AWd/dIGwVrDp+ennLw2NROy9Zus1Ocsm0Tvin3ip7OkRZ+XaxpW1jOSD0
S6WOI0nkszi8blBrStOBLC5dQT1OZb8KlGquadTOIPAWG6gWyDl+kFM3cpF6fljnUyvGanoLJ0PS
byfkYcHEvJkTPeKL9n/02OoZq/PZC/99+NlTNqpjsqTvmODiKcB13YjDDSgc7QGBGI8nMPaLEW5+
ec96EhLCjGHb8s3rSuXBGH5G/Sv4JXC8YaVIKvcM9Go8V+cgr+z99nqqpp/URvE6tGO+Jg8NkjYl
wiGpmCrIzEBDZbvZymL2pS3aHE+395CW1FyyROn968UEumEmWjdVu7HmBTzJVm7iQMamK26zWiCG
qGWtEz9lAFVIFPBr1tHJCIwJRB+y4h9SAvwCxJ370aoVs8bXhUNTaEhuEVGArOqbrkoyiHYLYnTk
cFsU1XltzleBr183AaX76Q06UqAikYWgPokfGmCYQs8fI/WX5kdn2EW4IkWbwaz/n404IBNZ/Wgq
HLAhKTH/hjqb1JxC7p16Xr6K+ASGHP+XbZPd5fZR2TDMH6nRfdOYIXx+dzdoVdMN4dfYdoQhWIjD
8xd2OoImEr1wDV506KaoFQ5a1iHk+a5ELT5Br3PjtjLHfKCtZRA4GkA93xD56AtBXDRzZzrUbWZC
uydQiFsb8gaOTj2pvh3DJ3G94TQMHOAAosKbqyS7X+M7FAE+VpvIFU9k3ofsIpSh2y5pWOEpNM4T
v4ftqRrBUis+KoQTp97SLolJtgFDyj3ho4proRvsNozGlqPBWo6ZUMQJxLQ0XyuCuAyzQ3lvgD4o
oECt4haadJJ4un8dyoJupFk47nGbGLjWIPXek7mjX54XJpiQoVnvU1tXTyCaf4v5seog+0hJ/JY9
zp9QmSS8+GDQeyMVFg1MO134YkQ4T4tbBfWgaQaXG/HZch6EGFd1YdrcjFIgK7dx9Vp9QkZaFKsp
MNZ7RPP3T0WADz1+Q5x1D47WqfQCMW7RQLrtRQdP3/IQLl7ZGv9T273Tpb1B7dmKjMetdWhtqAIA
+/2IyHicyQrrXuBAMdcGlrZVMrjhbD16sru4rZ6LA3WO3EgIzlghZWL04SGCbrEGrd/yLof2QgJz
ps0supgtvv94xRu+RCkOluwydygFBQwTDZWjjWzJ3zbEHgp7QY4UUCAwSlhoFS9FAQzaNSsX5lAT
ZGEA78pqyC8imtBjmRC0NhGLvKZwF2iA9rBTDuRiTFYmj9DOUh16MujwfOxQVh70uiEa8Kq+T6B7
BBTjWRis3wzAaDPjZEpBaZO6aLuP2AmLy1ZFIo+Yk1ErcyLpcAVoJ4ODPD3p/sd+Qmqjny6mjken
Ke8HD5vTzzJ/ffjuy12134Jkr0Y1gy8zpiEsKkb7C6EwOzw7itpAtLp5wtvs2Um4GsO66GQIZjl1
IOYadVcLMIs8OhB6GygOxmWffUSqMe1wM4nRyp5ErMc6EhZ6xGNPFT/CwdRAhiIBDLwAHtbLgIfS
bsZBtbh74ioC+3aU4WR74xeM9EJ7bRVzxgKmBZkavvJI9s7qQfDjSArjumbVsWCpCtsdgqXHzEwu
9tfJGcvtsHDMU6IL/Y2sOCGP2kCmTxJayriFyeOGPiTPpyAsw5pY36equ31k/r+d09UkbO9fG7XV
LK7wLqlLe4R75wP0Lpr6ut18ZvNKGKsujoZkBPHqI2tieVWjk/dsBYsSIRG4jjtWrYpDoJVHcVqu
g1dfd5tFgWGALy7wiX4AGxAnizEG5bjVklRFnJd/LBY2qPRS1MXb82c4ybBpNCTNL/ZZ8Y4I7Pyf
k8TuPPJo8LBt6nAY49C3X+N6TGCWELqaWWBc/s7WLGffv8VpxCTp9aEAPAhKxYz2rreJotlK742O
WS71a1RQ+w9GgxHGyry5q5BTzj7lKTDGW9Yo+trBsXbcj4bxuEPQRF18vI9rUhBMDRKj1Pl01oMx
1ovPGe4lrpAyBZt7wEWF1U1jVPQcpYnffaD1ttygIwJoohVskIJD6rVuR3BS8ImSouuJsbkeK3zF
M/dS7XXi+06Hq/SMTH6pAfQPqlAQQ+yoEWUuVLzdlv0H5sCdIq6R5xTN+V6Z1+FV2/iSqsyaxsAW
M3NuJvI1KtAXQQcz2IAeFZ4SiD3IUzoHrSn8EraVVvMVU+jplJRz888Y2w5732PWUPp63GAREbqg
/BSgJ4i5yqBorpg2we/vmlQAYHKf/hNFLJb9o5U5icUtobXlH99npwGVZEIB0HUKCAblWP53ojKz
OTZNW+PDJjoGAboy39vCoJqLw9MBT8CGX7b0U9U5t9Av632VLmV1q+2yVhYle0Wg+EYV3agYesVI
fNr3701ACWx2OOa1ArpztZG+zQmpuXDPIMkQtLRQWYKS9helXUFyTVzbA+6e/LDqtuws7n1LB0bB
fHtdkkzdqUr6fNwIci9mJttLnvlsOGzmzeJe3S2TaLwa6k9oG+3Mfi1hRqdJEKM3k1KBER4I6+Ca
DSmQsJDGwoxl2D6rNKj/uzCoD7+1tQSz1x8/kZDT+p5suLa984fswV1v8QcL0ybUH68Q9wIeEV8Y
YONw7INYdOnCmMpshcpJpPAA1FLMG3I+Z6YUeaG6jC5/b26HCErhmJldMMXA3zvZZ974rLSnuTFE
5JU6siXy/5q04StRaLEkyRlZvA//fDvHW+n7QqyTgOlr5LGpa5s2WksIAYrw10uTe4SivYsUbIuV
eAqIkDch38IECHV5W5AK9cihYKZ+iSN3/ESZD+Kk4I0IEVUAFysvDU5TGwN2seoc4HIgG5npjkHe
lBI++R0OH+hX9/CG9aCa86+1epYeUKIbJMNpz0j0coQAxpXgwtohQZ1iml7i35k7Hu0cRIeMyfg1
M7AOwC69L9HZXKSqYU7X1w6U5D3cx8J0nzBo8+9UklaSo+lNlF55FokjQHy6LxLcBa1wjBNlc//r
xSrmSY9cnUsWqX7P8vgZw10GGLxjjzSdEAOPiFGNPlPqvduFdWrwksczfVzjTDPpibWHV/zUAS4w
LZj9SIs6MzwyFt4U2qm8tPvYc/cs2lSnEWDXuYQHLeaP9r0mwqWs4y3MR6ncLgyul8gKMygFpYHt
gDHeuJvN7EwkW8SsegKfT/nO5chT4kwz5V/n9XaE7+d4163CJqdnVtsxfsCYzc6RHfPzZbmIC29J
U9VlSYlMGmA6cmKbyA4jy5hahWRKKI1RV5zmv2onFX1I4JAs+FShX9j0DuwFMMQEEuUIt7a6fKEK
1Wb/grW++Vi9F/6ie+KkAOeDdvSXAwZA4CvR7tyq24AZAReklOBpRil3vhiccaZIwY6P38N2v2NS
WUIONJbbJGkhRauWuHQ5IoTMQRmDWVMLb//9NaNYl/2MpLbm4X6Zd0udtCKM9fnHFdf9w8ueo0v6
7vNDbw69DKNQDyOERXgn/xbol1ARJTYQGkFIPuW829njO5cNxFcttrQL3HuNBpw6XqQpQaH1SoSq
zCdltTmZHhwLjUq7RX4UJ7LOmeajjtgjF+dC1z8WK+OzrIs8mqmBwhynE8RBIMJ/W5WBiZOPO+vc
bHXyhQgwW7uK4E+kEPTpZWuUe9UulFYrPb8i4rZBnNw59en/26YiYkIjG3Scx96iM52s1idffP4v
tmyG0r+Dg5CRMG9hvdnH/cBmSa/+ei8Z2Lh3CIs/rFAm+0GiO7QzEMnd+9XHjE09zHj06UBuD8Or
9k25IcQA64A4R0X7xTSOcJ269qpG/8QI3lzfolBBInJfkyJ40b4o6bXTgOo4ETNzOTVTR5jWYcVC
krvqLTEAA1UZrALyZzEYk9r0Cqh5RVptR12lHaXv9U34Rxre4TKI2Qyt2l/3KDUEMMAUMZg7sj08
Z0FmdJtte4Ld1IxsnVB6UwGAXXm6/B8psmOsF+k992A6/GjHerLsnzgDysQsJwISN6WyrVGC1/mV
bT3kqQjiscsACxEwNjsy7jaqP4LhO/wfIHpqSZgl2cHRmy4QRAkfqPWLanOJkZmj8EoX1qHFm9Cj
N0iyF77xbxCnud33gcQbisTy4RxPMrlLIJ+Y+jDf+Lt8SuQ+P2Iy6WPrwBiXmkFT/roxeeBwcRhk
OlLVQFfQ5o5Vipkb5gyhR8gVME+2xaWfOluagPXqrdcW25XtjpxmBU6atFnegVlYYYR2eATrS8Yv
bbAp5glHPOz4zII8B3dqr8VGxW1u3pokafxOrQKWrJLWOO4BZhuyK98q9KhiU/SSAR6trO3QXj72
sP0cLwKS43Wb9nNXBHlzr37xxnH9Lo60Vtkq1PaoX7iXJ/jxoD5mSyODcbjWau1A8aGakPMpq+dw
5uPmQkVYTVegTyVdbTsNkzTrs3HM/6vzpojDxlmnUlCqh8fSH7Y6EpJcAZQ/D0PtFbrWJyCEU/Bz
DD2Em9z5c07xdAWfic+b6ZdEID4Qdq40k3AckSZ3FZJl4GSotUCfvF3Q4ZUvmA6qAsJTGFPtQiS0
S4HRZhRPoCy76izIrPWZLn6stXsrC08Z8KCo5I0NoZruogegIsyVqSE9pPb3i0KAp437blo25KyC
npNhPaUgw0WUzhnEwYpb1mZaQRpO75MQ4R+g96QOhGGupG1i9NyhPLDVExUxVPXOrVrWM58Tk0p3
yekxxFFtqTXTcqfsW9xicSB9ZpqaMNxqLylZ+H9TrbvyRZMPBoZXucOu1cyNxdjK/AlsT+ULdmIH
i8hY2mHB4+lG4SAVSaUH5P/dA1mKxW3O3WSlGfULo3t4vWVOslIj4KStIiXdn6+WwQdw3AtWWQVp
bQhbiZ9Ng2zEH19nPABd+NYJTNh7DpH7cx4IypSc43bcgDP7IQ5xjtwROyQzxhSgOOUzIOP+oiwr
QG8KhUPtTziciG9nQuOICJmuHqIuftvCMd4zL56/FvNoGBwvF6Tjlkz0b5EFWqDA7mbdGzBtbeGh
e3EpRD3wVYndbF5tOsn2Z1JtiA1RuWHn6EjgcGOCPN63cbWwtCzie91HndiQoHo4gAa/Xu7g6S5d
PbUC+WJaph7lqakpTuQb6TJTGUnvEQMVhKJHGrOPt40Z0qFoivpWEZptUyE6KEAqAexVhCkhc7Fr
ODz3rHeSO6H87qI5v+P80YYEct3DIi8cgDnND40trkRLS0Nx7L7xPzmayo8FWXeZEVg8VeIgZzLl
+catRmrciAnjhs8MD+6cEWipXIhc9v63n+GSPAuLODRMsZGJbeqCzs8zHOfb4F6+R/VFse4JD7BF
zcY2b7k5aYQrVm2lJhUi5cDovnoVcGk5Dca5LJmorkmGtspMg1KtFL7yaR3301LQ3RA4PJX7MtX8
L4bAwEt1LyqopeOYT46QFo5DmWEtyEAYK9SyFvpLsKN7sAX+c6cuCXHBFv4YSczT+RHBnyF4hzqL
HOzBCZumExioBWEM+8lH1Yhj4XhsP5Nx++CCs8+GvzSMfg8RKKjuoF1w7xNevt4d5rlV12xxo75h
Kcp2t2nvJzeeavhQHOznIrasKvMwPGj3b6tVRcXGbN4axWp9/WvXJBFmF00H5O2hW5L7rGrS6fIf
1GAzK0ZV0iXRXstSnu+sYUqSgKpW8+yhTpINXOQPulkX64RUL2yhCBVC10jVqnltregRPck+Z9Yj
l+drurUq1p44IYCBw8qEFGVwAiUaFLC71HSlk7HZOyK6JZz3YSaA5RdotRjHWAYFG8MI75O+pmji
aY/fLZA948lXS1xipsS0yST0AhZ3YTm+1ghnMLjuZocdVCrhRtfUmj9wZEnXpgwTVQuHzFLtaKyN
2Ut+1gQnyMvrKb6h4V2em9MwY+O9gQ3lRK+g4aVw+jDZ9GXlRyQPHj+5WMTTixzxQcnnA55jETyc
4o4Ldz5Naii35cE/H3m5mjRhRoalphE7dXNNatssU2UZFjhv003ga2GWpliSoiu3Ho/BWfoHb9A+
CEVlaD58OiDPEMcdXTDzmdzuRhkfxq/ugtADN92NBqkcQtuDOud2p1+0D+UabKgIEGQRn3x5pglW
NR4ym52QFtHYfCm8Lo4D4RsFGgZD4jzi8fXcbuxQwKScuEjVFZznOdG64aSFg/BfDK0zBGmu35gL
t+rm9J5I6m3fJ+UI0rzFfVLzqW30nJpoplS6dLvICcr+bKhICpn6BohsZDazwav+IVTIOfing6Vz
ixduEmhmE8GXGBLv11tmV2is2V33eSVtGDo9+TgNbPHzG58v8LnZtvBRh+dChmaCm8esc/SufxQ8
eDnjrhv/3V2NYafcN0Kcjv3/yxhTvCwkkFRm+6NG+vDhNvGn77vlZtIl50mherOP63CFaCJYNkZW
e73lHYkQwzrdRsNTQFvdy0EoPsJOxr3lVoBbGiOXCa/JoEKaNWFPREUbsADDmP/g0ENOpGiqjmPU
RObInPkhin6XH0P0XPQSYjlDOzohqem9lWa2xnOOyGkVhFcHyST9zu65kF4Ouh3KOXmX5m37AdFI
SiMxT98w72ZPLHvmWjJoJaGkir+vKuv++F6Hu5EukA386G1AikS/+wnX7EPMkY9JHwwQkgLxvAg1
LxKdhoSnRQTXYgwHjFR6pSVhlZPTrPAAsSdJCg2OeowpfWJx60kE3t6AxPw57LBhHuvIB0bcib3e
983T3Ct38v9uCd2w6CgGb0GShIRpEGTa8DV5mpXPn7Kn8nG3En/8wYuz8Bvme9q/6Rp5lKDFE680
gTURuDxxYT4Ol/aBtK2zWpuTwL7qMRXk1oej4wpI6DdfQx5wdJF3KKAFLSPLlTLyYn6TPXTG9MzH
jacEr/RMaBK6i1FtsLhN/WoMbNqo/UFfY6pk2NuE4hpk8OAd/FaGQC8jhE0P08Y3Q8lylgHKTFEB
L6CNnRhzT09hUSGu7ZCNsFa5QvdoYjC/zf8NVCjqytKGWIXpdTXXBJhSkh+zx+phIdCRgKf3nwoW
BnxwhQb3b7Zt6QdmsxWe6jzU4KpaZX8JPxLr5lGo5AzNF4a1Bux2kGBK8Y6t1bptDclIe93svuso
MBLSx1nLMDBBbS4rsdLRKAxknKWI5QRK963CANK26e11rS0s9Rk0PoOUl/NHtPb9K6lI/eGVpnM4
HmO7RN6MGQ34HTgYwEFvIpNoAdoFAKOrmGfTmwsUIvS+sSg7RMpcLAMgnVx/Ao+ZMnEiDsVD6jWo
at+R+csJP2ZDh8jiDSnarIWrECmQ6HYZ9AIVttfHHDhJbRf199qG15560XsgZUaxHKDalT0TLrS8
uDYsg+HnoudieG2wmFNJmWzgp5QGzZhzrU9rcob81qJ3uaFgb3JAm+6lIs5jot8qxnpJRhb6uGG2
rKs0OTBq9gAfJROyMwyMLIrqx42zfkd25t0jvW4fdjRA894Ecw7vqY5CgWyAEwlv9hZwL6Tmb38d
V1Nu/OpLX24f5BzKl2+fiy/KQsWpwmUL78gMiXlTN/bNkSe39Cq9d3BQzf9eTo8gKf56SO26uyYe
a/Z6a9bbaB+G5z2PDU0ysBnjtUJnROD5dtDv6ZJk1WzEZ/wuA1rEdxIccVpl0DQpU39/LmacemTe
KvhJgGXnZWN3nFxkWFwLizqDWxTusC4qPnb5Gp1sE/+jI8LM6dwkdjQadorhoKkAlZnRDL/ehNiS
Yg2ub02PBBTeuJNrPg8hMQ8IhMUyK54ULZI0BlMA+3crO8vg17qFN6JlMsy1KpAzm8XcXdTkujs5
EiQRQdczU0VCSvZETmbQjceZtWqh+qs5GYCfWKyJCC5Dcx9S9xIrqpAkpnjxBS6QV8ynvxbmep98
RF73bsQ69UsBt9WzvWcw385qZiioXPlu3RrobDMWVBrdDfkx8fb6Wy+a3OM8ScMNURzwrzfHRSf7
PWTKORSsxMt/cIJDa6qddA55u9DF7EZqLfn2IzxftBQ43FAeD5KxvOFIzyh7qYCSsUQr8/2mKB8Q
VWOmN2bj/+pYLC1y/ouL2TFxV7qKYrI+/DbvgdEySKjZa0qENz0IFRPvPJz41O6CpCg/EssrZUsu
rpgM1PuPezDrJN2ardYpe1CbQYK3FUqp34KA+0CIcOApcNhqN43Hsa1BlKK6PpIt0aOimWyS8LYg
ax5l8BXoeD4yOrN/ahfNfat4exXdOPdSxU0xoTrDvFbN4ift2RTvejoUZukLn4D4ofNfAXDpCMaj
ldZ4PiKGT7IuKgG0cRO6MiDTUiOEaHoGn7qpJCpRDf6Da/dYeksLXx381PDiFvnFrc9WVbwg0ylS
+VbNJiVSQ9d4IOR4gA+Lk6fbDbL0fBmz9sRRWDgpj3N5uN1kHKsvNRnyBTKP9tjIs/Z2sMYZy3cw
uQ/M4uG3wtX/Qjc2YnSqq64Za9pAaxXg0O8T8MMikQEiqLPkptGisi26FQv6BXbhlUMpu6Osj4lG
1lLdyP+K7KtpoHeLbzdDQqysbSFaIZ+SMpX0q3kN0Me60st6e+OSrXRjYFPBhoZ9Sj6hx6bu2Ss+
vxD7Bi24yGEiWMohtLfGVXGn/S4H80DrvWnMLHWLbG5maImN4Z5ApnlcfywIpVfIGCGTyyezYJGU
Uj4rQWNGE02QKh4oY6PwHsflDFW9E39crzkemFclHq0V+YFIcut4X5+cAPmPJyUaZtQo6QW18SdB
QilIonWcVUk6HyKaYvWXDNCtDZsvTLZoqJXFvm8PMhAaFAijhwWmVC1+JAffyPPcGfTwDYWVt2ud
2os8RGx2mM9LYNNUkfjxX5V4MEUlI8OKQqs4ylOqtab0vtJmbCpdUx6vXPppL2BdT/HVCBLVurzg
PtzYJP+Dog1uggn7agdHHyR1Ucqu7fGYb/CUstpxuCnA2B5iJ0OGI014Kq85JIe/SgFJ8X6r4X9/
tA/WCjOVWmm+RLFiKDXi7z9dtBAZ39Kyy4MM5s/mkMG5Z6+YqZNIzzkUceivnil7L64/sigxxo4c
Vl1sY+msnTXSTc/wCCNg8sdmgbPtEDTEJa0PhvdHzj78lPPMDfwyWr2SFQX3+E4uZjOXe6f6o4zY
WM4vIhaoLZ9AW4dgE87XCwK/adDOEUFy9LhRfrCrqwxUDTsSkqYeDIFPmFLykHVdmqpLYCCnoRL6
xZhPaUWLzDlgZNkfVfv+mIT3xiLqgjCnjsuH2zN1YGIL/53BNLAbIdBaX6qDotDFLTsXSsWjWGiV
63KWZT0XjlvxBQzD6cUGbM8AkGCFY//3cmBkcmfb5TqR0LLzK+oXvJxYnNRb7qViAqHGkKGe0Oaa
hxRSDI5DPmriBuG/CRnttZEpPE+qXJw0RiVKj4pL3P2mc3dqfu+svHiES6f9CWn7kfdOwJnTjz+I
f7+q7xv1pUK+/HP/JCS0ktjLJ17SvMiDR5Z7JSvYNDQ00jCMcm2XMOVPeALC9u4kcUHlwrvSHKph
be55U4FZ1FZC6WaZriesRRxmCD5ummSlBWcr12IDVIHI+oc+e36nyJcqrgzBw4268iX8JjnOYVhN
VW7ZfYtf/dac1AF3T2C/BRXpEGrp6OIuouNiHUJkhCveDpWvxtUODEwbsvPFipxW+3kLhx+Vo4dK
ZYMg+PvywqTccpxUyYF/vlDlXKjDHuF8hZqtv2SFHUmgmSi8BbMYkTkUuLW4GtjaXIa0V8+UPczd
+eEnncb+MGuvd35w7E49bzLTT/NLY34pQ8RRpjnZ+dmV9qgRXS8XD1Kc+YHDCr2bLchwi2z7wbs0
s2F6rfpLR0sjdECevuWBDdvLk0fb8W3uD69w2apr6coRVmRXTue6OQiAogBZuyasFb8GUNOY1Hrj
RNj109OBKlhTOuKNpH0J5/89Ps/szlMsTPiAIPm3Kv9wpmujHRrRvYeD5UDlGQq21H5ifV8h487g
gR6MmQrWaqQItlz8jYPzpyt8kgk80qDktSS0mENQPdu2DM9lGfebmGsjE7xRCbDXlVka+PFSDp/w
1JNPhtzpV6cC/yMueQbtJTpuLe/zPCb6TODepZalH2uirmT/Gev7r1OM4MPN44uWN5gmKiwZ6/jT
aMVxcuH9/tHHXpQoX+BrPCvk33eAwSl1CVKITgGHv8+ao64CevjtFUbK1tqX36SkJji/OofAuacG
MrrhyrvaWm0hMrlGHFE9ljZ+eCcxBE0XsZZpaVmi9KmLF0oNJMDadzcdx+85hQOrEhMMQwGFdlE0
SfnrZ8BzbfZy7EUQ6gU2VNUiidUaHXIEDdqZjowa5FR8IQ7xzbCHhB7DW7kXUtOYNATfVpKsqUTi
cokyM//5RBGXyCP6mvtq+t13R/izFQkmc0QNlgquWnbBbWN/Ocfhn4DpiA9VgRnzA7l9WOfZPDB7
rLcsHSDAFgdFeLMIS1uBaezcoySByLgUD3XOAdUlZFAyxcSW06dKx9/lsidTYxt4T8tdSVHTbvxB
80/31wsAgEnmKnEL3TrtwK8LoXfSD53C/70V8kvpAb4Mh0AvOg3t6mCi5vl5xsabQeqsQMHyqc2b
iCVBLxGs+1WBRO9u3RIfHduStmg76OJgGWDd8BlQlDCTtGULgPPpz96TJIHTuJozjccXdMr1H0W+
1V41N/HGvnq0Lx1nBzu3YwfZwFubsIavDU+onSa/5O73nst4/wz9ZWRbnO2tKKCNLi4wyw5Dp1lu
0P8x0/9+CstG+eD7ZrMKmSs0D4HBXQVaEH4A4vXRSFcb7tAsvvlJpJiMwEpYDYD2BL/76X7VQspn
uVgU8cLWdrQHqs9w5+YQDkBDiEAtVgSpvxN8ReRzjuEDJM/Frq3dKLsZbPDzFmPs5T910Y00NRul
RWu8Dj3aO5uy0/ZY7FsZ7fBzuRjkqglXar4hN18x6VfZj8bWYnCsGSP2h/Rr1Ht71jwLlF4/z91X
eRayjuW5arOcPcg56YEp8SeA8+AEgTkk36fIciujD5W5ik/bCc8+oWv3+W7qQS1RcikYameGvjTb
SxtnnrkQzQDvd4V1BMjUtgtYwuLtrorGcEkLs6C9OJse11Ml9psuvAFOXZIk1V/NrXyEgu0uz306
BULJ3TohDCOec0nZ4Zy0B0/0tVgQNI4dT3DAlJKiASurOKlxFlb3URSPijHRcLjdF9vp4UbHvL5i
uFG5VPThMCwp19R1vYOISRcSAMRRjyAARCNFjlF4KNU2EUIgZTQqwdyzULQQrcQ9XlBiCUz+t9/l
podwuYImqxZfbJPqZUkUccdTbHg2x19DXy+GfCmsZrY2pr2stUFh+Mn5vUQWwThTp7qiGmFB6YER
+OcrlLdFWVqrph9Avrm7zyQkijMTsr29v6/grWMVPuP2WMMEdkhLT0iogXtvh7E42Bv5XeSQ9Dd7
v7BUXc2x9IIeoFrW3kLWbsk8ByL7D+HeQ/E0V2W8EhJlNT+i5NKp0MnEaDvkEq1wIJVHRFms3rc0
9KOg3NhJAuw3l9bRZFbWjowv50xg5Bspi0bjHS3VogyV7JNp0EFkrgHIlv+8MtJrBErmkJ28d2Fk
CPXnUF+FD4lgOSESlU1N5r4NqVYJH8AJ0aTpkrW/duT3seoaxKAGEv+yEnQ4s37VQE1R/fWvwzLV
Ft8cMmQOoroH0bfKYW3EOujo0C6rbYi8TWPIaclQXWB5tEIYA0fS6QBn0biz4mZXI5eRDEaJ9rNj
Cfp5I2frDCe3T1iRF4SYbYIcbG6zzaMbUYm9AxZOdVCb8aOewHXTHxauiX0kOCfZuq9uOdZKEdkE
Dl2Cv9hHlneez5ERxIovJU+8Qu5oCogZuYJA6C+N69tddxMa33GnHzPDpVTR9mslMniR/uY/Bazn
GkHqgxGOJaBUHLNRFLsNDEvNojdD2w94iHB3NG26IwXHrFpy3sr4uBYOZKqTBPFU9dtyETRE+p82
TwT3LCRqhF7GtzxHNoWf1jWGRjITsJ7Gvab86yCQi55rZ+2hO9d0F9XYFad+lO5DfY0YiMfiYG72
lEopoOANzgTfe19zPSrONljujxgYfWXBGYSzHr+bG2QGTHPUb9j4jsXedWyYHqp4ChAgo62DMFJn
XFtl4wTyFZoW3tNtU1OFVxIa1B0Jon48/b/PUf8Rta6m82B2H9dmTdWnhuH8yggiqxzSBYroPrEl
5ZyuXnO2o0C3dAcIEnhiDCoR8F3Gip2V1Va+tLOEbcFNi5uxL9/EvJTLdtBKd1qPhTEq2niG9P2w
ecl4QErgVI/47fR1z1DohSFzv00H4iQreqZdNPL93Ob/ezh9uwTRDD90bl71cnx2kUnFyJ7VtXlM
SLaH0hkG9hXLjiGjAFIUSgwtXeAY9gWXKAV0Ou1cqGxNMM9cpcqiMLbBgxrSygcRjQb7pq9KSCrS
vtlZh5gKvgeIEv9j6CfuxApvxhdqNUWHhaFWchJFLd9APJwEwSPZk+xXbAv2QUpUxhTYe/V7ME4D
hcVsZajoH7dsXnXrIX9clUYVuck4Mu+uM7cec80tNos1K3Eq9t9GLDo4dH2nVryJ2jKlGnDpDr4A
6nXJ5RRm5aqZFT+/GiIFUFQk2eXukkXtJfuSK7nOB05UcTLYf8CXWvZVk5+qCIY/r1neY7QS2wuu
h7UOO65SB62EUdO3GJXN03wUwpx/gXNqy3aBoGNJSvbct8cn2hwiQg1+nAtB52PzaNd5t1D9Ja9q
jde9yElDfaXTVYhVbMtOgdXz1DgzpJ3FhWLD7hPwkAvnUnV82lGamuFppMp8CpGYs9pkbDfLgUO9
gjNRR3XtMc1m1W1K9qLB7MaU9whCcnWbHxoo7ixcFHlLHwFLmexGFHjy1mi/Yc+Eb5AHGSvdjwr/
Jnvom4aa8GWo9RY/Owc9tC8VPV16qRhgISrQ3rIVuzoo66omMygv16p257ZUYVeMruhzbGm/pWAZ
PJaWffdhTVpBaW1zCO9FCzbNYpesAnrhlgTedZMkkIwcNFk8FbToNg3q3PrKacTzd2sUFuNk55On
1sXeeqt2h0RRI1622xlfSJqKwQ1VVhlVq7vFJ27F3mU4DU+EMQLFOubDgBiMskCj4A+hOf1iaO1l
EYZg+kDJyUvQbZs3RRhIPLqWp1591LozZkJ3sTn0S9tqwCgg+ak7Dv0J1x/O2Wi0fWZhDKgOyWpo
ZppXeWdD2DuazpmNJRIHKM37U8Lj7WSU2YcV5BPywjqaq0Wz1369H9VZkxFx9asGoMZHvMZPparI
0xa3nU7y826Y6eT0mLlwaO1fuyqjfnrlSRaaMfDS/8iSByWP0CSQnoDcW63/616ZJmbDEScM+XMG
KQuyipIeZiVSmM5aJsW/veBtk15vylrQWftWsjLfhfuPBH6aWUdC6/uw5zWTx22b7M29GganKa8Z
++GFa/DvKzkj/g3AjkWv8rXrGjASrI+NSO+X2XljfxdWPK2zg8qCuw8ZwAdZ/0q2RfnW+edyABxc
sGFVfpbQFg9kH+k/Ub04xuXk/XaCzKsf6XAQ0tT7VBUtOCWmSVHfn5hCbpHK5NdXryQZwv22F8vu
WoyDYZqUUxUAn2HVY/GKy9wMsJCW+lOobigzYAWP2o2VpaP5hWN64r48+oPUWu/lkVvxg7XvAApE
NOLf4ZxGgPiOUOgwC3Nzdud3F/q1wqNtRbTnuq386XzhklLkHnQqyfsh1jl64NKDA1RxjAt/6f9G
ClhplHxhdCNOH8qQzbOAGysT+OOBGBc/Z/siwTUxjdZgWidcXEJJG3rJZls6UW4r9ZmaIsYo+jpa
A1xVTcTIOmm78JDwKVBpS+aKpjSqGzOtcq/IjLa5CCTvXKf6AlByaVvCm3ydMjeTdlz4126LP8wz
Ku1CiY+36x5rAeH5eXYcuO1JIMFilmh4BwZ+bvLu54mIguL2pF/+Oa88xNrCUnpNjT4LHR5rPGuk
uwd3r9dMfkKGAyDHONuTaaZdZp02/+3lQA4u+EpumP6qTe7qoUqhlnJncFFwTUtUB3TG2soZDMt9
2DgLxazcQWlsiyeLy5V4IbsjfzSGLx2EjzE8RK0gNtWD2iFFDlR1JPiTdiZV/KS0cKEWWF0+yYaA
7729u1dUEuvk3CtNZJZIj3ekoJZ3DsU4tujezQ+YHXgbt0//HWyumHW9naxckG7YYTpK5P4j/dZY
/Nsm93vzn7p6VXQGCZR14aeXfVH3gCOu89LLDxkRlcSHoAOEM9u25Ge+OpHcP69JMEwoK/ZN3PfB
PrfayHDzneHiL3XFCKqlzrRqpiZQielX2coKwRF3Yl98EfL9erTWXwfk6dUzOVoFuz2Smz5emHJ4
pw9Vy1mTXXjSNNkT6HVMNGN2IfQUec+lYcRhwLd+YN1K8ILsWIjZM4MZ7fzxZy/CzQROOv2hRf8n
3SmYzoWeIl+cK0BrebYxRODdU7I4Fw6aD6vCyjL7u0y8lSx6lqSRWjqMxuPJ1d1+Vhrw1Qe7OvQQ
txzZSp5zxvYpvQynDqcZ6ozYlS6Na6zzQffdmVPCVnjJKf2b2RuQJFWqEy/zsggW0zIXN8YanApv
9DAuP3vYFGk4vUVdbL1XNa7kDMP9yeNRuIQWlp9yF5uoD6MncxUMi1dsW37fyLhoKsqHqetcledu
XunGbsW1P/ULfPOwbuVXc8+GrDyCrbEVRZJR/EnvS3TJLhqQlcI8ftIUE/WJpPiW5rkveQldrTgb
AWKJ6h/n6gqN3n6gHYqsH3b/sqIrVWQe8/epTgEiPhKJfTpjPIqMSjJnuHSFk7fjx3IP29Sw8QXC
ZjVUHYhEKEs+/LI8e0lSvtVPl9CQOrT9r6roiADW44Sk3RhQcDZbwTEwOibWktSnzmI1QTiFpoWV
FcczPLfm0rNrfpKQ7JvWvDuFKN3DmB/wKxZ5kXEgByHNJ/ugrVQ1WIlW9sdNdCThRoO7C7dQRSOp
Zrn5owIqDRyNRqgxaoMEMsMuPOVIO4f++ReOHOgJyQgRr+ZTAW6NwBsc81+jIMQuNe6PbYEa6Ug7
fbSctdDfxr26ZMexSs6yXdDELoAnKnNA/Ab/AYEgX16X4eEqflPE4m5zCTCLQlrBJi60DNPW6umf
8OTFGpqFwzyAZMSgX25fcKGT37PD7oq+7wA0E1CRk/ExQCJS43gRRLgCszRSFHpch/MQRW+Zkwfu
yWlxw+SSVAqvYQcVnHHe+yViDc+0kP+EcGEH6APRbjFOXPLBRIG5SNv4CEDptg7RuJ8FkR+OSqV3
8URNZB/onZBSiOwzj6yw9mC/O2Gr7JCoEU2Ek0QAtbJqlKBrZ7gXQIWOIxRZiSxijFKSdsTmq8RO
RL/PAPitbLHWRF89zbzbTVU5Lo9vPxEsfuaSh7GyjJiztVtQsTiMfyzq+41WdtAhVELUMDxoNwX/
Bl941CrBV3SOO7gD0FY2ooXprf2ikMsDt/fClvl1e1jvnfDHGz/8UMGcOHcVUvywNxUcJ7p4uiIt
EEp+ViRG2iGv6v2Tcau1RhQiNTA5Ca4vfC8C8WTI5JsIJfcozzn+FbL+F9/RXhCYa4ADQPfuttxG
I9pDY0pHONGLjFMk6bph6U9Q9IxrwOZFMMofCkhd5u0jZMcWKMcNhl0wHHZ8UVa+3A1rT0RGA5J/
kTAYiQa5NCF0na14xP0ZY36fcfMGaPvJwmXawBhCvNiaIbe3thLxIdHS/91bZJadIaQqYiOc4Xd0
3KWAMIKPTg8tiXNXY8uW7Usdrl8HVrKUH4+eop/MPY3PPz1JRrRNr+7BFGZi+uyqaFLCJjOCD0sx
t3RdnQa8jIn6IB55IcdLVkkjfxm0Jmbd5E8k+aj2KXo6T86sA3f1EEzIJ6D5whmNlpsED1YcPta0
ZYCdhe+oo8tAaKvEWyZ7T3llXVZCoWx90TrZ9slX7dJdJcyvBuCWJetzYmof6TiITkp86P0nxXeG
Iag52Oohyot4OjSY6KUjlqhXAAObOKkkdrZWKvrBTV/qrCOyzg12anh18Vz8pTAg8rUnwTnxKNGV
kLWkm+3Wifp7qFPVhksrXDk1VTTIHj7YfKhxPA5B7Knmc6Ic5PQ4hqm4L5PxSe06WVufkFxzjtJw
uTiecm7K6ZVJk+xrYm9rwZNSLAFGUdG+gC4HM+XxyqjjL+RTl8fHYSEy07RdRDsvXS0Cry/CB17C
3N2ZJlUVhM+Y+4aRJk9i/90i6t7x6SXQ+l/puHSon6a3GHYVggawH+/rPP6D996H2GEDPmsOA2Wb
lpgKbGNr/phvzfMRLi89ZsbtLCjsqGJx/hjNBbsFags47b5J1wGk+3m+Zu0cyyXX5BMM1ssxRjE1
wnUeC1aiG7eOAS73J7pfP+4Wi/v09pXeoqwKhjaCcVab8Em3cuaLpV3tXfpZiw9AA3KZRgHf4dp1
ftIUamu5q3Opkz8v3wUiZ97AnLUEqlhzJYGC9NEfoo4QDfWmM6CcCUVE/neFH4zA13ikqiu9EdKg
1ORFD2H0/SgKLB9Mn9IwZaT20BPrtkD1umREj7RDE6W3Eq0Kt+U01GFyocN5158EBG48Hmu9jtDJ
j3BSKCLnJ5rWoe1hcble38iZNT+ivG129dpdL1ryFe62YzYVaA4yfmswseYt+FAjav9i8MMoEhg+
34BsSvxyHMbv2w1skZ/FJw0xo/bmomsQxxm0Y5ERZCsgbZCTA7DK2erDJGvuWumpErb6Dqi4w3jE
hXbznECZKN/M8lHyiV7uUYyosB+5lmIZ24V5RieIdMiu0K9mFNWdjraH1vrO7qr79uFSc9LjJAJy
OMjqdCoqa6bVozZs2ymcdekrBcmAFd0MKAbRMEUuIiCBSTljRQCXMG7Ro1rjkIoWFgssLG/NwcRt
UWrp47CsfPQ++fRxXMjseJNXpb3VyrPBd59epQU7wE6dS+ymm6/JX/tx0fjNGq1E09iGLPPfTcfj
vX2pZbwHmm6Tx3oTGcXW7vUlgmgconC0JWK++6900ZwF/HNDyw0HGJmoZuScgkiWPFozvUWnhdtb
vJHqZMS8wVaof+F1wZwkhTgIiaHJgWlKF4NFfCD1OofZ6QTfAVM0cwWBapa/m5UMhtrbSxC7xinl
xQiNYvUX0gC60nhjoZ3iC/s6c1UO+4Aeex2SdQUE1ARZ6HNNGcCQeQgKTVCy3Q+44f63GCBXWmtv
Q1vnUDYiq4nqH8zFWfy7lF3+rRbgURzmCtusgsvKTZfT3LPRckAx2G/pFAccTLF3eOvPPvKEMdcC
/Zr5wHFTDfMSqUdVzgHqR8s35b3KrynEzf1x1jQJRGkZAI0/gSLjaZoRAtAdV7LlWJctigjIIf78
ZmXcBLX2qNrcjBT7VWmm5ngzZJeYKnk4IQAL2Dy7SjPCK/WIjDAekAic/IndkwhLRC43MsaJ6VJJ
3d5lOlqiFrONOWovf8Uj5omKuDSAf8UORS5MAB8JCcx0ei7mW2pLh1ABzBrVmb7ALKgIvGuuVz0k
Jh81V4LmLxiaf0kN/Yb4uUFfd2rhPAyHN5YK0DvbZBd2x34u8HmufMhxWExvbZxSJ4xC3Tofjhnm
Wqs6NDwMF9loNZxmFBhNdmeaVmX7RAk1P8RqraDz4u4hEdfag+OwiaY0915NJypI5NHpqBDEM7tV
54crfJJ63/zQHCOhOYkgFVrNiTYoJWPkCF0VHmyf0EgkKb1NhZ8jmr/fRrd8UE15oy+2bd1cZtpq
yyOt0fnMEgC0c6LgpUOhfm1dbUDBY/gXCQ7LvW9uSLLWP6LIpDBh8kU8p0pTev+SEGbARbQMN0sH
2UyCK27gkFT+ykP9/T42y1iz7BAEYUDcvLUNxJGhzXzjasj+WWpAbtPDP5NT5nUgJrkLiswR4A31
qja3SQ0zscRH22zqfWfdfNmOw4P9T90n4VpRsOxCTJ/tS3TTVM7Ac/l2NHhjwXG59ryo08wjyHVE
HVfO//CRTa7dUaK/hS8O5xh/YI6ODzCPNYRGqz3do+ZDkjnOE6eQ50OcjhYnrgar6kHRjhRJYTDe
UNo8ffI/ewN3RP/E3ENSuoGo3YVm2Z0HY97/M0UpVNzCPaMUxJKhZBhJmVu4EiJ0bkwSsa8hXkJU
PwTMJcjIfD4m9xSUZtpsUsHDCPoVHFYx3AAV7+Vzg2tRbRsx1d3+O8D64bmcnMKpPKLwRPnDXE5K
0fVFqwuDFz9EdkWJrh6g7VaxTXzNGQvFla6RiwbxZtWe5c0dNKcenhTm0IfNKpzHH1/g+BbZEZA3
aQDnXpafLY1LR+3b0Tim6RyZIxorMi2+d2CtuMuWURo5mrj5ubWgwXLiXEy305qnl9mMJyniBu3B
PBHiGY2JMJdLMXjNqT8Fwbn/uinmJmgXnnAD/awMTbEaFuoAGtlFEmMiHG+ltU1Ozbyew05ESrFN
XD167uhlsXGLgeB36MlH+mcBQryjLmotMwHaW+gDV8wqEUEVUqOw8GqOCzrGimfC/BzXMqWnfrdX
74pJfMD8TABr+YHXrTevLjYUzZsJ1KIKDgUPJ5CtqPkavxUEx1h+R/3cvuSsipJ0/CzJqAZ/Lvtc
q+EyhWWCWVZskpLat7qHhNOksscka82rRgitCCiGG8WZvS8ehRyzRtt0zVLYu4pTqYLX8MRAscFg
l3kjm8Ziy8XDYLXMdQVnr5BePdn0Jo3ILRAwyKTeFzeLQvxa18xuMTkAROjVycoQkijZneBd3Eky
NntCNRVWY+YdFDsi6l+5cj7rvANWisBjYm0bublJKZfaA3V/Glu3KeqVPJX86g2c+aJbVbl77Mc/
ztC4WFz9dcjCHGGCGtaqzdtjkEhRiTQp6MlG1qAaQR8r0YaAA5b073vQUxhDZ7I787cV19vP2hgK
NZ3s4TByIGztw7Ks0e1Zd5/MmucfCfanA28gKpc7pFFNJELhKTdmQOzCNzuzwNQSARB7g4axKiRh
KaLN8FrQBs/glsCFwWTmB8HXGLesCsO+dG1hJU0Zr1O+9xuu8jlNx0f0Kf+ACbv9ODC+5e8NAl8W
NVyY1n8y4PceQjcaLClm/YHdnEf3MqKcWFkYakxZiWqg01jMzvFw6V9tYDwuSxCwM9Nmb+AM0mkm
GwMIpImdfI6+YjEeon1oAFPmtRRWB/25z3soElnLdH5I1DSa6zn7ePaqwYt4kBqjDNv2W9i+Li9E
22KlqoGD6WLPqZPrx/iP/XdxxZkrTai7eU3kWq/jW9VGSaN1sYJIoFGZnUXUC5wMgv2D0r82F7Hx
CFONK09+fokwjdY2gb87UKgPvYoVYtREafs4vLy2l0lyhYaP/fzJYNjXEo3Xqf+BogHHKIf20BUC
qR1GexqcMv7AGB0uMNw3hlRV/38Hc77G43+TcJr9hzAtHcejEEiPtvHXB8ZbOsgOEuSeuyXkihn6
NsfMSDX8M1Lb7Pj5fB1ovPX4URwYDLS33YQ61anSMcmhLJb5AGt1/UpDetKGRz63NSjx8Hu4Ni3n
n+RsJFyYFzT4QJh5/vFjqF0ZzFOpLiO4dghthAkPOQUpO9IVZo3xNLR5dQ2+7lqD84v/tapjyvQK
+Bkmv20zzV5tIDouEFFJTMqjANBuYdi68JtYyWughleJ7XsDtsg7Z+N/pqku3e5ASkVICMxgCAkX
CcSpgX3SiZVkO81oJZ4T2I9BPj6B62pobJqzAxK3+ozBcrfpDAUvKM5GCdcR9eaRnFPkCRUqrHg+
demuGNdqOsOp/arsCjB0nASPdhzxJVlbqxKHOE44EWQm1XJxfpBEQ5hvF7CCK+t4NFZWHx+dwrMx
wKQHC3SFnrySocE+GPzwwhrzzF0JwZfmONbXBwxG5aRUlagfEuBDF+4S95DwlwtlmSJhi77ebhlG
Yc6N7qFNLKLP8yM672uoxV6XdnF/kLIDkYYpE2Q02D/PWz8hXSrRBUT3MTez3OmeAtuURJQtogGd
X1zqDGrOPir9aNKF+cQPXKhpIExL10BmcH+JqjEmtp4eS6gXu1Gui5IFf8nLfsbmVzyfdEwHigTK
KfnqAFBrT1+PMtfTExcjl2Q2yiSEVijJKYNxGFAbeWAqR2zW10eBvc93fVOgtLmco4+XVfxiKOWF
wnKjHuxuwUbX24HNN4d2cVWb1ly809vrKzx5WqpgoMQVvMF3Hzw4alWkk7fbpiSo5QWK7AYil6ck
Lw7BHLAXzH2StYWpb9dy8AG5JsKxH7CEXqMCX7S5d2SqLrfHzPwNEahb6CB9aHM3Mu3PCTX2UvB9
gg9NI1Y6bFwm5E+fS5fx9R2y22iSL7Cz3qVgy7S1R0E4YWAHGjaggEsD+Qt9PN7s/z2eqIXDnJ9/
pBzmZHjNLS55Mqiitmt2rARWj+OCfIpw6JkjB9jm9NHuZj9o0I9VO4krDs5SJKecqXm1OfXwUb01
eGjvVEI8D5MOD46dTFvxW7yZjy9qe5M9ef+bDAdY1PhsI/70UlVMaD/i8uaAnIliefHkQrJpUBsY
bmprkCR0CFHwqLGuQnjgPhM/Kt81/goQezWqNWeJE3K+f+jqu7MI6TMLYVIFf5G/jwpq1DIejV+C
B/4s8A2K/AvRKz0sce77zZB3YpdAfJWHjK16J5qR2KgImejZ5WVYmMrrM8dCYADnqpn1zAfjrMQx
9/aCobCnP2fzZQB3/BmJfTIoRb5cwHEIfRZuqbP7EmYQ50fpkj/vkc6icaJX4GQiARAwJIKWNuVJ
odqQiJFOFh2iR1JlLdH+WlP2pY4sagN0tk/jOzhAsBU+Ppe41hY3fz5CRBrNVv0i69O2gl+vAZzI
TYi1krG/KZozR1xPmMQ+1D9aYc7R1O07wgxH5/as21+7oI2naJuWIfviu/uoCOKGAuv9u4pjkeq+
BlgLDhJWPGCwoUiLHnPaQ8LvEFfmMOQw7HTzvbSyqWhOmOYXUJRjGo62MHhw1ThFUTxkR0ERyV4e
oUzqW2EXGC6wfta4aV/KLJAtkvk7USLhyRD9Bd1FyO4G4t4GO4llSz1BaYhEiupi77haJy0AJOcb
xOKS78MofgUlYduVXsHOxERhz8GYIOWVe8kQRY5l0w6zugCjV9IOAQqDKhTdlAxJOD5663rRUVqY
jKe3gHFvQIPVe7093Ihtc93wcPN7/o2flRMJT+rfkOapaxBsTrpKqBLZjRXnYRpIM2HYAoLngkJX
DptO+zleQUPW+X3H/kvYw9gp3xJCWPStDDgH+uV+vv9c7rPa9i6RPynysOSSqc7AszFQrCJOIUpr
owTG6uzlIWSfZUIxQWsJJJsotX/zTeOiWKoQb8aSIGq40ed6cgmLDpYnq/sjW7YprakDBQDWPo/G
+rJJMAL+hp1WEJ3Zma+WNL7T/Ww1FLSDgMuXrRGfwJTxYvDJMiQ2qWZzHMXhwIptoPgw3EKF6M4V
VbXDwmfazuXBkg0yMb1wAh3NROf/rU0CQxnbr52JWIV0UzHczjxy6fzGk80tfQwKKHe4vNGIqrYx
FSfFQSvPTOj46K8o7Ui/R1Us9McVHK+TbAL0N/qThkmNpyHl2/deZlXPojpUGjh6lTSat2UUg7sJ
riiK3z+NOjwkYmVnA22OFJ2mNyPkq7+qeXyraZx+QaOXPsoPhtQQrN0Q9sCswdtuL3oeX46S1Vsq
7P1fL9PKWIRFkG3i14rhb2C/VbSfRlUbaIrO9AktDwKeqYLBwr8lXrfm2RNhar8NS77fh8NlMnOg
Cs7Jq4pWABzl9KRL5rjZtG4E9jLLe1ZeJoSLQBbc1M8284zTjhJwBb2GPM9KzvAvq6hG52t82TZy
+sjzAKZm3dmZK/C2NZIbPNXdiZfjpUjq14FawAipSY6X+PAY43YOrFcghgLbkNcKgfiAhyb1jkpr
V+DcFXgnTxj+yInrckmiAfkr4WiRg0sXHUeFdscrI2L8KiyIB94hYs4JkluCYyAZD3Ij7E+IhKbG
1QwULfxtJwGF3qi9jfUaoIktigSZfFIF+y1AkAv0DGTt2zVA8eCdVwvWAFlHDYl8SC48NU4dBDtQ
aKgM+pWtwDvQePObXsYs853g4RwqyvCugTh7Oiix/B0jLtJkPiPGc9fvbu6ClgI21s09kD4aX9AH
FPqSV1RgqxEnYXsZJzjgI3RYAojwDqJm/ni3YgeHfSGOBbCaENIY7Zx8DFr6r/qzLP7RuFjvVwGc
+XqfMSiduRjArQlpZaPxbp+eklqH4A0djoJGMoM3PEWqQMKsjP4F+mtH5hLoJFbE4ZD0O1dMrZwo
6dx8ZcnVx2LPc2dX7K4jkp4gccuMMIqRmJaF4iimO2NOtpXkAIF9j+ouHZIPHcYGO7Xv/uDRrmj/
Jlfv9shosVLIh527dgeW1rFzf/2wbro2DF+W1pzmBlnTnKUvGviY+JEraFxigjqn028kkRdHQWhM
Mht4OZCiEHYmrlevV9arT7LNKUs3Toh/xpy/PWcfwnH1s2HbzaJMegBivD9OtObBm9B4M2UqkVYn
EI3jSSYYBRUEisCGMrLaeFhMiDA1HkTGnTHh7n5I8l7hiFfPwY7/FYDKFoIeXegaNydp2fEaBmwg
5lBVvFm3j4I0+5vWLMytjp8gDRZqy/TxyOWRThUWz59Lf1ftQDT2JYr04MuNIClfgnIjSxKf7NeF
thSpEbrf0Uk1X0/bwRs6lwNwR0LtVuA1ghp1//dUrTf2iHrp2hQB3ID46MhzL5+QJw/59UtNNz8w
eSAfRhpYCbWzyiJya/75m6AY5OwE+UtizCnA3v89KT+cv7e1Ew54UbKUcHDGAXbuhhBQqjCCdc5A
N2id+zEhWo7WKsxtfT2bVdxnOALZib2BMvuwavnDY9QDPx7gQG9KPH99VUyYqupXEUaKEVVLh7iS
1Gic74jKLiNQHxDSBnBGIpLhKbuEnYVw6f/JbqIeawnxRp1o6pnwsjTJLwXHSv0IoAemBlrFTz09
KymZGS4E65gT3gmyUXDgqbYErpqgQ7UEwTt8FRqxBhHQ/klUCdk+in0Bip8ntKgMqSHS7Npxqt8F
jhm0SBUnIO9VgMcWZd7dS9Co3pttEdd6YpNn/t36EP/4mhWisrpLxBju2TsMYN//tpuTx+opvYHo
AFkykz2/FGfE8DxjwcK6vShgjtMyiCXhwRUUNeXDUl4lxN1zw4Ttls6AdtteC3tovgR3A1ytWm9l
8Dl4Ch18XS/aQqBMgn5i2epbfCILrgC2bm/WCUVvlsWkBY2j8XoPl1O2Lp8L4GLewJ+otDzTSK6v
pPMJMYj/huMYiu4F6thDI2umif4uaxC6w7/uW3XX4ZewxstRV1aIHbV5+jJHyWMkTOSjmmS8/Ck8
7BMVwuSUXB0G9nd55sdv6JeAewqhpfuoy3EWqdr1hiFz84chtabnKRchQS1JCqa/GWVJDUo6h5ZO
lVJk1aRdu76+VIvrx/VCTUzi9azeF7FFAWPsWN2gE7tmFWt5+jVXMJ2NW26qi9CoWQh5HbPYZFVS
UQxTsXwt2Ts8sZqV+aipkWoYrNhId/DQABIAHT47mw4lbxvFM4lS73uFTu/RVOSqYMgBOWX2jn8W
2EiJ05BLPmjJUg+AVG2AHkMvnYRquU1uVsu3RUR7oyLJVodrBo5m0NzJ5VFjMlNb+08OvS5Sbe9L
wmP/QSTdmEQMOXku22gnz8JaIwlQ8ZEf4kjuaCAc/J9iSqq+LaHyLgmpMOvyrO7MBiW+hpoMf6Bk
gxGgX6gcCQ5uvhOmhmNImTutC4NMW4FFUREU2Zua/y4EPGelX8hPAFc+uQ+ggP+Binwla+JbCoZB
iZwNnJkJZCewTYFBS5RSN6age56ODMGKZJlBBhKH+QLAPZUZ4DlzzZu7RcusOuB+73ezYDZR9lQ5
hvdbW5c/OnpDQacrCBwTtoy3x6LUwr85tdULsAvyhCWiCLMVgd5wgQ4z9cLCDf82AVn6wWnf+2TU
jBLrhsU3IQW6rbLEjtWSdieoj7+kTid6sk/XU3+7L9aMZw6NZQB/jrLFGJSi3CsRBR8SW//in7jo
IQYFIWTRajgn7tqqJSoSdtY7onibqLTdyB/gh74f+QoSOM3MIKUCIzradrUwcAf8eH386DXf4l29
2xX8J/Hkga/DB0jV2xnYO1lRUjDGgfIVxzThuajyYBxnUxhVF1kLvMl0XVsWOfc0LI3W0EUeoECv
hqg1jWe/kxkdAOFjNe/DK6otIZ4xmKCqnJ7bQ0IgGVqukEezL+4MrGlR9l8cJLWXIW6b/3xfQMoz
v/7lbveJvo6DGa3P0dTZQRl9HgXM2gIPxoK0DUknbj0EvKi6bi2DFt0R6PEObZz9zGzqoTbbFGpG
IQnmN3SqTHVYzqfiHPk0Wh1lVDmg1+A6PUnIvBAqStQYxA0swfRwDPFsHzV2W/IVU4xJyDABG1Zh
H252F+dVHA/NQmAbAGt3UrsdtqayiywHQT2XVONezQT0S9aR/xW2enHD2eo90GGgpBgcG1H5gwSK
ESaaHgGz58HrHv7t+XorpVFOlWKMsLNFqVp3f4xTCtEYMIcKXNr4+xMVq6J8LFJ4/PDifm/28KsK
X422gbSHabMBtPBGMOvQfKtUuRnpbjm0HlEQ7D+E3M1MC/fv+oK4Pz6Bi4b0g7YTsNc5vMt4lc6f
4At/yOvLl/LsF5U5Ets4fb7RsSEbs2VfKI+WI25D9QKFePI3au/b6p71Q2xix+aT8B9W4hpZYRBI
zsl2stWAn7AQSMKf0j8V62nTn0ZqGat5m01c9iy+rEM9wiW69yCoyNpy6wwvL74xwiQca14gkUJh
OrQNZWLilKMG0hNG+CMcBP01GFjLbibjmHu2JimtwUkaJAOCe/OF/qaM6Ma1pSdByRY+A5Vay/y/
Hy5CIrlRWX3NWnijIOmExiww78E0VexL5OL1XB4qiuZgAGv+Fh9DwgvVHlr2fkeg5C2yL74vkmea
rQ1ZCMuhcg/zLBkpYwIH0en5SeDybuuNgXnCwp3UuSfQ+svLzuVBljsQx7vodiC55AoJBmAVmOL+
1GAFNDMVz4aanljHndmFzFx8FPn4JsO2K6Vq2b7nxeMAyNgt1vdb2yhzztO4nQ48T5idVcI7pm/e
rLwe2+ejx04EzH5W3AQL/2ZoDidtz24+tiFMCo+Cy/4F9zUuGrzQNSapiLUg58Eovk7ftADHDHPB
/Fa4h5YvjhCRnGzej9NK7dNXmOiyY1aV2H/2oTe70xarBHzL8PsT3JEpWS+A3mc01/GShZHhcTGg
O0geFWlsXbnP/BCxzWYKX8p26h/9PwMiJfL1CinpZW7kJNswbaA1D3wDxEdEQplaw+yDOHHyDnuH
kzgXOVTVc4t9qdYr7HXXCGo6XlHkl1Ry8FygWwOJtVt21nhIhkPnm0DoUGd/ry7Z5oVX2aFRmp5r
jpyAXgrstCf2r912S+CUxvwcArUlZX4TPXDgMylgeExRXZmiIuvxWnoNP+Z79vTGZeEDQ+oHjP4g
vAoUOHpoGETXXc3qFpRo8VBqkul8X6cxJ6+A+d6dNzKO5jk8+0qp1HfUst9DYJNhVgTX043YKExc
3jFoQUjwjjqoeaATmwRtm51hR8CA/OSgjn3PTrmruXeo/wHoZNwX5gJwsACQJmT+soHfiDN8pQHx
DVuJn2UgmdMJlT9jKNbmPazUB/YzOZXNNS7wOKjg3sodyv4yeLdXAMvJPR4jR1MUG9bXNAzpEuUA
VqexochFsQYe1lP93gr3gDbOoAJ3bUWL5f3T3Q6ZKmMKax/86P8AT8ZOzhXFYShd2rmPny1EcrM4
fu90IZoV31gosouK6JtGOrQ5DakYTv/LQgfGfJnPKPokuJ3WFDWGiiHvzGp2JCvEXuHZMZaKVHMF
ea9bEg+oOuikOqieXQehmi2etJKWzfFTurzIEJzgY2YDvCsVjohJXFc7swEn4Tq7QFUGQW7wRYtb
B9On7KkSkEJtPc4/ksoE8+pxSR2J61gUIzsXDg9fI/9eAjjTkc2uD+9eMqdlsVG2N1/YMKDR11NX
yMci82CJGUnfCuUypDnXHeQe5UK0SACbrBBDJ2E4X7iZSrjjZMBuKVFL8aCtxWzryrifWhZSxt4q
fcr6CrDxYHe6iGFMhYlmHJt7IUJ37dXUx/RQTc/VUdI+8eppmXNy4nuPg3Jk4Z2tSiJnduaN7OLf
AKixoaok1GHIHURi9bfOzkXRAXbtOoo4wqPsRvUjZg2aIpHekz2eeTPtSA66miiCgxpr+AzCMXjW
NS/aZa1e1+Xm+SeMJfg0k5srKDvWG5UTOpz0FYWEs2gDjFiOVcKnPxj7MMEdbahVr9F+eKk6+LVo
gou7NizCBBHgQPzysbj4+Hp6XBzMxQX3AIr4XVty7rLogoZkjbw+FErctj3EcLQ2cMjzsK2E3B+g
rbe0PZgdPfvrqRBc2ZtIz2UyE5fLy7HuP6ydDbOHFAjY0CvgweHUFB1n89mgaal0eC3ENuADrpOb
Jucy5sQDYJXUH6wj2tErJbgMP7xHbKT0zfO2vrIIrOZDTQl9uYGFRUEzX5WeBNp2ej+ZwDGKBcG6
cWgtAnLugZMk7kD79U2o0uh9yBlsQhM9M6keU9E+nvPpLeqoyl6iEA8Q10ZF0QsRM7U97QokCqe1
KGCaT8etocAm6u+UWIqcjdQHhu/nd+afYVjV7Z2VK0utDK+yRq9J/A3WGaeKSDdudclkzj+hh311
4DVYCvrQecKJa3+89LY69QfJO4qzaFpCby4doKsCBTTSIQp8J2sgIPZe86DY3Bls7uXPV45tKUxZ
OqvLmibVUKNr1TzPhr70ogwCiXAT2csTKdhOjpNLvmWYwklgKx5ZfE9xI/mzR6BWVRjWvA9y4kzu
lzyiXc0oCSrTSaZcutqgIF5gpHnVc78LWQiEPJ+n2UNxTscxt1uXU1xvMdrHN+Y6I8Xf6ZICkRAI
2B3EyljxPj6eSDjzeGTxTXLoBIkpNgmP0hbEHr2NVG6VU7TTcahglDl2TAuXXUsWlJFrJiHPppWV
Hj5BJR88kkpp0Do3+zas0DVDHWM+Es/o70FYWKlLQ/mLkv5r01opoqDfnJ83QkFkHExL4QfZ/neY
thTUehXBe0IUPMvcn3c+sHdbaUo5mWJkGYymPX6I8PRaU/m/7Q/Wb4CPdEmprXXN0tJeLtczz+Yu
SP6DLJWULRTAfpuZ88k/c0khjkFR/70/x7+FsNjja6WAVrqYCUFTPqMBu3pMSd7IFRjMCSfhqhe/
47R/rda9EjR+vkqk34/fPi9ZC8Zc0l/i4GZynfefvjp2SoKRRzo080pgFy8bCIFGdfsHeSdmGIg/
abOCDIsKnTwfnicG3Mx9au967fBspMM+lU7crRrTV7jwpNv7ZIVB+1nTTXgnJeyAg4Mmdf4DCZ+V
Btlsa613qNBVny9OLFE27yiX8txye6F7S32OJFQevto6bwWzpWkqO9amKBnF/c4qxUmNRP+H1k5h
OkUI1lbxSuz4aS+FPpbzKms0S6T7ZkmM7gyNNMxu/zguuNpH3oUewJhqYWjR7RiUiJ3YFBHjCal0
fK6WOSsizSawEyU5ObgT4NxrpQmEc8fgR4t1cRMnh5nlKQPMKn8hENl8Pka/sGoRlBXcM57034Rf
XyaOhah4xqyRz7qF1ek90y5GMOgUjRVAwGJeDa93BDr5eRD3NLc5E4lPhH0LkuAzrGKG3M+EqZFE
z3AHnrKc9uSuy71/kMxEcMEm+XJh3RQa+Oy1clFYXUHd/VX2Kof7CLvsx0p4QlETotb8+/XKSIQH
gerBTDjNvh28UOcRFp/h1AT5L1qh6q6uwNvqZCwcNbMAV9vaZUUS7XYnONxOqAPFm/wUyMxReIEZ
5gzd13GKjqwcqjZFBu9MsYjIPgL98bvnmBOok+voAEfoOP3vG4lurScPJQI1S9Mvz0CPMtiFGFO9
6Gnfd0xfo87I63G8rgPquDHOY6gOhorxRCjDBxWlfpz/ZbRKABsFWwLlfEG7aj9ryPYS9K4ThWr5
ZM46XekVdaYHGhyIQBJh+hDslOrwimILon2EEglK6Auuiu/FOsg1VH+rkFUEMCjxj94Tr7KJgsOl
KhYsAqXeRv5OsjmMWLejx1r03CokA4T3/QGxMR4JNA1DR7lmHrT4U+x0Dwp3Vg7+4X+Zm6b9xlow
ROCbLf30dB2GUdH1jymY1Xw2i4KC26lH4CltkGV/e8QTWryaQFYrenNhKOokMgW36lhAdVVPAhiF
jUZJhUpUkAshNJwfKjfxGVBw7hwJFCA9YAD5GxEXNS3dxO/BDGO3UZJcmWo17YBaKK5IZtfbxlKr
x0DjzAURZOWmGnlBSnROrsy3oCUdorpZt8kzHhOloMAouIeZ+T1UD3YiLdK5NCSpI/kN35dD0I4T
BwpX0cGBIxWqZ2NwR/4TLvTMhN5FXfaHusPFt10Cn/a/OE5CGOOuGjyYzlzRCJAc7yGjc+RnLSGA
IZkqLU8PAx9NobQPvv0VmEFli2QNTkUe0fggntxqi9PjOTHJwBARAJZf/utjbAqnFTCCtKtfIDOX
jBRMIVOoiSxdtY4FL3GXLmhU+RaRKYfQkGVdCg0SOy2uE45pIslMAspv9tKQvJMwt9cTzQ2MUVCp
8gW5meyxE/DJhpzOxseg2EiIgGvIx/2Suadg/JUgqaEOcj117oBkzFgcKtMgy1DjzZcginc2EK0z
3XhXyMf9UI9BAtbGKVqcP62ORgDGo0LGYBNd6wJTXw6aPJS25xM4mPnXYvxXPQ/m7XtEdB/+qaKt
AiIO/kidgfPTJC2XKZ/bc4xU08zU/ljuzfr8Vw5M8hkEzN5j7jlv4ddB3ziMhqCX0mAkn8IGB0q5
c1q/tzlAdR9y1As7S6q/eZYLHVtNErpzgsRkGd8EGRpNmO3eIflkRoJmZwJsKn3tNpWnKd7k75Z6
oX8Ul50yPaC5o5xohc9+1VqhPqLlog3g/7K22Le5nhKx1Em332BWE1J0Txf8qgDoB00OsG1VVcyl
5nZFe5wITQueOA6ZpAQ5lvnVjclCUvDpQj7kVz7z6sGMRFnfSlGP8tIoELoHFP4QRCiFyaIzZpXD
zsBHRDeu5sld1G8MaJ5CLpj6P1TyXelJU1wxYnBEt0Bct+493QYYJv83gXznP9OO5OfwEHXhS5db
oAI9ZJ8IU1tbErBg+Un1nab4VThnQSkoZBOjJsY2ZZO6703Pnx5abBzMtj+31a3Jc49a7/ZMtnbB
rfCmmnQPtT/FMnHzgWUNAvXQlwVaK/uPtVVJ2DVDA3GKHBF0xa2x0tqgebDik38YRzVsAcM3q0lz
HqF0wMY7bKGq3/Gv8G1GgdORKkFxsYDgGAnYJl36JgdztyWlnAm1xxmu4ku9qOn/IjkAeJ9tGOJ6
Apdz8JkaZ8zvQVf8kgOZ+B61PrP4zDHwhLQGr8PfrGbDHZI2geKPmq8bVyOpEuYrUDULVf7qOUa0
uJ8jnB3NUXP2Xy6V3eTQEl1gFibsYAq9k8QkiRnaBXeHPtl7E+fdFybtqWKk/D9xpznYIYwCsN02
SHZJLRAX9Y9MLLYUmOmZkKmedDEYMfshgl25nN/H/qmp8p/apDPH66cAQxITk1p0npHVwbDLOwYE
X/hR407hDd/IJAM+WC1dtwYt+4W+34I45PgR+WsF6qfsk/PtqrUSpdWh5yLyWrjwUktISSAND/Ll
biqRxuaj/HtBQ2UrY8rkrGBwJ5i0GfTqvLjEB1F13aBhRiamVTB65TSy7oMwWA2+3SsGKVLm+nUA
ao7jjPIUTIJ3hHyHkJqevi7Pzyjf818OUPNDl0GgOgBw7cN8yhEy486oBE5nt2NqF+jMUBBi3WuG
kUr6wmWgb4BuH7RG/TiUU844gNN/QwUs8DQtatHII02qmjIP2ccr0BNkyUW6ohxkgJSW5ByeaU+z
yPuLYoIwcYmm12UJpLlV3xSbkpW2gXWs7tGDS6u2nclt2lsciBKgc0s/w/rxH2UdqlDyaI5F/2pQ
pv4H1y5tK2NaLGU1yWaMoq1ll7NlQzEKxVD2hFD+9G/dpBafg0NBKUJNHxkD70kLTvxy0p3Qk2X9
mtcNaXS0Shssv8anytsx+tsZ1xwcV+JZoct/5iEFtJoBX9FJaEeLNY6p+rH9sDETZhWbAqU3bGQs
TPcVgy30g17KAAQDARqiJXOpPofI9Yb5T5Acwv5kwWbNRXk38PO0ShlGC3YCWnxM5OmhHRDvcqZz
FeX1uDg9zVU5UmS4aXkXvZUzqve0LAIxeZo+wsyKHFIKeC8RUiUwD/RvS+Grkk6ZBNNssfb477tf
aloarO1IwDXGjk65iAEiJYF8ke+dXMUrUlbOiA81amAUwMwp7FGxTgUQAcWQNuzKkapXpnJ884kB
16dut+hUSLTEvKWVXhMzkYB6TZjcsjrZnY21ttSHH7mRzqCmZxksdieEwIirIjS0DxNkkybJY10M
PWyJSqV24JH83aV/Hqwv+FfHmnQf6MFbfEGDkzRbE+66nsQ9HnQWjP908FZ2SvHmZzpsqAzG+cPv
NWCmgGSTN4//628OuQ/e6VZJ0ZtjArJB43669m6ed2ex4GNVx1Hc9YdmNEzv6e6kwVoTseqTz+Ol
6tD4pI1GIHDmKDCtMdm1VBzJmSAG+UK5OWyF7iTyupTfGUs+zaNQQrhrsZIaTPx6yI5rtpdBo8hO
eyfxqT7XzT+aYjAvH2VFHU5RJMjlbV19FE0upo9rik9dhlUKWrvjXl8WaOvE3LxvJMHxyjxwfj7+
SV+ReEllqT7S/XmVjgsgSKnTl8jA4pEHcbSCHSX968BLWXv0iCdtqXSVneKfDjuTYVO4cpYqBSa2
CJFmLTVV+X9A63I1aqThDGgDh2ALsIkXNCEj77iXAmnfp24jgvZD9OAuC8H9VsUnFd5TpEd5in4n
3f3W3pg2oL6w1rdeOT8RGWcQ45QpmK4to4jweakNqLsrk2D8KSkPDvrIeF0iBsiGk1mUrEQvgVbD
NIzkZ1W8soACijAoanF+hijReaqhS1ZfTCbJ9Yb+t0Op764BsTF4cOrxK93eJ9tzDkRmtq+g46nN
Y5BRM7lCibFQrv3fncWpvqXyXWCI7FUUaKAjC8poEYhZ9Q88/pOIdw6LFfFvbyBmQiDuhTJms0+f
69fju4UfKaBq6uaS59dW+nkVE4eSiUi6DTW/SmLPXW5NRqNQ4rXHFL4JGz8AihaGfa8J+JvqnPTw
ixqOljVgyt6Vx00R8+gyr1kl1bJxv0r3ZUJLbEOnbkXFEjyz1AtmEuUzWpUL6k5qqF3xpMroy72q
FCFH9iRuxotpMFMiOHQFhaLiYH5mg7GZgtXqxkctC5Cyv5okPqWcFxOALQWXTOvgTfrZmScJOIw5
iSwpHm4isd1ss0qLPvJ9AXnrc8xBF29f69D923OTWH27x357LP3erC6Lx8PYkjSrFyZJl5jhQW4j
cxYwTyFd+ZLUqkGEqQiat07JzD/JwMNK1EtA0j4yktUfu4bV5IgTxasgI8u+vE6JtNhxB7WzpB+D
3iHZcqsJAb6aMHRmMDMHUBISGVDsQo4zP8TO8LwdZnxSa2Ija8UPc5TZibpO0S7axyPC1a86yhMX
oXUqGvByvWzeRAhkDgcunwe/yUMCdE4bTOJAYcaPFm9+rka4QmPio8uIxOxdKyw6QV8rArc7grjp
3O0VrvXOSM7SnmPAaqkZX7Rj39digcptcNMK+8FkQOVU+nnSEhiOJGz0TVQDyoC17aPYoyH9FylJ
lEMgfuHaC+WxJqhBHnR++dDzN+ARqHLAhG04587eJbFnDLBLvlhRPV7EfYNfuCn4sfodjlf0lXe0
dpHwMaymkHQ82ep03+pKGTjY4+TYd6SQ6RWPl8wKv6XJrIGH1p5k4P0QZXJr1ZSO3rFXSAVtgfVe
MGeXz2YSJJqCZM3suYPc95tkmRxpn1/nQYKxGg1fzYabGxEp1V/F55i0ExPstqKhRb6qMk6HJ5tP
zv4k2hLPaIeahCbjujhYHlLDxEslbQLbN1HaGE8e4Oz7W4hoGQxQ27jyuQkThRpPTHQSBjwiMZdd
7tBObql2fH5pndCPZWyqlM+uKiN4O7oODQzUuyDixsS1sqd6cuAjbk0Z4TlrgTNwTF3K6RbE6i/K
/c1WOIbfXc7wNiPKMXnBRHia/z7zrxZKjH9P1gY6G4qyKlCDN6o81ajg8CJ2mGKi/A8TJiPKiAxy
mFiZ3pv53xBZ09UvorfV7WAmWg+0SvZG+tvIsU1SletB//abvHfD4algkATK9c9iLYK1bn5AZOav
NRcT6gEOWNx+koV1oVeyZZdWmpzxby4ncJuwuc9OQn6RF8DZH7c4qyB8lnV9Oi9V3LPkcWdc8VxI
r3ReRP1mgqY5ILDGGDHEqV2zxaY6IAUyPfLSf83zctUGn6i6qokomdSfGPeo4rxopggtbLkzBeZm
5uUvA80D2mLFSnb0mk8MforLoAqrdfhXob5sGH9gEMVBf+3S/TvBoOBkn4s1yxCu2FNa+DBSkdE+
UDRRy97ej0ftSoSTcL2HmRIj606u9KI4/yAtNfY0PGoVwcoNmlOrgdJOXCotyd2aIPGiydHdQzlT
NQxgMJXpkWgRrpdmZKtbunt0XFX+U042mA9CAJlBzEPK5/XIzmQrnltzBfXzg1t7n0hZPdgiTmsA
mGdooVZ1kOwY/ugAGMjM9K2kiMqyMywLAc2c+4ZGCcgpP1Dp5gWsEs2rXf94imYE4Ul2vW8pqQuK
COtQWN/gL5+YbRxuuYYA3iYNgFIlBG8iLxQ6HGxxtX6IQoIVnwXzi3EWXQM3+n7F95QQjvg3Ie4W
294Hy/pi/YMjCn4lpcufzuwgm3CQR6v+tPTgPujAs/UgzNs/Tf9e6EKNmdsNUrOsXQvSqfpUJOyK
N8G9V6lHsENkgc0YJmGgQ1trF9uNhJ3uZTXvzROmj5r+xPhXxO8LNZxJimY8P5DNrGgE23CTuKm6
NUGas7dMVrEJGSDahpaLXJ0fnpEvviiv93ehe+j7bE6bwBJ4KE0IWVhNAGSGhe1rsV5bHytW8TrA
hjDaZjcTyk/a52Oe02XB8MLGemAYtJ9JDeUGmzqC1sma5dPnnAdvbfvDEaouNzWg+YSg6MQ9OJmq
Ae0jQLWT9HYWIdP0lahDn+sCYpUUIpqaKwbgQTZh0FlSW3pjjHlltL8VD1+qmnypkmJaZMbUItRM
pBH46FyEGlLAd1AiW9fl0FvnEnf2hkcK2b8aIRk8HMk5g7P1Wxeb5DwlJ8T/oqDEE0ZEn2jdSpmv
iupDz+ZmqYmPOQn4Pd+rJ7k+6e8s7/fu7qPM5rqq/ofcBf5pNEDjD9PEy4II7VvvFXWkNy8j9C6q
t1qpYZmDoSOurMaEY7hoB+TF/tBlD9Bf/rbxI86eqE96TKXSjoCRJQ0w/18DRwAMYSZOuIzdoLj/
v/K3aX8wTFyFi7tuzEFW/hWd8mBkWU1lDPeubjMgECiKDzQTR1ZC+p2NM0bFj8mOaEI+ZnwAHhjT
6mR6767i3a5FfdWFwqyriX19JUncg7rKceTfJj4ZJ5qq+Z7BvIeGpBmqsG4UeHwNw786t8n4G5vd
8+PX5LMef5DItAb/VzPvhFimdeeeQX/U/9d+cZS668VSN/xiBzt4osZudLGj9kxP4TbZvqnxDvu+
n8Bwr5/yIfrVsaQTzYT7fMG9d5AM1Ne/VrKG2m11k3tNeI6KlCSFDJT5yK/7rXqZieGcQ7JQ0jd7
zNMcFgtj2tHn/AH1wc0s57LZK9Zn8zJzRE1UZ1in0SDYdIv+Kr1Bdi7+Pr0RD+v2FeCWC/27MdsC
RvmURj4+ZH7CjS1MlcjeFOTcb9KJPjEA9cr4S0Tw8v8BwQvTUyQUo4r5dnFWnvy1+kyzfnbqUYYA
FYPy/gIz3iWiqvLzL+y0fX6CTJURXBJ6s+vK0gERODl3a4VTq+Y4LIkr20gvOXjPRJ3+W9WbSsoh
6emgLciO/giRAgLbItwoirlqnWbwYs0ftc0DeAB/vJlmT+fRWnKe2rmFckKFdZlzENO/Wfi/Xjac
rtcHay8IKBMBJgW56eTuHUafYVtLDJWVSOL9hTtkRlqR9kJ4OBlCl8UXSvIEj14PUW3NOQB8T4+A
rMXo+qJK1aXIzotPoCxD8dUWuMj/Xv3kzGwv6aDJHsjRj0VrJ3I9uwFB71qUHIc1iHz1jkZYbVHC
L6zdAOc9A4YEZxrBhH2cRY9j3pddo+dGtWS6ITsACzWsdTfj3USWcvzQ9sWfH46N7VuoSopjZCLw
9UlXisOxz/CEQ0EPzYP7zcROAaXBXtq2YKp0IpOxS5/TYrSIaT83ApB7GAcfDS10urE9p8itGYfI
Fu+zEBiGKv79QyWT8TZbwsFibsbdY5CND1942ZGoeJr4CN56vBieaD5e/oxzjXk4wTkYge6E6Ohy
l9AMpYkdzZYU+klR7R+Z7grkn6THFdkem83kv1cK/utS8WkGeHUSnuQD2zXshi+srLmBFj9ZvK8D
8ESX44L5bka9zkTFkyzgNmWlalWzfk+TbOhiQtfMyWQTKupazmjylNogODOxyu89IKKafvRUy8CC
VmgQW+cNc+Vq2pjW8bYGJxj7zACqMqGYWlCxMOUZ5nv49n0sLOH7qkbSbbFq223CqGqM9F8kTUXV
wy+ifR0VLe3BGLn2pWHgDHcOwUMiC+UQRajQBOu5kTRtqk8LzqZ70vHjbD3iOjppoiNcyd2zyrZG
fZmaolMbwVogwc/0eGHt8B8GYHE46QKXOWy2xdNh/EdtoYLzoDKi9Xo/5tF5Gb1k2DWAfADslU0K
empJ/hhigARMryfSrLYu/LnMlNrkrR7Z8l1FbSVwOAyxH14jglSamVQYXOo7qISN5p5u59ynQ0KS
hQZVyGqjKmSJYzdRhQsf2oOnB+dsPBFL9pY8I6GW6zJJqBUqtwSn061ZMDD2XbF9We1LSpJYjnaM
yBQXRFse0mx4vi3tS4LH1fOSxDyE/64MLJYAV14OUnsAicawytMRQza1ieQI0VTJV7iel0JfwHEb
MSp+zcB9y5Lx0gbQ5PyBw2haKMYUI7LDyqulhm6z91QIJv8h1F5fKSrr1d0SDZCLC3XArIU1pZIT
ogQWbsmN2D7WdYpryDbjaNjuKKWZFDAftx6GKrKH2Jdna2OnaaroO70QtYfWn5RffNk67ezZV1Fd
7iFob/IeV3vbImAAcR0qq9TcUUJEbU7eoW/BL2AmUHidOhLIXACRwEIbryZjz38fW2Cdz5bRkEVM
m5lMTXlQpvk44bPO35+yOtGjVVYjpCcIAkouFKK5Tb6Mpfm8qjZ/wKI3p4eV6EaLW6nU5M1UcuBT
KVevByOAXgvJ+GMZVnXQhdzhWBXCRwuBphIWQz2fDO8gzxa+5nSZzhYSpnYnO9dNhc4yLj2FAiru
DmJ21AZfXtnrOJGt5Je5GRbFQpY6rKzT5blhfFswg3AOpTqvbKqJ2zbcY3srOfNxotraP1mgxDnu
gm5+K0euhfGgWNlwP7HMWAybTGYWBdpnusnTU/3rwHeJ2fi/AYJ11cp99pE6ccip5SPw8AULEczJ
/aL6/G4HCFlX8ZmCcebGNYV7A9Ke0ArN9RalBdFTTFmVtNa0KExBbR8rtGkydcUauaF8R3b0Vxl3
g/1xtrcew4+cJUKVfM5+6Ila2I2eNuC85KZYbIVHutUbqtYN4XJ2HLP/KcBDThf+Uyt1zXcvl/sw
MoIiWKN3BiyGN2Uzs2fxCvs7Ajagi3CLkNwc3uGxv7mlMB0r0NLabFjIUyvLFcDTqYmN9WVMj3VR
wiENnnz8VZQ5NVDf2IhDHmtytFHXk+3P/1ayt0JY/+eiSaTprIKnscEBnASTqVHqMajXPKr2Eiv7
j/BsxK5EWPKIpkwxmlseeGmrRTlsNcsDYb0vo/Boem+IuzLN0/7VPcg3cv2H/jc86urhtvvHNUkg
Df7EgKvaMnA7sr6ITEcScePuQ3xA5MxyaIp96sQHpr3jiIgYcNh9tDS4bXlEGPnxoNBpOv4CMKKk
Lkd09vlYbQvxnGU1f6/+FZxpaT9WsdD4vsw69rtT4VsBk7TEbcH1ZYQhNZJtg9xWAexy9tmoFOfj
w2GEQOwGPBp91e/BUfA+STYzvQDfoLf3rfM1KhtSkhZtPA4hQEkEazzQeB/cbpZKIyqnDtFE1WPz
BKBCGifg48R8Wu+SyqKunZ5hoknM0KP8GpC1CyQNlMwm1FFj/4SfqpeMLL5jmrZWPJWCYWVjh5wl
ojwS/4jemD4AdXGtjXHfYp1ZSz797Dmpwh+CVK5CZrqVFwEAMY4RYI4QETjHXktAFJrcLx+zfUiT
Uj0wfpkuf8s0Hp3hUTQoUxkPTZbIycjy7Xx6l2jPyjHUKmvJPT72FnJZOE08sdzIeKP9ZfFyKF6b
eAGQd2DMviXolqHTfd7eb9L34p50Z8+CldXyNmXdpYNuXowyI/JDyyWtOSs0Oykk3/9d5oJNhdHX
zVrpT5v+n047JnJwZJRXjqky2jHUdYwjJFB4GN0gGY2+fpcmoiTzO+zddO6cWCUHXJ7lsVKfwZVP
5nVFhX+8Tb6AxlhUKxMyWoPvEWqnlXGnQDB9rSYl1KEhHPoqdOcrakNm8SsUb90/EGrh0oP6jTFA
PmYggGceg1H/wxhmYOzGUrCBaD2WNcTwHENkIZK/xUqNUhgpl/gpSxRuFgmVBrDEY5LYtxKmuZF2
GVmZFiGy8gomPsaDV/r24pGnLnZOHW0lI0peK5BSpSykI2GnqP8+iluMsO6558C6oMUzDP6oUBtm
6LWBxeMAj/9ACMyWR19EHd0jhZM758gYgvnDEQDYxwrvKLP3ToxWdVxM1RaFNIRbpKbdNQDo/tVS
6aE8WCXSDI/e8jAosJ2qaPhzCLTGFbCc7UGCIJ4YNpROw0bBusKOd/APp+kcCZ21gRwMI7lUal7W
OzrFxuZ6+EDsAfaNPIaUJzUu1kq3twysSWaHNlRIhw7ugti2BA5aqnYHmB9ul1p6dB0T7LnTUkXJ
rxUvXvy0iIiMU0OV1P56myiYJA3xMAyLBJJfpL3YnqBGhgFxBQEU01STaU2NFQxRcUR9GNh8+r9x
q12SJ7w7Z+g7+a2262Qs5t5lr6SL9y3OXrUtoD/dKXekdfq43X1FLsMsI3pNyDmmRgg7rVdSzYa/
tXwUpm3IUdLltzp/TXD71WIMYcn6sGr7r+ttvDeXOoJQ6O7cxt6nl7iAflZUhbRRAGrEDefzv96a
PjX3UQkBxxfLKcWoJJdU2I6xv6VQqJC4dMcCWi4vVCMGozyOSO1cP9Q2Uwa6KjRtW0SFgTCeLasg
rFEcn1TzuVci+e0cqBkNvczC6G49WuPMLpPtJWdvLcT1nUUrqfw3QnKwK9DDZhWmCVJCzuyLDFUO
RW8n2sVA+HsG1rIqRac9ZDk+bkIJ9uVffn/b9RxENmU8Sl6aGVtbgeYRCZ+drVO4uw0hL5vu9HCY
HHBGnxrHTZCOXSDHMvLvpHd9KRkpnRfA6gGOI5b0bbCFVhewSlo7p0kpywkzZKafnSmoZLVz79gi
bslbY7RLzAW2ZbsEaF3a1+zxLPDnR1YgustCPaHyRoMhUjpE/qoxrCDeVp6DC2ZaSVw/+2Pkaf1k
rQ/VCoBmwZ66zx8Ou9fZrpdQLrncJglHEAWdLBm2vj3OUgtj0oWyisAU4Ymcs2z5ePZ3jIUv6SBU
w+UB4vHgr/0P2FN280BkQGc8LdAUQwPl/aqj7qjx0DPhPPsq5gkb//Nb3vmCkFp+ljN+XJgEg0TS
PYqRo/ibV3Xt13d84tdE2RZv4tEQA/PMcbxyqSR4ZxFgZvUbpew/HgwNN2PZiKLvenTQCNsoq0sR
opVpL/D0LIubirpvDjc5QQYhuBttVr3+OTcSauVJy7qtksDyjzny09sWs78ma7NutOnnZSuz4r1T
5U+6UBU+xYX3EadLQz4Jqj/Sl8EjxIthqX0UsN4LB1IXIF9uCvBqd4hjRqIeurpv3A9ZeJDWrhJ7
+Vrsgr7PORCWZo4+Zc9Lo586h9BVFaOmJdTShWgDB2gn97GR2MADmWiOoJ8Pc80iz/dSlgKkzGa2
Nb2tQ51FVgNeT/MmR0gf0y6VurIK3rXA3YcAE0wg+ol6UkP0zJRLUeJPEwxCGlrmXjaA+nSaF13F
VMzDQtde85aiQoWzv8sp0MSMgoMG9cqDgFwwpOdJDevP2+MyU/RzdGrFkanlNPU6W6msLPGE6WLX
HJBYkN4U6hIIqIkJo6XIihdQS7R4MutocbVrjgCkTKvd9t/gygW3bm9PZmgTQiKTK1LwAVWoGv7C
M9jRTCjUyXIql5NFPw3k/7MfsSkJ89u9083+YNVmpxKr9SIhxg48aPkvDDjGrSqvB6Ph5kUqAsJY
jfvXRwm5nkHHqzhEU17P+sJsAvjZEUMuHHGJ0xB57eMzbDZ+IGqfyQwdBozCwbphKQR2TYA4w3Zw
v5NqJHECiquoA0VJqQAbFRei5jLaGbGqf2XfjZRYSDyGdlLvbW3fwd7tHWo8E/1QLoU8nE1Bkipr
rn5ZTGcRKOUp/Lbjz4ALGgFaHqABQ1PnBRPlG6prS4D+EdmVMNrY5kqegPCWRAAQHuS1M/CVIrOm
UiLs4dJb89shBt+qzQWrfsPvfKhjNLcQ0TrABtXFU9Jc/77a2wmbY8m9r3DHurAb6ser//CZYsc/
QoWACM3XY7sWotcTSi7t0fX8itsHboISr3C5GrUh3LxmQ5JCNslzbjEurofyRZDekOFP9GrmkwcD
ijkt4ty5Xq5yYvDCpvREUOvSZlXSJFu4d00wDw06ozz1h2Pw8Y34UeCcDgcGNZy3f4QZJgW2M/nJ
RXNe7TXvXBUBVJSp0wZZy/pg/nY9JlrXroVjAKBQ6n3DZE3SL6f7+NUff1ReWWWvg918wdKJ40Ym
Cppk98gI8yXt3nJBy74a2ZlQEyP+duseO9rtRaN975SwswfzHClikskXPY7TWVzar7RP0k75zkpI
Ada5B6m6fdKwi8A/N9sbDU7EtBiyYQKhKhlLJVde4cB7M4r2juLyzd3ew16WzVzuIjFIngRW1vhu
vooOwjvgkzmVOp+nxA0vrm1SfEMCQL26MgIXsO45dZXu+uQFfl+w1xpv2oD9iwNqUE/a2qJOIW67
ceRwBbCE2edeXv9+cJkGsjMVwBR239GadGAlXP39XZzqXEsSN/8iWMOsPtL9zTjnHjsWCAoCvaMX
i3UyKUh1nHr74kgnFEEcpt+R7OnS7NYD3wFgxxq2AAUSH1E/uhzT3h1SjJkVdxZjS1IU/ZxZxeXs
ayNHUNZObdLOqZvWBT2JO9eUphSA5gewt2cv44pqWLBTZLNfOgq9dsHstps3qn93S/OShW4QxGsv
0e/hrEKw3vBkiUw+JqtwjS6xupRrYnEg67hm/vJNkEsrsZjen8IL5pE8rjOsyxTmzW8TsG//DeE8
MjRXBd2oZ5EmoPpTlF81eQbSFoNbD0yJqZnxgRzJfuG/yfGs+Rj+EPv51ErVIpiivFzXHARoVIrp
ZTrwPhGFId4CwQSaQrvHOmxwL2g5SflOEKCxiRD5Ehjf4HpXjQw8c5FmRP+tP5BX7P1T4SG/4jRq
U3tmjVW6ggDk9zUfvesQcN66uu4q4Q1aJB8+Wc0Ge1Rf0EmichB0jxR9qmSyipnDQ1ZRxokeYVTF
cjIoSRwQ+CDxVqGkZgnK+RLrzVtvj/CdxkHYnqZzbfW1v696zAmX1bQYD9CLtsMnj1yemE+LXSka
U23SIMM9Dk3fHVyRLS4cnDDY1hIpjUKJT5dzngVDmJNQlJ06LgSgoV4uWe1uC5vxDZ47BLtbXcRk
fnLRNHDEcnL4fCweXBuUUXiBBxhsHv0FdBDFNADA/i2AbxFEOJuPVdGewrHDzFH6TvHL3K/AlzjI
0TfW9SujTSu2uV/rVs/mA4dKpeKW3utkyu3kX4noxtuaVrBb5peWdp1lwp/8IYHK4Wbcrv/qg6YJ
lHkRoOTnzgrpdjfd3dGwYKLW/TEbH7LNd8+J8z2XEkYc63nwGyp853AKE0oKbniYUctZ8ab4JWKI
W7nkkubEIqYPAByi3bhQUsxx8QE82BDbg/JasYcpvOngxuHMJsigS8uie94HDdSmqTFZkZfu9YwX
J5D25S1/oxMQJ+zXiE1mBGL6AbE8Vfi65QPt06QTbQjWQ03AXMKrqyFNWDSXfdBmZkAZtAf5ikjH
otYN7nb8cuQJKYBp4V5aQrBfTGDmo/3e6dLmnDlGT4lEqRkscSH19GhNCj44/7mPxxhv2RJv6/KG
3m9U0CgOTPHb6+PLhfek/+XAbsUvtLRb/fj9jmFhgjAitK8HWkZwwpK5AW7aF5jJCXtEIuDwUj1Z
m/FiV9XAg2ZDvWKY3t1HJwWVxJuOGJW//RTbiyNzlT+Vb926A2uORVL47hNTr9cnf5iWI9Lmefzk
AX25NPFWAOz2qs6i/iuag2ff3eDMCIF2kAD/8IqDD6QMgDonaCLh8JzbFvsi2qBV7jJmxqaNeWnu
mIrE+H6ddOWWN5bget2qJ2XtCgZeCJvW944gdnPKPceVrAx4K59i0BSah5Q94DHkGKYfMyJHjg7O
19wgEqpCNlptyxIX5OTqVB3PqY4i7/AYUoLsP6EJziopCZ15PnHTGbkm3xBaL9J6T4ErtpaCQzp6
H6PKUn7lVGVq/Y9ioZVEiBwW/jcW4dPBlL1szDH6SzjoplupHouurioJ9ErqgSUJV5mKJViqLHZU
yTkHrIx6OlkNTrFdX2b9hn7eO/ku2jubDfGodLQ/VGtVkdQcWXB9ql5PlJ3cQTC+7giTjK4nsVhL
xNVRNn624y8fIjmcA5yHiOrDeTJ0RCFIH/a2Wf8xTw2mv3JNek+oIYxSXwXp8bicW3BYJOgnpUna
XLHg2SnCcnWgDxw8ZtdtgOfiPYisUn4F+J8DcVWu4wj5Dv+V9l57eZow/CwOBKEZh5fHyaikQI8y
4m6HrjOSmorWqTKuhACHkuILPo1POZPK3jTtJL/Le8vsUGYnHcMqu2V/JmMElMN9AdGNcHr33W7Y
F/2eW2xKq83oHreuDsVhCWVnjnGga6szwMLZlVmrmPgpAYxbsudbpIx/OLgEW7v3/X377ulTMkjW
kKECRTEcWP9MA+7q872fH3XjPGe0SdzJH7hkPK5EOBEOhsrZoWphJXpSw5opbW0nwDS+8pVCSN5Z
RuohI9QQR4oMGLu2ToOY7n+wts5c9OsufwFcUh+VzwNVdkXM6Z2ML+HGGFAUsNzdNzokPLxUl8wb
gLByAyYjY7B9QPr0RDIHaKjcLRLyWekMnbQ0g7YRpKVIZuihkWsQMfhKaF20laQW2B9KvHpZWl2I
VxTEVWwfDp9xoNJZWOVeXfWJCMMkx9TwVpI9u7OBtI4vF3N1Xd3I+bqE483ApWw5RaBIPGsv890+
a0DqNsAY0g313krhDZ/QK8VRMc/iToSeayK7keJAIcUNmcbyW+GtKny0jc9x7LdmxTfE8Hg9Z9xe
nH4BOqDC8ryr3Tir4JjztV3kFaTU6QJSDHkEL88eG8X+N2Mblqh4GlntBw1dKJd3yXGFcLqfRNjS
T7ReWne7yAzX7MZSa+d8etSQm5B8KHwoW7355EH2EJu8l1+Bs45qBn71W9ce0f31Z0W0tiHk1vFD
w9s+5AjNZuojIsewxvAMffVTanxY0GECRzQMpwvjEBTAzuvcXljoeec45u5w1DanZKEDutJHMaTO
xlIc7lB0FUD9YSxcGjvqX2MikguSH4gJivum9/9rs7RAaaGjI/uirpgnEyLmLP99DuHyeIF4kY2w
1IGshIdiowQljQ9z9lNxeac6Arpza8aIjwhiHloETTNvA/sWh4KBvKUk7nYRI2N0A89ODe9NJPZF
Xn1Tznn1AIRztmYDPqlv4aXFqDDKNlMe1BS4/TJizBwszLLt2am/s5AfYu4rvV6S5l5AgyvKU5i7
4UW7c2d/U58UXBBsopr4sIv+Mh+u3sKtY48nQDZQDN/NYBe+RbKwBf+ibQvd2IFy00yxBf4VB7jX
5XizjyjgPH2EEZvqGej98lyUv6qWPNb86FwvvFihBFF7QHO+paPe4dcyrWvotGxD3Y2oB7RH0DGg
jourONG/4nvupENaSfQS9Sa9zLM6EsF03mrDRf1pLg+UpU9z/OfG73KISliQVeJeq+DBMTFvjpsO
p9M0x94kXZ7NkXYcrNjykeV/R+0gpMM8KT/wJJIHk4rXBBYBwcc5ulfpLXMQwPTDkhoifkuSHb2Q
Yud5ordUnGJj9O/uL9Q3WYgnpOYYY4JXKfxW0sZR2sKwTVHCITkrWQqP6tkpg/O7tcpREunHTRhY
+VQdxMsTmdafE0oJ8Xdeh+sMqV7AcMqD79gERQ/0kWn2JK/ApVgR7e2d+jUVXDpO7A4VKKWRx4Y0
5kIkjCUMyup2Bl7AQNkqc+JQAbpe889p7SS8hLGJReRFsHXrqGiPSEWB6MH8gFBNP3qtMqnbuaal
d2IRRqOx/wX8MxPe3frQ/1Ti+s5mfyDI7TqtxfubcDdePJbjg8/l5fxEBsTkpJ114WdMXdN7qUy9
wEAZwbseEJ8dKEkDYv7ARn8HzUofHIgzwWTBFw+DmaRo1Yhqbazac/rbp+H+4W3EPEriQU+aGbE5
ZW4nIaRFy9vTgrTcscYYyOPSjhWtrKAOttUU2n1gI7wXmHyKvJk+IIA6Pj6YGzi6TZvmowrjHVF2
jEKwQAqXNHqTVNLtnY4YAUsDLeAIHIHy0HFyEtzje4N1NcNrMLhR4Znb9Nebf1eMOOxMtt4LYgLP
nExryOOVXoFH83EF2Zj4YVMMSBcwCtjwYrnLZrzEe+mbKOnvLHlv+Lbn6NaBJwKc3Qy0AXdCq+6i
ME5VNXIeuKaTO1WREYQt6Ki5iQVJeVHvyIj6kL+CpZxz/AOhOJw7dRhA3gerw0KRh89KpnIUD0Ci
lRAj1dPsjfkU8NnbYGDJAdXH22/X7u1a8wdkfx77OUKSE5tWnoKaUnE6Wh7YD7mQarsTlg54q9MS
QWgzaIqDF+bnmM9N5Tz08DUa9109kEdP4g6h4+CQavB9brBRBst3zbqpOrAVaeVkLiK4h4JIh8Sa
BSKRtlKPfj4Yc065KUUCBVrXVU8RZPcHwsl0SO6vaY8+TlNoqPTTN9YzVTuQmH6xoN0NVOB3hfQz
zbRW9DhJWZ9I6YqgKjbBuBMs4S10GoWfXpIw2hB6cRtoAV5OHwoFIIlHc5wbvTAJ4z8dwV0tsuSA
2VFWPc6KTAiqnvhJh9jLfYe0DZCa1FTockvsOjwEgN2QoMaLBe7gom6twpGZhQfsSNNv12f+KD02
XsupmI6dXJR2fbxvkhW69gqvt7WvOFKH9Q8ziLmwTg7uUjmQ6gJv9hPvYQ2gMVvzIlyokpg1ylv3
hBxykiwNeSyFS7KexX+D8XFIlJVPFVsf5EpJRhjYN+X+xZVE0Q7kGT9apsfqXq3rbRhqMDBBxPtq
VxD2ZoECbFwduKTcrBQ8MaOo/wM3AlN+Qwdb+hkxd/Tciub7lPg8kTRb5GftHG8TT4ceQkg+SfLa
jSqkLSKSSCRCOIoCyMSqEX6Y2D9YXoG8q9WVmf9z9ST3iYb0sW2mvCdvBbSejclEWbp76q65jXez
/QRgb5Boiqr8Ehedk9UkHUp+jABACOmDodmHEPt2TF0QSJ5Z2+fXVkBJbRrya7ZxUNNa/nlBH0/K
L7GNL9su3hYXfQ0QA+8JlggdkTmdb/LRtBXRF1LQpsgmhsLYTcJOl8tMVEVstFND9KMIGHrGF//X
vBd6y62hMa9PjoyWZCP7/8SGt/b/1cOpgpfbLAnpW3hXSOSCJhfyDW6X99HBhl1jPOhvN3kXj01X
v1QO2ZJmA8zV93JEB83Oc3Rm+pK6jB7RlFcu/RSTCaBmMIt0sSfV//8yxGkNNRXs522cHLzjE/Da
+J9CQHx1ofKAIozpYhkmteM+f/euzHRYqLDFxlcchVCZ6KEpDxgmG0exrzqiDcujtJUTthuEv6NY
uu0JLRYUyI2YCDP/QVAnPfbyIcJD4FbDEAqBjDVQy+UYhniQX3PgD3T23/8THzFmmiLBayb8AZvj
Ay0mmVLW4AO+EpaZQcDqd74Lu1rNBEmJd98r/63acjacS2ftJsd5ogLl/2F+U/2k763WrRZXAE+Z
QBVSWsQXC7n7U1xjEBFqbLHEnWirALvfzTvXX44x8tGDTtyt15HXZJhURoXG4kON5fauSph65HU3
LEuXX2U2Rv4vVzShI27v7UR8CoNq+ICNXOQ/WteaJu4vP/lzrUyzesxZiyQXnTfpnQ1SFFqTiInC
9K3irBlkUW/tqSKO2cdctJNnhd0hmhsAZDG8zTPuReZeKTEljaG51TEjLPEKt34Q0hRlIaIaPm8C
Jq5rpBttkbPCmnqfdKZVfjySa/gPVDMkwxpn9rN2bKCWVj5YCG1x4jfn21EpOY8infeNjy3fNm1k
6t0HfVwqsBAi//lXc9mHdlUXgqz3gzeAjni5XQ97+ogW6GSyQ+wUd0SQCjwVjum6IXeYLAH578OT
OLabfb+92g4Vrikb0XoTE7tt+H+6uL3yyYKxFTiFUKSjDzZmQIh34yx/kLQQE6wdmIYVy3VGXjyY
aa965dNRvRv78dDUvSzxpQPK61wXENJkFLzBAECc9GEQaykX1o2aYA92UapK/7OEM6fJL4dZYT+5
1+owvLKsnknVVIEJ+1ndoH5ntwgxAA/P1DyWpThBY+45L0AIdHBVUsYG+VrSOpjO4BozFjVG+lJ5
5IaYqKcCoNmEyp2yUH0Pc5I7d7j3Eolx32NhXh93KHoe5TqSZ/LzBAhHYtGD1rZk5RbgN8BKUJ8m
r4r/GPG2wzkMFrQ5rEa3P3zHW5XlPyoEW9b7fqhCenD5yFSZ+zEwB09GVtl8moZj4DJejkKEq8Bm
ndjOdDYO+jgz7wtlplyeojmmmVBkfyOIxGOFmVWcilpcaFo4Lgu+QJs/eIZ7/KynriNP4WX0RQR3
J/SfY0DY30EkXTx71K5a5ESuLl/IkSR2fS1DozUvvxzlTFvtCgCktQwK8/uxe8PfcrByHTKl+3SU
x8mZuHMKpEjL1SYzzZbt+Ocp7V5XdLFn6mup9XqiEzRCDHrkiZGszkWbJX4ofRaNKH+PuC//9b/h
50XxkxZevQNHKNpROEpqxAF/gRce73u4wCqMnWokW/eOumdL/IYxrf/BXQk9JFWjJE8/oXnna0S4
aCPK980m8/wTyHVx90ka38LGQgZfEH+Be9Z6Acx8ReJAWLZ26WkE2/qbmZLlwIGp/kFB0BafOgSM
lXNtH2SpWxH2kaXYD0zA4wAXvaptFiDLO0dnPRl9cfIZzMk0di3YnNaTGG3fE+O+I40uMp6wZGJo
j9/qzfFy1eARR3MG6IFFsCpXnCS7dOun3onPXrsHVbSKv7vKx4ZMiurXyAEfSSaPV5vt/oODa9cD
jptNSPiDYe4VqXojGb+bKlRB+oW1JktoDdiZePIV2drJG60zZsbZNdjFn2UQkkWfwBIOZve4nXoj
kWLDKWsqjLQ8wfl3nn6cJz9tmufXA9/JBxYN9GeubK0Fb7fwtVGiVkbwOmxb2J6hQpwU5hTJxmTk
vssdjEtJVSPBNWAkWrwDTymRW0Vha9Bz1Ydzs3IaGgTm0tqm07Gut+73/GjE31eEf5kbuIi5eUGX
OH1vpBEpljr/SBZ/3LmDnwCYgSdpXhuNWmRzU/GBx8RvoUDTUDtbZUemkuYCqjvA8RxiIjtL+GBN
4ibv7W7s+1eH4UMozxwPovCjJSDqzGnGb3ceSW86Mk6aprYUkm9PtgtNNh0HyCQznL7lCplW3PkP
VV1+YA4Tnj3+kGTayxyrhe8ak65CPbFE/10NM3JekEHkHhqeVJRL4sv8evIw+3F1nGzg+gtERff0
1XkmQpzmtX75egY8AQ4FPLlaOHrx29RgFNJXqN6lgxRglewAZOIaPy64OkWf5GbTLfuWLTjGtV/D
yLz/WG5KYzRHHhKL/QXw8kWPbejirfhGwcj6BcJRXCYTS5pZpatW8Qwg5+4BqsBeAKpyqNnFvged
ppizDip4bgjCqX18eCiUofajvWYBYuaeW79fHdLOCendLj0alUQVgfnB4mI3q4Z5gZ5rAHb7ERL6
Z3lcYz7oVki2pe2upGomA7gx9Ov2Lqo3WRB2ynvGBZ5/rsJdM49VC/M8aINSMPBWR55F1yb7IJ8a
dp67HtxCDJuOVtWczEuWnnkuC5gV6XCcxYBgOorMjeY7DeXUlLBe/BMpmxx5Oo3QcVQfIT+k9N3e
W7UZ/j61jDBzl0CFtHfKzcij84jcmlyNBoFCLaZ8g7hDyU0hDC/C+txvbckX4vtbxwVXyhmHtwEP
9+PK4+G6C0HISbumTUYWLpGRBb6giJYBCc/RB8V9cL3EyfXfATodcAwBbHaQlW5P0d0mo8qwUcek
0dvkDYS8u1wGEq95t1pdNOIXjCLK6DVElXUbRl6KzYQv8dwtGsIj7AjyTDEFRVsqZRnQOEjDicHd
kr3GhSEjXEtNTmXUP1WSOMz5z13ZoIcRSvJv5XDyjKzIGfXqRhFXybNNyH3qIJgWqpjszot0h6Df
0pGuQjz0Ogw3qybbdF5jyYZvkZXsICRqkCIzs8FxZdplnTaCg+wwm6D2PlEn9CXjAj6Ja4MykupE
er37jHN41RNVcYOBaKZUxVnGJ4tziRFAgB07AA1MWvRCxI+tXx8Ho+t89gMH4iLz5wmPs0gz0Qrp
ZJOGrueoVIO0lgCQTbjMlEsYjBLV9jTs4yQFPoB7xoGNkeV3qR93iHftUT/iv5T0znM5oVuPP1Dm
Duhsex5ActzEfoFdyuP16S+bQaNddnc10nl3vQL0mOeuH3yEGppFLuoXohnPf9LIYIrRRw7gBQSr
2AdSaxMpQibscKZvs1eMa5bUp4Y7LQDGR+RwRQvGy288Ttx2lyplMAT9+flXgv7jbgnzkeefpcrc
u+ahfg/brrSRBqKHCBVe/X1ATMOUfnqnCRzZwA7IKh08RYK+jI9/m6S9fa/GyOvUlMBUR9pCKRkD
9hXNmZKukFzpB1ZV83YWMwN2rIq8ycYRu9AF9s+2LKOksMojgKdwagN9T2Cmj7OIgvNP5uqa7Hwk
4aORJAVmHncXZXIEzZhGtlDYb8PKPI7HvxXTrfE0829MikX5RKuMK5y68jANJc5Sz7YdGGaP2F0p
pmG2DuMAbGtPohdDgabM5VbFEGq1IXvn9dPSEys4Jp4s+YgHkv8s2YhaPlcse0LCUh1FOY9t5gJw
cDDVqNIqHF5zlCvXsKyD7/E9dIUa5fl1Xz7Z262NrIRkWV7b5lEKLcZ2qmD32v4kEtgb/P0Gt+GF
51EQ24dIB4eDxuTObQPs7oyVUNRcUDS9bYhhF3kC9o1vnzXn1B52KN8J80L9TdsvdG4eY4yx0fUI
jIiS9lc4Xvm0kCKJRQkIqWO9cYT7Na28rRynJuoq8q2G7ItQnsXO8DLecMLJfVRUW3GwtwpuzgBB
6c16v7WU4gejNo2N2Wp9THb+FjurSH8081DGckcoPm/yp2NeIdita56jDguD2zpqGoW4CFyA8f8i
wrzatSjZW7muAeWRu+kf0+qHa7RVlmnzVrRer8z9kTRuS5s0JqfJA7FqZLit5pTefFV+VTjc3hUi
99uVkhsH1AsD0ZLaJq5oSeD5qbCVEOnNtg4K8LvVDJHg4Tg1XDXeGgP9aBsrI64ei2lrKBMIf2iH
PnhGq567+Su/zCvBn2/3+DvrLYIXSTGFAMcIsSR7SUIvDQEkfZiTmjo3+RLhCrIF4DlgG+KftoXS
lqXNj3xacVGUY7EB8qopRSlc6D7wiJWsqocRsAyCEFXV6fMCu+VbbONX0BIb2bvHjII4mS2d69+6
oTP+5PytOv576yP3wsacdvuQENpXkGLk3O+IFwhdzEXXsfug0/1BlCYOxBhbARwob2p0drSr0Mr9
cTfu1/y85faYymBj3zUSg7DQLMYleT+ct7zrBBfiUgt+Pdp+Z4st2lwJXfZxBJiTKVoXYKjk29IC
B7dP7F2aEpUg/8a6qfVO70woN648602olXsB4ayVsVTI0zoXgvyTtfWAjGzyMPcSjaShVXSvFa1S
oF7O5A3YRFd6EpnYpDsBBtDpIFiZNBpjQ/xPeOCVcgdf01jbiRYZg2bJvLpFmd0cbNsAAwvkspvN
Vgrlkx8kJccGdqzLbnry7mRXcxqtDURAl9beB3JfxWT4ge6ocZsfJAcKF3dQrBvgwFI8Idn64IEM
KSzdOB9bz0wBfNRywwl8+LT02DDTF1scGfujCDBayAEpS1XMIMcFTEFnD1zAMZWWmSuaAVsLTAva
3qVcXRYaqtOzwcO/dNeMyqk1Ohs7HoehWT79QGg9rWwSq28yRrmHfymR+wquRAskxcY1F+ghHf35
/zJ2SZ4p/ekicsd4u5P7E6hwfmaLY9KvOBItb7mt0nPBPXQWIAPXdL58uCIq8KNEdgR2hbyCqNUk
vKzjuTAbfhdyV7xshiFcYkUGVb/XyJQXYXMnYrRdCtrnklEvPrQHuRQoUD46cUgSKg+2u1mdZpbW
h1r4xbOgobNkEABTUTzYtXryV9j0UhDc4+oZ/ND3dauplZp8Hr4es3vT/qQndxQjp893hcxFZ7bd
+EZtV76+FFYGa5p3rXAGEgCiCZ9kz7XiqP3WnZuBLfsP9YLyvLbVV3uYNlFZhyz1q2IVPHChHJ5p
JLhwHPGbFNobhUvR4hjq1mRKRmS6yH5blAqCrsX8tGob6WcZ8HFi3Q4rtRx+zLxD/cf43kAy9yKR
Nz1/f93W1CYY8OjysmsqKG9alRLKz00MsI33lbExPDgPR4/KAeNpS3nZGKgFZI3kceGuSBct/ISe
UAKIz13P0+XacMFipXl5ehlLw+Frdnb3psh/6xY6b74crWRXYtM/DE7RiFF8/QMNcN9SuEZ6W9eo
hDmpfUV30h080Ckan4ZqXYbpH8Yx06nHpUl3mTb1ILTbhmYvHXvVtxeNVBpK4OFRZVtppRCDk1OW
htmv6MTeeD25Q5JhTkDkBVa0PiewDzON03HJtku35dEptPugwXcSCQQLcWOU04JLEP8EHOxdK8ij
6nQP6++xwtn1Bjuri8SIdN/bKnb1xy4WvKlI7q8yFrrgUXBSH5L12iWAQU1m5v0kACfSYxZ8bZQM
R3DCi3DbZ1jVAEyzuWtVgUlUQnzw+T/ETltrcjpWJZ68D4r+aTDXqCJOmWefDlV9qlNUaCIoe8YT
o+TQHa0U39CO9/pcpqXLQV5m08P8hsmkXYVt1akwU74FaAMyNJMQqmNWMIr37pioMM8NLxg3dU4k
K6xNzyj5Us9o7uOuLiHo5MwIS75xRP0HSycs0G2ZsSu9sF4FAN39fTtpb9x5BY/QIbMaWDAbst55
gVqaZFNTljdTzA5ko41HE81Ji1gjW/XQXUBiLQmJAVUeighK/2tGk1L/oTsN2OooF1B+11UN4q7w
MW4P/aSLCQS+LAUQf59z/HHMWf2ZzQNmlcWxbjwRS8C2Ko0+cWhZDqetR32nvTk4jLxCVTH2Vi1V
avtIxQ8EbnWDAJ73aVMvIojG3o/jWEAng75F4fKU+jnQvN9BCd9N/ZNXN8mq44iSgb1aAaOrcOnD
hwhC+CZ2aC5DgLLTW/xNiWRcig9kGNWovjx17MGLfBGF7pKCh31KE3M2cjoxTmOJ4YDJxHIui1kr
LA6oPUc+/GwoYb//D7KQscTdtjiWFHKIZ0nh/vwuq8RhX4tRXTKrto2n7o5+UeDNxluaWNPfWwsy
S96CUfK29dtt3R0AbhuRrdDWfIKWYezlRYlX3lJVpEixvUwP2FoW19SXyyfujyJBEYgfS9tR2XMi
3Q+A18HJs9z5bjDce+2uLNPaYHppZogO73dmvFknc3HbcLGA0wYdf69rVtvrpPnL1g2TElveVyFx
Ft9MqaGOF/BFVwFF9kGixWsvtzebkoCf5k29Mywj0fZ6TFrhEIohaCiVvoJU2Iogz47MmK6eaQZ4
FBXzkehHKkffD/igoZhdZa8FvTRrIpBo0xUtRxs18WFRj7cPMUjWy8bKT73OJdJGVmdTvI4fohZ0
ikEWI1S0JVdHRtXDTJsY+6Y/G+B7SLWGeEA2+s7VF3vXh+v1q7saX0txI1OAOOAcEhlEXHd7zUFt
YCl9K8y7kBXrwT8LUJq8H9k9Gm747t7hJWiFJn6hMJUH1vyktRKVN64hs+Abc+RS+fE/qa8a1gGv
k38Xt6qtodvQdEH084C9LPdwUSIieYK0PngQ9IXKX587XiuJpgLLdIknM+kqeuv0//c7wYf8at4I
2PIoWxjc+1DlUzrilPQgF3o2P4CQ73UIJNM/W7q64rGntulCu6VS4HpudXP5vvessqgCOmWI0X3Y
Idrmt2JKgkUD8407g9qqBESm7ABdut+CNXGg5GwHfBIxLga7qfemMk6Kmi5t6bhbLmRE+y3bh8Qb
vAvcvNx9Oi5y8+O0wORTYzP7jvQf4kqslVMJB0hmv9te9qNtTTXfJlv0FoWvRNxrj9polu8gKVa/
pLvTTbVn5BC7OgO8cKIKXFki/q5VWU0V7LYkEaxLrxQsGuNwBF8JlonICvrTdvxiZPqcLLmKjUb6
HoQURRfQFyGW3+2t0M4F56Ie6qPXwPHtPFSChXl/pswGPfH37hkb06DxZ0hvnD2dAvCYjk5ZXf/M
6NuVCuL3aMKVhmkei1TWuG/DPiQQC0XnOC3sgWsP1NJwNoANzcm3EYrur8d8DjEHTSJsOiN64Zln
BoMv4DeoY90uYud7j+2SeJdW87mAWjA4egUzRWtFpaFpstVuLhJzVnDKmSbfSQ+JpOYoMw1j5hao
hqIxbpqM5ux5CkbAgLqV9ohKwKR7CQdkOmDJIh7eaXIguDVcuccsvAOJngEYmHgZGJZwRvBMlQ3e
PpQkZHeX9twtBjx8hoRv9+bwBuunNJrjXs0aQVLWmLS7hzti2w37hOi9UlJa7MnGW5KG9Wc62NkF
fG2qDnD14qYn9lJvQKRzsOP0hhwt20LY85pB8Ceh2JSFEVd+5ufGFs/EqbysAY3xfaiaxtH/oz71
oG7HHwS2Nut3WkIvwVVxjhHF3WY6yVlBtDb78CXhqcDOzqlBjhEFIKzisF1V92bReor3IQg04n6t
jIXDxC8emd1s7SoCa9WnKHbX2QOSZuwwEeD03XynBNiWdsy4EQArkZTVLekFKHrL7CT+SuO0YXrH
hXRvAWBLT7vyIzfmJnb1zNWuTx63yHT5XziHi2vTo6omGPK0Bq08IRnxMOitbrsTexP1erA9axM9
fmPqjpdhWiE83gJoJPsKGQ69+2UsS7sIvBCP6t5Xrh2EolKzf1O2dYaxeQ+AYZ5WwJWrvd3TTvQK
95JHG2G6ld9qSguqcqd4ge9Llz8b3sqg8ofnHvV+PUdn7X7LWhoZWpsd0JtM7AlTzzsbjmV/Rpl8
XiqhPQJDPMeo/IroV1p2LGw5dV4FEfgbn5pqtFv4Cz53wcSCqeA7il0AXM8bf9Foypa00DmlLPeC
3eLEO3o+fxD7NFizkczjZ6+y75A/tojzTLddGqadCRvFwFfKrD80O7nfzFTGUuYhNNK5ypExm5Vu
j5aamti0AFMgMQGTHcETGTHJTOW3SNsbVhA9vgbnmmcoHHQo7bW/HBsE173lVRr3JNwxzwzceL9c
QfBVYJGavRWtSqp27S3dT33dN+TTE5lErBhPhd55uqlXCq3HiSXn9SzwiBXfw3KUXWYNow+Ywkib
hYn6PTcK8LBSsORbspli+lsJjN5HCBfrJ87YVxvbRM9cN9Y2ZIBqYwTvbklm5mDAKPsxk44xDlHJ
F4Rm4mOKgW0jjGs2zkj/2glJ4GT3kblkWaFZrQxaLpYKaEhgdJhO+8KbIiToYXNIEVX19iQ0YMtK
6OSDir6fdcdtYLJrfSOOJV8tVucLyL/586kdIDaqa0yhqm6TQmQ0Kd66wH446aT6zX5bwWS7WtFA
6Z4QFYwEjFdOnZXG4AJal56Ope8IJdiEWfCoiWDTcUIvhISFkenfbv0JXSD81HPZZIZb4s+UczF/
IOmJudov5a1uJ3RTLDC1dnC6eLYso/JIXwZMse9YI5DWLCsxmsA3W7OJDsje1UPsynp+Dsrausfq
3AxqGgNFTmuxqrKu3O0CPMbLpRdSU6X/ZvAAE5HxxOhHhMt1bU8eHY6wnyaaAiAs4WDGvbPjR53U
9fLFGzd94/DOIVqfBO23LFifBhrvuIfUXquT5ydRpIOoLkryL3pci/ad3vqaDorNdVW3xIDn38Zd
83XO1B0AkZOm+gbweBrlkL1ISqRyOqZNNsx57ga1xHh7zRXG1MAkC8bQ/1N5ohXmX6UrQOiiNmUs
RPutPFCA9DuYqyUlPK8ZdLcBBWkjFSwuJVkGrbSZrTKqWazSMrxLFALlusvNBFjbJVv5BafL8NO5
x++a31+wW9OcQka2QHRmgtwzfwM9ktiqXJZas33RNdGftQXfggg6DyJhNh4RYiPFwGyk6GPVS/m7
ijyPsWF08uwOyL4E94ehJziJW76cTR5T+O8ebBvB7QNKmWzssuQJnrHSuzRnUWWapc6FfzAjlCCp
Pk7U0a6gF39fFFlCSCLAgXPPb5cBWvuqUWYvrzaMYyNl0XtuMcC/8bgBqiUv3Z7yzFvGACDS+Hsk
MCXxYt8eny3MXh3I4w6789WnECxY1pyvbp2SrN41dYEMPLXLEZp5NmtsCLNzLNWbc7+gqaxmmrFe
+pC0Hxc0VV2J4W8/swlf7tDDixZNhCXmWmRmWTmlKxEC39abP6alIoLzk2Qs3l0Ld3QMiY3c1hsk
Dhnc4D7+n3u5NVVhcSAZwx4Tk64RYafXP1RTrZrUBn4T+yPxksJNcF8deFpDegBtCT3zYcQB85KV
gifhyCUYzjHid3KAYmSUh5BQFyJdhEN2YL46pgklYWvvgi331FT3a9H+6WnXK0NIQWlF6WyTwXMt
j1iF/IlRM+ZpmKL3tYn4/wBqKc2IcdEdZNuh2tRDzgCsllcJqxpTaSKLi5KpnCr23jftZSQzWySk
TD5tv2FwOLTegZde/7T9pnviRimN2MVpp94qW1c5r1JFrqkYGdDgmrsd/dOKCbh82mhxXd3b/rOs
EW5ISUfJLqcmS+auUL7mc68cDnnJmWg1N24t+129fdDMG7aCFTefD3l4xe4bpuXkG52qCC0t6QYN
8pF3fk/rLxyv0d+pGuWBbDo1xf8vQVgWE6WTvbrSB6lPZNjzBxuHwMalcdwIpvnSTWRZaEF4yLm7
FTlRZuCC/WKSgw1qQqt01qoDN7/h9BoSrUsO9V6uo+J9e8MS/x/mINMWfEg47DuyOwH+dLvtnJZQ
NZxZfBpVlOkEjatDlWMlc77V+XvbiUaK3KOTcM/H78Bu+eFIx0mA+9dc9zCAIeDJODDTVWiyCuge
LLIdsKMYIkrMCXJ9qh9KoXtM3ra1/ALTF06fEkEbefA9w/6o07OPt5AaO8aDVGV9pfMJxoS+bhGY
Fpm3B8homPTimqA9x9ouV6ZhUN42TrU1ekBmLZ3F9sQVKr1PY0aVAu9z0YxzIgSGynYeWY9NKbDS
FzB1+t4/t0i3DApughQv7ymdyy6SJWOvZqQuQNb6Fffnuz8u83oedfm0xMFqJfIMs9cY9UORAQiW
4qdLpYvyZbr5OAF7j1AgKjIesI6LnZcLhZ0AuoTKwb2XXjIl6FqOFwmlNlre+Y32+5NJRsNfmPYg
OUAJR6IrAh8CNln7n9apVsblegWc4YJfk6CllIMwm1agbn0bfMwnLnUgxgdibW39PrcHFGVUz2qe
CIx0HDFoUTOKjW8r92Hc8jA3wD1nwDVMSDpIM4QSYUdDODRLPujFwpK9vSWuVmM7vVnf6Fb233Qw
w21lLILoxBpMuHIcsRbeg2HT4cPJQWlRS+yhVdRArvYuKfcr5bpYH5H2muRN79SckSVBgV2aPgTP
bjqSRzFUWd5uz/3tEbwyaiuI4LHre3nxYBNf2O6ZUJmRuUe3ML1rv/1x45sh4Xh7ejp6cZpYfmPg
mbHvk+6plVBF4AE+wn88PH/IKCQWDvo2EpC0tHt02mA1OAOCMyaxeCX8e3vDp9cYOHa9Z/bA/9jI
cx0pkEnzHbrwR7h0aCuLorCy8txziQvNN/P/9LV2qw9klI9Mc960Byt+9+hSLCWuwqJcTz3iqZMZ
lRLf2RDrYTXmgIN8lRyNauLZ60McwbZdekejE2IXBQBELz3JCvNmdkDhxHhgJlrMLS78VdBmRk1h
rb1PYTQ8vDBoP6tmJu1evSqUywccBcFAyGsl6O5pwJVst/nY5a5SQfbXVkmelw1NboAlIiSDYPCx
/VIZbeOzrnD0Ab7Jb/vAqQvDifAgtUZg++396kUK25qgoYLhy7Px3c553GHFHV6ridxcvTo476s9
hU7VyzjPHYQleB/7djLEHU8rOgj2Y46pqVWVR+Zlcjo4DtXltLxIuZmPYmsBitsyPTRaBdN2gJCr
qmoxBfUTPbfbhTO5rpuJatTWwqkMsjF0Ewzy8Tnp9FFpCCk0wh62fuu/Cnls0hKYkCNC9+98Ocqd
tZvTzJkNf4q0Bit4CpsRnaLdLCcXoVytrhQ6aVO5rb5ck+ExnWFkIJ20IYDBXZgokMUoU74zK7Sv
6YlrNgQG2STqLK6l5Mk7VVGe0wDEMZeaA/Vc+eb2nB8u5cJStM/bHfissvALjpS7BMaL7wAdBIv9
frceMPWKKxNDlEOJ19yu06L3W60OUHrFTaaoIVX292k0rV8/OIkLRWYPIwb2FECeskPnk3FpwO4B
YgJK9h0pFgiyyR6ruVcxnXDnTcHl4F54c2nAInR6x058B+d6/tJ2r0bLBFc9iejG0hMbI9AjOuun
ORdArNlAZ9PInpE14BR3PlJydfBCTGrT+0Hh3Ni/PIy2KMSh14fBhI/eLQfrhIcHt34OkM33FTrV
9tk1a+/Ql/cDuDfpnURBNPw8AHFcISoq3IUz+p/3IQppSriAkIj7QU5lpmgO7XOnn/QC1jSoasc4
CvPuD7h4EIqj6r/+niYY30mrHFI5ze9X3F60D2ep0eYXye22tib1NRchnlZaNXMBv2qIVwA+ZClg
tVPJDupIHjSKPd+8LL/XtIlYPgKSS7Oi0mqW9Y5mk+q5iYVlS/1f6mLlYra3xEq719f3+Y7KgfNT
1FoReAS6YrkPtsMWMozUi+Y5hQLOiZoVzKfCtk5w5N9uSg+CnMDty16l5FP/37W1xrG5VBQL/P0q
0QvI/82SNOsICPA2abDdjKK6Ou5w6K2XCJIjTEIKrUMxjQDz1EQh/DNzSe/aPYoiMXirIudr0U4T
DvpglA676w44exLl9YNwrU5+HdfeYkGmJdAJwMmiB1IBCWtntgtjLDeYlEI3tQ73JXpGA6fa5nZd
Z+NyQvO0DVnE5m6NYGVK7ND8DuH4/KH2eSSIlepRsSvdtXH4D+Y+93ePfbBhbJ6Lf/lMG70PnQqw
uuqr5F3jOEaHjkA8KblXR1lz+wEurhR5wdR5LRfuFxbiKGayBpmAASmySmkOcAky4J9igcBw6IdW
FCo0ZlkFI9BDEDsM/dtStVnMdRgH0T3bvZKUmJ5yNdzGFdge25XMylG+6eQ3dSr18ysa+pDvGjsv
zxgu3IoXflq2BlrmjdGbCxNwhQSyX5kxMiYBmTRHfVauqBaRfqp5EWiwL6CG176lBLQA8AlR0/My
a73qnKcpbhuClIE7+K804609J7E61lD8FR7GhSWQp9HvH7e0qxm8s7DxLkDy02g2E591m1VPkjne
nA5Fs/3Jcygf8RXleuLp3/mM136mjS/RrNVr72R41tsJOeMgBVEHb2mc8HonKEzFSSvhXwC9VBSs
xpNT74+FVs5HfK3GeCghaKWX/Hw8h+swbMa2xKIjXEM5O7lKHoGXRHFTTLfhEU4id4pPpcQ9+3O8
PRSAQKavSYd9ZynR5Sjh2QVj3WPfE5A+GnYVSqsa7kQPBVBqh0hEFHy8LPpPauP++dGx5MY5V2l5
tGZFAsZboPr9uaDeFna4LlCh9Pp56ea+0CMee1CdJMIg5QSnANAiMjtGSFGHg8y1qK5cDADQdmrC
PMVOnVjizgrkAG1Do3eqWnK+sr9cXI4830FEA4XJvdCI9d+u65b7Gls+7g+B5ivpdZV3gmw/wgvD
TxQZAIFnrsmQeCDgWeLpLdMtvr1mAD6lABYcLobxojrS27khEYn3ZHd4viPYtuSnRswVUoVkzgCj
FW/fiB6D58sw/jfaM0unYvG96/tZqMk0OHLr/8Dkar+Wz9siGJYsc+u78o5v/m1emYBAoFpRMgxY
dWT5bt+r8qx+DuLkW9xVyih3pvc9osifosuc3RaFLGcudviWK4FBilt24A9WyozwvM6NahfqoC5H
35EhB6fKrNd2BIipxCAZ2tUTrFKMkYEL/sHQlKZFgRdwFbZmxF2MJqh5enPUOFCoA54phD7wsEZi
p6HsZGri9NjOLf2qsufMqvB+peYe15yO8kHLT1kIvQdzC57fWoVPwMQpakUlLhX9txjA8hAfZyqw
3VOGPUaxfk7q/aS+sYoHDKnu6iX+wSIzZS7T/i+HX6FN594S0Z/RuILp2QtqTXACpkTAW2buR7j6
s9Jvaezb20qUZ2iK0MgPH5PDcb29GPL1CR7eq7yV0erqh3KFApwWaAV3dxKTVMt8Ws2WwmerMXvJ
S8SICSSFMk++WMkPw9Q592p8Gslqd8vkVz5iI8l0BCONMU3g9EMulC0pedtyrDot9G1E5f2wrugP
dEH7bAErKqNUbnCY2ybd6TeOUatR6xj8eiuPHi3L05bivnm544Ks0+PrUPr8FGsva0uHOQq0noYB
QAk0Dpq1KR3z2hEpWilK858YHmO8jUqGHTQOnz2J880bEnwYrNphJhbBU7ibKVIWFPO9lsw+21SU
IOBcUcaQSdOmuUBOmZWD3rjbTMyhv6B0kqkkv2YcgTPa7mKFxAIsvwXAWIk2gqsl3sisPdRPW9eE
h/rpNnjvKNUu0f2abstLHgHDEJr1TZBNpHzCq2pX8D7P+T0z9zkoLQNVXxnyh2pBl3VUURnYFBpu
8huxzVjl0fv4S3ivwCOZ5+wA59lGyXBLAjYv40AccCW97r7wRQvWEaqscAmereJSMheZIfGL+Bjv
lnj1yUc1QSEVf+Ddf7mUK2mxh6kulAeiOeeaR2uWIVgfrafsOQ4YRe1fWID21aXiHRiowJRd0b2Y
Jjfi/rOn6L5fJ34RweUCYZvKh8yk3Ly0bq6OzR2ZQxZJFKH+K5VXdcn+/cg6cFT/oX2dq+VDtsPp
hFiR9yGe8QrXOe2lEgU/hukP8LP3f+Fs3i8AGODLIlmGzYt9JlreJG2ZsDKqKNCStepBGnJTJEsJ
bLi6R44ofPhlgnfMFnt+55mqhpAy6N4lJ+Aqxpdt09LsUFblqHy0E3lfyd2csTPc26Ob/ndsXEcB
hdzBP1QaI7cAdxAXQ3dwy3ryV3zbi+Z8Efd3M235yoLS6TC7jcIpBDB5c36J0oB8YjRdmtrbZNg3
XoHATp3Gy66unmcIAEpTLFPz3wVJoWZUkm2TCnTI0m0ArFGoMJnISc4vLNU5RoSAMaYnnjoazuR2
gBoP+M8RDe+a0f0YBQW/cnAuwjbcB0gKVHJKw+VN3I9LvwwrnYoDTf5KBUphyddGJRomv3antPO7
J59iEQZ9Vz0sZ2tLkPj/zeMFUXgB6c1QT7BmT4tuSf5PaYzYeS56lWmIdAnp5rjVGvkNeBlA9ONA
evZYXJbQB4d1uRdY2IT111zWpoK1xJIxzcsM3hwat07A6OLo1pXqygoaVM7eIlxqx9+XaIft/leY
NMqnk31USzVxWm5xqYq7VjN8lO81q9L6Czyhh7siPhwW520cGfSmMSfdOOilAabCWQH8sH/l/0Yx
iD8amy2rhymVfTtByWuFMODsTewYWrS0DRh9J4lj6NcmyUazMXXZqF6mpQOOvuVObGGh9itKVsiY
PkykEH6n2ENTTOSfoeFvT/KHJpFoZGGKxa/oa+sowWOyECx9JtWEuHy4NRnNjffewOTSD8bqQtQC
wu2iDCzuQcBkQX9sK93HGEtz515E13/KRyKBPFIYHm1+w6mV3OCmLA/Nb+7aTCzFqD6NJGTkbdxW
DbJ2SCosCakQlxs286lhoP1FvszGIv5S7B6WKUcQGAz7slLO1QcvhhhANgtD8h3XdjBefk6IlHzC
tq0TJ68OJLM0T8Z1Wv49ReGxKqCaM9izAKldSHnXKzGFDh21loodiJRRu6pgGHqGvysGon406yot
FA6mbXvaqOMyQETES7Tj2cEWK7pQ6wMebQbnqCCGNsXtVMNDB/7LFEeaulObt+Kzicu2MsHuV8Op
zn/1+Z3/SI6gZymzPVKfCy3nHCfdrl3KHgfaXKLxgxuKcSK7Fj5NKxAqQM6QcdIvBIhfLr7gcZGO
fdDUxmFPRBgyihHDC20AT1HS0PNN0gIlUw+GhAo/a+3gCBsqdPuEevFNnJKyU9mntJQDIAguY56t
Uz8I07Bcm4mU2X8Juy/h8cbV3rWX7irnMxUugT/kCHh3xCgKvMeA+BZwPqoXZfXyMDo2AVaimPTs
36cefFRzd3g8B1kQEmEC7iT8jdEt9xZD5f2pN8gLsL0yVXh8Mr3/W97LSTBLEqgJuma3IntGOwEw
Hi5ddMzWo0gwYiEGVuwuvuP9WdDDyGA8ZgDLXqPN9gCvzyP4UXj9qdFmpJR1ZNgjJg8xzupBVz3C
fsWIZ+5tPspct7bpOblmVbAia1YGXn2WY7I6MnRlGlWXGNZ0cCg/XywdJgPicqmLfDlsDVBSNM0n
OU/Ee+kCHBdoRDD8g+W16RIfzYQskyp3eQ360hhta8sPTJpk5DOhDqH5BDYSlmTUCroSIXspAJhf
2m5aC9L5u9iTreBuBfWhad56ePC4HClqJb1pcBSy6GsYUmU2YP9lzQasFmm0H+X2pnGQIfemCRbt
jJN2MSAYZW0Mlm7yjV3xcwtfygqqtZGBFlaVaHsZvpaRahttlzA+e4s5a19MGoaWzIrqY1Z0BE2x
CczzIu2nJ+ZX6/i1jj+SkH4pCcHoCZPJvNWCtvXI1eyvTaABy5yJHcF15JBEgRXA3AjFC67s7bZs
MDpdEUOUoQRJC4VIYXB6wdoIXwdwqWac1qLRN14HheniBcLhqBW3841krK+LvveR4ngtyTkSP/aX
/cVy2yaIcDfpfeueh46Umd2iPm7Yi2Q8d6UtpgYtfMhw5ooxgwZsJVboJzAxbi4l2KNMfEVdrxzl
80cZL8WHA1ynoQ1gWkYTKt4lkmzSVDkzPLAiJaE2oLwsZVMfHfEAMVQlZF3Kks5pH9I1yyBGu+7a
EYNd3KX2jv/bzQEHg80UfGC0vPkET/WKsVziWqps+Xq8M3LNWWDsv+WNHL6GvHE11bfPE/gDl7Bd
sa3IpRKBpbME8U0rc21s7xIMcSrEwvCjegnmqUSE3ifOG56rVqHZ2C3hJ+WIX4quUXcWKJVfpM6h
fwvQqBlCH27YCdGH+WakuJnVN5zzGLAoy31sCjsJ/AX6KL45BBlNT08AlBnkvQaRh1U/36NCVWd+
jaI2TgkMljTvFgI0K6gBFVNHwOByn3P3RMOzL2cxFFTGBGlBDG1bzHiEKFS1t17q90kaa4Nef7CK
O4ptv4/VO5IuvQR4oYf5lV1SDeuycJnUPAbD8ZjFNSWikQXHdQqPqd++dU65KgYGJ1DVVHZrU9NB
pfmtrjKeDFRo9Z3Ktg+XsQCMUzg/6qAtd6KrhQy2IkTu9/Pvv2MIwdO1004R1FN9bnaoUZCmFlQm
+j4+bXo5xiD9qK4kqRaKdc/bZIdxxcGE53H7yRZgKTSGLifSDmEagbkIylxmbpwzlUQ317pcEqCz
vXJH5dWHXtWBrB4SGxQ3McMktx1aDlJpOhi0OpyvNdo3T983swSiQiHLAdHFsUSl9f00/sqbWXPr
fsgxsBoOgNIJ/mDtAmDRJve6Z9LfxVFfu6ROmyT4DrWy4zmnXZZC6qPx/26QxT/M6odwR+UH2bZ6
voU2ckmbaZd4+PiZY8BIt7QfHkqotmXIFmmaRp4OmdYZdj9WNFWVYa5jVvf/j1AWBnOTMjf3MyRX
zdzjKP+XARWIBHjl/XSpxungwLB64f/i8O1ws8aHKgVl84GWwlel3KtDnWddCqgmVeWZoH3IZBls
B+gQW98iRqPAS4dpG8eSJZmrF3l6CPnnI2Ed893rDOn/Kp9hWw87LqhBcDhMOkB5YOv6faIyawKG
QTQKGPC0BZVIlROlCLIHas/40M4b6DkUrnYw3SaB80NWk0Pe4L2RqoTwWEtODRjMmIQoR7LLHyaH
hhxbxHzZa6HIhTBta6+UjaUY+8TX5lVZi0jiZedtspqpHngAv3WA7DfPyMIE94yNPYa3z34jYx3N
/MRVUWttuL1FfnasGQRKZcCBeR7jD/GCu0zqLB8MEissOQ6IGlQRnt7/DO/OWIl55iseHltnyOLX
K/NfPOA5Dr4stQSjcE9jxFuGRqqOWhPaBiUul1OqNx86Rflt1g2J2mr3bGgNecZ81nBXGCv9b3QC
G0HsbVKdflnsXqNjKN7YDzxwTMPshoDli3sCqK3P97dYMcQfIoRy11qtV6YTYl8nMdZrsDBMxN6w
z5ztfm9/5nh8hHCWibDrFz5kqJ1dJvGfP2rP5MmG+mzga016zWgBhov3meFcUNNsDlGZnp+h4bJk
mTk57cOTf4vs02L+OErHBQ3nT8FUr8k252mXyIzM9CVwMXCWPZZ1+gEitEzzGWmien3t05vUPKZc
sfDV9VrHNtK1ErSMdjUj5BGKIt5SgdRgTUjIHEjYne57NU5IQotySB/X/AsC9ECb2RwhtSYXpA42
oXGeo+0FnVD9fZAgh7rUckcJG3pjH+UfyEZJUIg/OFC+cEHE7FJU0YKOWtQEwh+eSKVRqD064waJ
Boi035OlPeeWHsqmFE9yZ9q7Q1TTR2Deg+M/jIoAyiiXzdn+K70iPWKVaVTi4zz2x8Va0+CzQcDF
bMDL8Bs2s6S9ddTXjneoMCjqhbTPyEf9ROkGzZZtkqv5ymFhkXJ3IDcsiKpNJ+cF8sMmZ12P8nIG
o7j6oOfencvcX29psDC8QecjutKbW++uKDE1wosRkT6cTSUjGb3Tb/6/QcILi8fDtrh8NSRK1vcK
pla2XCSaUP6r6A0ZrCWs0X5ZkiUANeddmOhf8sEAnaNa+qcMOPoQz63/FnM8GZ8Cmrlkwo9uBJyS
EM2R5ttglkXyIGZr+weTDWJ17zfPEZq5jKytNxG8O0NmC2M77PdDNz8f6HczktZ0kxfnUadM0dXf
9bEec2dkrs3Qvzw9CTlGC9BelhFFWpgpo7UxmIEO+yspzdUT9qVVMlRUrRym28auE9HdnSFWVEUN
TImrsg+SZdCdsAUrJTJIr1HAFV86Hc6GYlGCBOKNehhR89Nbq4n3zgkwWFqw4/cgjLw5eaGE8f6C
yHM/ghWEkCAjFfSL3D/7EF9re7cEGHn81hOnb1J1acBGUcwpxf5HeciiAOfjLXo+39GhRMfy2j1R
az5qLpb/udAYmTko+NmCLUZ/lZbAo7MiExpjdM+7SdmDGePa4hf46XRPqf0c6GkO2P7Dlbg51s1M
smrmjkpt2zdP7KrrNnbTi7Kqkk7As24mF1QQp5usWuqvRWMqI8FA7yRefTrgSFLP1yWkahaqKqga
5D9a7DukoEyDI58XlP5PoeaqKCAfdqXnfV1jGW3i4/p9OIZFaP3OuSl36VpfcOBRzWyWCq0Ph6mG
3pG3ftvwRWVWHqBKx/RtyutJi4znunWjYLUApgX1wYyO+vtOp/QNVP4aexihffpR0iT1LtTakOuy
ajVbw5HixeHAVMIkBxqoDZPFpGKnFgTIl1CsS341xJWIFOKFPqv+7N2rF2nzWRa0iQoOvG1D+ErC
CTAwrlsukBMikbKAC3cposTOYqkqoz1oXpzbmGa3GmmY2J6kSKpb9Q4mFHWt1GLHi4aZtKc9kJc3
DnK22Kpd+cf0iluMTQYXzL4yWRyczXauHkZiBFxrpFGZyHTZGRnuVy/6E0B/zjK93OoM6kOKE+y0
24vTVNaKc+m7sYkNlD/nWW974O/evzh2tK6wDgldHpPtWOaVo3N67ii8mqvg2gCQxvfBIlIucwIC
itOAbFzOHTELH2frB8ZpFN9jIZG2O8FTWSTEt7hF6qsS6nhYjgcHekBJoMtj4yAuiviX7AJLllHC
GdO6DV6M2muxCmnKk7isT9i/20pNAGa3+8VAu5xMtZFFIzEDKoBVJT9fPVwUbX8I7+uyEkB1k9i7
JCseJdZZLp9MYOh5seaODSgKr2WJySS262Fn8i5vFvZatF+LTDsJYQAYncyeyOCqhPDsMgUv1ccb
NjU6zytEJcA87aRr62haTE7nVBpURVKSeWTFKDMf/PpfvgpvNYL1eBp7Ra3gpzChN3ZSm8fC1EYh
fqTO/MJ+ziXG5K/5L9YN+88DpphdmnZpet/xcmV8joraU2EFM/IWD37SPSgz1BV2uEVgdhlda5WN
22S2MZv5tjr83nC+IjBt2LQl3Uz7kQcNywlRSJKvKUHzBXL1dB7JZ8bzC7Eb0uyNzr1PH9QDdi4h
O78hi8Aw60RggCkzdRJN0JtVdQNvmQb++QbytC0SgqWx3dP3UWiwd8fZasqkN3VZvdCyp6U7tdFz
XbevGg23zKLh7+1KjJCfQz8MooURqR0Ub1zi3jnysXKN6uI4rsdxSS+GIjks6s5g4hzibMUQGZ8f
pOpokCVm1G7vpQO1iY6FSiAlJaoIj0av1CWliSHfX6ueXJhwa9f9C794yBOpHDSAYh1nxAnmvLYx
E89ohK9d/ij41yS8vVKgL/0OMsytrjSHXh6SCbozXXE+ldhH8f3MNHgItcz8HrgDiIgQZCO3Djvd
9UsyzL5727BD3Y58L5mHwnPUUb7g8FnMmy0xzUMHjdwpB+WWec24ptm823kMbIkuZPUDEU7mOsj+
tXnjaAviLU+rFfHufVrbwD6Xmfl0kBWSwq0YePX+mxmamPjrVd4PsdKNx0EvjOazRcTwhxrXLC0b
a5pyvqPlCDqt22T5SoEfMhzbSuHfa1vymBkVTckTqcGcqp6i4794Yhn71TY0266Ht315KscZQG+L
iZJIycBy9aVsZRoa/HVJCvQ2WJIUg09GmQ7JKQ/XhiIXMVT4wLMSF8yMnqQeGzghClCAxk5GSANQ
SToC0S8Eh74tHXG6etpHacnEV+TsMIODoR90lGxHMCq/52K410MtkD85VBdoU5M19InuabVS6jiG
ta3Ef7SoYfx68uKymhgnaYvON5ZSL4X6v2aDUFMacP6M1V0NwzhA+EpeYiQw7R71apAL1KRDLYnJ
zjS772eT6Bu0RV0KCEnzYfVxgloKJrPBzFC7+j1AikmZQwn8q3Fyc0i+3NTQevIorUIw3rqen3Hr
UBZLHZgs4SknM7FhrCbSO2HkZHEmWkyzd8ZOyUV2cV01KZWxJJT2nxEXwSF7OCLpFiwDqNbtl2pb
n0eQIZQ31Ng8FErQPecA9o2n7huN3P5ymqRwcZJgb/umaehkIFotN+Y9AUTQFEWS/M1hUypEzxGA
YbiSmkDbx9cmkNHOou4JNrkLyqv8P6tPJcEOzJqPQeMcwgZfuIPqqS9Q5URzPiSjMqwSWVHlcKRl
FP2wHLvaFkPr/l7C+yFjNg7MUDTAlGNA+j45UYMeti1wqRpP2BEZIhjoXfAmt4T3dhRgczCJfqHV
Ll2fgiz1GwjfKfBRFCRAorqDtQzC2Hy+ARCZO09M+Nx7MNmxKU7E7yVA2ZselvMzRXN5yZoQLDtN
Pnx++SpXPvh/78dGB31JznSv+xj7GAWR8GQauqS9y2UsAgOPHRLraod8NPE8Pek0uB560v2q85H3
6x551Gd86D7rvJ5ZjSExT2jUaiAOQsD65s7s1dCSN59gAuTB2GEBL0jyfdOAznAYUFUZBg1MWnSc
Q0H/aZEymq/D2OYeNOxVSAhIXU+No6x+laOjt/5qd+NXp18Yiam4F/O6fyyFbN7eozNnbcKb8zyt
kDQrYoRMZnWaSqRziFDPROBons/azSCRpNn+TOV2jFPj3D3ihC/EgDrLajfkBVaDkEALTAhCamiF
GLXl8F+gkP5yURSDTlUsWDmelLQcdhLtW/IOD9vOK++KyCA9ZsnJ+PvbrOCUF17dIOCVP0sn0BVP
7F4WrE28rW+hFiIwfbP4963bePTLsQYxtbKkG5kCWAkJSzeu6TrQH++CZ+Lf+Wajz4/SxQmuqbbl
uil9UwFnpnE/sYbrndj+jTiTvWtgSA1TD7c5h4gzoRiNVnhlyxzGN5Nju44/hVDtlLZBYvEBFvo1
zsXFI+laWb+ZUXiPBPKjeG2fAUAvjmaWco+B5PaqzKH0A24FeoAHUmwK0Sk12X9nZPmmhR5Wd7kc
ZiLkz30/wFsS9P45Mq3jFfjyPMDty1NjIfeqRl4IQOEDIN8DzzUOG+aEerjpIBOzFflOf6VsMW3Y
OTrKupDM32vjgbBErlWm77GNEwWBo/paCLFno2tu9CgFW+3qP3fGRxZXR8YXZgf7ZnVFLFaFA3Uf
3ho+rv43hV3kPnMj+0dh40JrYR6rOoLQB0ZKX5+0YCt0laewDfH4AAoAHT7rPDbC0/c3N95CvZJ+
cN4K1HrvAabVibP/EwGU1qt9Cy6xLWVCHy2cqkFkYCK7LM8ftqSCWerdqYh1K5FVQv27uexhFtxc
HxIMOjJ/oMlHRwRhhxxNEUkmGipayfe2GosUyv/S/Hb7ybjZ9pUyT3AFSv6vf6zDZ2NLehCecChA
Lff4i9NYJBtBLCSoKQrSOFaL2jEXWkUZb4cc158wdZoq0xELt7Qk6yUkMLV9UWNcrOUjXdaodfFN
jixkb7Hs9RFAnAtu04dhrIFqNCdsLa3SW4jxgCD5QSpWK70QSdaBAFQBa70SMdkOMXDyZ9gkR5IM
wersRY/0S/v6gA/YtJCqlpzfS5nykAkI/VxurQnsi7KNrS3lT8XhG9TktU1/n2joerxlbiif01Pm
uBEudoFnSsipHIHlhShMlqKRtVWebfRcYec2zRZLg/xnjbBkWygMav72La9+yHDGLeg9aBBqcqK9
CqCsOnnPo/k2uDfG0CVfc6x+07/DwVE+ud2E7xeWTNiJAsWhIVdgUuFJInvQMB06Zj2TBMATpSH3
nnBf+etdvd4zxtZpVoGVIIMsCyhFRx27y4KfPtbZzZiZXR0QVxfyV+GKkEJz+qsdBzfd7WD99Wo3
E/R+VSanp+ie0+ZOO6/mdbYEYWEarWW83FOrMc3HHhbAoA06MdyJq1l3I8ren9/rN6Z9Jdi+3jBt
b20MM6bETT23BkfZfcRyedenp8GbADyg3DtfWWbCzzCEYRJ3dFiBJZMYaeBGCEmvMFlXAvMIezYs
bS/epwknTaJbKmDABdfenj6sVUp5DFJgjfGn73rvEN93dSptewaBrdNEguEg01SDNcN9HTdxAlbe
SNs6F+qhS36yWKKgl/u6aBtwjA+uvPxcLsrvuYGx1euNKZksxJsTri1PrjK9RzCghaDpRehMYAid
J/MrVZJIh/jWVhYKzP8z1/4O5ycehkZr4TfnsiEuqRxZJX/akOs8MgzZExp0ysSogsvMS3uXDg3m
7UosdFzq10eoBMladkzbdytKrOilChCMMQnsXUu4o0ALgIV5h43fidJLNdtv171GyOrvyGa4hCej
m7GWiuvkUs3v29wC+rl/QIago8+V3rKqx9heT13n/aR4UyB3wDGK//3f/fNsspilZD/HGGOZLZ3k
7zRrezwVVmpFF5eTehAFWYxCiTBc98rSjcs4Pz17o0I65WTRiVM53s4xV9pOPviB/ZJ0UqpoWNB+
UR1IOyWJm7c9G4SJQ1Tcr/0R4k2buJTeoCc90LWZ6ef29+NxIJ0LlWOvgYLKTKB0ErKIyJGiQiqq
TrKlCiuLzIA3QB5X7kqfp2/9df/jd3b31r5nOEJaRsPs8pyxA0YNMKdzjurC6ooQ4K8erx3jFJtQ
RqwJAILttJ7QZkQMU7pSKZ+Ip6+A059ZDgYow0n95FZUjMHmysyRobCkg+yG1NT+GT/KCGZz+wx6
f7xMj9vP71VDJRtdSBj+4SJ4TyKxebhMbQoKyGJD3Bri6KK37I6VpnW2jWJJWI/YhfZfybh4CJts
b4Mx/FpNo1VqaMntfUWxZr40rOoqNc7/88C38AspL9PRfyJ2SzgUvQBcPqx+cP3jsucspEbFXS9s
MbNSpof7C4ZHeTUKGtw1tgjNoaPhUKy/gw42THckPbGgUgJvZs+BkppS7MWYim383oyA4wDFOiar
FuBTmgFxzsTAXurIrTZ0Sz/eNU5TCGMhNXk0NMuTjvFLN55+2vbJHxdRZqIF+0IIkdve5p0kX3ys
7aafKSsLT2gyqr40Mvcb+2jJf4Lh5OZh8CrFGFfyizpfgmzakdgQfPvsW56RwOEhXH2RsMK2zn4K
7TGlmRvWEBOiVW3turLXtwtmOcMnV0fM9X0LBMe+JxOhY5SO9/1w09oLq+ryXBI3vqhPTuBF0Flh
SKDv+C+vlhi4lenFzI0wyyZbAMr5b70ozcm0ciImIUJ3iQIO7fEU/JBn2mfsCFcGnPqGo8qXK5XL
lby/MJMYvuv6mg8WjPDdeQHojPdUNILS0kEgg+sC1FEAn0lWx6rSxL9y4+fGR5vsEjmHTH7nnSZk
BdLsnW19B0NAytGrsf+RUF03cALmnd3/mpCcKS7XbTgS+R92vDr1y94EScO5gsxUZfQZtQvknaSW
39LDYusd84PbTFr/zbt0Z/ezz5IQskNv7Dj0uSQ2us6M3WgegCq1f6JaWXHHgXqIB9uGYPDZDyrz
pexSv9peHyOe6Fpdr93NychuBRQaaf3wR0nlIvZBQMyF43oYrkFA75AcWKkW6YxEo/vJno50py83
0beqgZ099aQNpTJ1MdaH7Mx27bIoO1bNxkxZ86ri5PEPHBFRGz6n8HybbDCiwqQFUer6zY6du0T1
6H5oSGuwrOXmUkpDz/IhnHC8W3PhC5u8tmH6DKW6ZsxFv1UwV1FE3NqndLRNbl7VQy5mvOpJhMt6
m89Azw25SagM0Y57+AB2qj2w6rBvK8TWsenlkwgpeRd47cyzSUZvYylllmgU9bOzXllPZJcXoIS1
8axQd0q7szh3GIlaf9Gshei5ZMEqysfiQvcDclrNH8phXL83gneZcrvLyCMLO3cg1HQnGhuDpuTM
nEFSlCGBsjcg6hOXN9jb5czPEPDfX8acOwp5Mmp+2B9N/mgbGA0ISmLcwPS2zdZas3ePYyROVKp6
hdxaqxacW3n+Znqkpoa/zUq9Q90sxSaNKQzSmyiEa1lec4vx4SEaug1UsCBOBcLepwIe7wE0r5Eb
ZybHfLxNvt63zlTVG62AXCQeGAmQLkfqHXpFMFLgXYs3f0HDHYImRrsw+d0fn72po2AlEfIZNfKn
1B9wU6Fx521sFy1b6+UfMEcilGaCaUBZ1Vi9nRZ+tFcSDwntxin0aaFtyLbpOrTAVByj+lg5s1Ru
NobFfL3V3q7+crK08Hx6Af2GggSDcBDZnd0v4ULgxBQVcD8GCKdDx5EV0uYww+Lpuff99SoCthel
COUjDzjiyh9I3svMPZmTrW7ogKXM5K+84/y1/nxKhNfiuCeOkqEoyPT2UNalasdLREwP2sKRs5/j
dFfSd2qtvDXbt4OF+2lQpqJ/p/QE2JBJdnFPxiDADd/Ym2aov7DIqbwU/X1CChjylNcV1ZuShPJk
Ilu8OjeiEseLr/Xk+Gd3uu+ukGYekMnorVvTW6tu12jSlTyBvZV2FmkIGNqYSXZm39QioPgBPya0
iIxO3EkNB7KVZUQEsOCeidxPzIRRim/ww7jq/c4oioIlGY+h2Z86x0cdri6DWVv2iVnf0jnGFhUM
wSH4Dx+3IsMBsSB9wGmUohhsWOwEuFxY7/8q7RHjMlPizkmudnq8OyvdTMLbr/F0d+I1jdtqPuoa
lUQBFqmeHkgM9zWgyeBvuQ1ngz3z6awe5zOWr5jQcOGDrY5aAOif4ed+OGe+5gmFeePp/EHx6eX0
XUtYQV7m58/H9u02UpNePjXjC7diX+CgR7YYlSnFbKus37McczVsxv04FuEJCIfrmFe97/SmwhR5
mgKJuaNOWCyC7RVpZskE2cJkJwR2zKoR/NGUw/mxrb+uXWYbrAhAL9IzzMAU662V+MfDYs0j2p+o
eeEPKkIYENA7WOnYRHBSQu5PkVclrK1YW+JagZDTVa6xHxGxASykDyJfMTnUPvVNv9661I+d1wEg
E8u4tcESEul5SHDX/u3TRv5eyvexznHtx0eJWO1JF//dX+8D/XIozPHPH+nFLSwkIu7lWrlIVP7f
jmm3vrns6L3bDNbsaDPRvYZraSlN6qS9K0EJSwB9OjUe6io5tJKvbNawMRw980FR/qVhLhai84ZI
wzyBPHPvRon8hVoZK3frqZvrgtNLw6TmJliXNbNPthqQ2F5qaDl3ifWwT65RcomSoPC+W0wax0Ct
///mY6v9uge+mLhiZHyyeBVnbiAryHeiIy0wIUmvrzWyNgWCeLFVeUI9ItF9MY0jhgAxRUPV/0/Q
FadKYsAvD8HttMXXgetv0ydpf+jrIyNXW5wO9OrMaPWT7J2wlBLDJli+VHM349y6PdK6tOP4DdOj
iLO8WSKGGaAAHTB3e0b04bJm1JipNMbB422YB8YLy2fdc8jlb7x2Bf0uH/k9Qz/xT2Jcjf6xAwvh
O8iELDOaAPXqrsLyjNaxJrUI0CXKKqRQWffx8HYm1VDPS5rttZE9TI+gjrg+ffl8gTW7LZhNUcVe
NL/U6RKXXj1l17Z+xUb4n0wRPgid4okhTZmQ4Ik3JdBvtXmxbveBgYA3djL27fqyY+FkjasAqUjL
DGfIFF0HxKIv5iPWrjna98N24t8MjniYkDrhDnVbeibwWWTyn1TOGaOp3RKXi7rE0uqbCeivnemR
cPkSfF/vNYyvIZTYLFimE1Ijp77i1BymUdRwsqCUjFSx7BXYHMrK0brJFdhOq7Fo19kCvB4U32u2
iaJFCMkTKxfzY4bvQLRebA0TkUNdM2P0qQl005vo0jWX+MgmJrj0Vst2+aM8f1Zw2CZjPAGgliID
WB/UBsSXfZhJJIfXwGr3ijKR5RRq+xVivgb9b5hx+7v4be9DWeCcqjyV31w7Set1FIwWSBrKZFvM
pbm96lRwyLatgyW0YDgK4ZJc65f/cvbcUxNtc133net7a8RihxBvZcgH3dXppNPliWrR+rTT8xKT
dm8fU7cRUIGrRgEXzHENqgB5ATBkjE2g8b1Tm8pBZx3La9qLHEhGdjcBIjZGupROhSs1swoxCKSW
qciA3uxFaGRDX9LJgnYn/zAyCxd5IH6ky77zMqf3UFazCfHhaJLz+655IPcKIOGSxx9GYDhY/u4S
I9Z0nLB680MVf8YwQzln5wi306UrUmzXS4QH0MbChZUw3bHgGjNv+EyCaICXnjDvG22xtUAaa1bw
1kRLfPjsLUwM2wy92Y3jXJBskLhDR1GJibmS7IjMgcto70qJxP9Iu8kbxbSy9np48WD9oqtFYgXi
o+fZDwR6WIgSMUppSjPqg1Ha7trvGUb8pPGL79pOCLpryDiHeqdBrtgEaNnpCdNE8sR+6qyXbHkz
EDLzZE6tVM2aLjG8a7pDkfWVRjI67Isinl8lre00KLbG0orjLDLbftcttKqvk7HlMmfBKfd9xaYp
x40WFQ8GtxVW6HRsoD3vAYOcl3bdt7uFNICwcMtLs797la+ZlbtzPYbATHXD9pchU6L6GWsZYFWO
b/5isz5GgpDNW3qekIYcVLqHN+3Zsli/2HURJU0Dud5jz7hSuLKGJ0dd+MT9PJjSan9lZfKNDfsc
OTjdrdvOUviIGLqbCAp/hFxXMSO0SYwIS2eNTeLCw2Vvup0/W51ku8rcYWiur0AbBdawLPBHvw9x
yI2t5dLl3abuMtFDnNBv/4AETmtIlMKTk5NKXXZki9PQI5ZA3y23HTdX1IKBg0OvssmUR79aRfhf
U2PG+ObGyFFEn9lNQs7DM6v0i1ycFo5NGPMcBIhbjTw0fedfwoN2AJi1SBeOIo5fZmKObU/kStia
lW/kYmglKkZpLfhetGYBbJ786oBlLORwjB1PEg30mutUOpszzeh6bYfsBvhcFo9M8MTwsampySFh
jpgf6u17VCjfp010S4GzeM3d5o2GuY/XnJKWabTmGhj3mcnwIcW0Zcr+y504fsdDp+acDYe7pTvf
LoCH6vX0gtBGCODPKJKHN82uvhfvSi8uRHZ82pA8rye3SSwJM1BQlJNxegrNiWw6xs2Z9K/aj32Q
Njw9AMY6cNp7SlU4jj1ESCi9xOgFHfgZwSJLAVrjYwvxkTXhOdnJzjCN79qbk4CAZD0h174pCNdI
8uBGbHe1k7jehwOunirqiBYcEXuaAJVEDt04zCeHlxtPWXdGx4jKJcxzXuoJmBd9lE8tIHYXO+wz
pfwiTyQl2GOQz4AwbEdkpVpjDoBGGsNE7ElrrV4Ymr/ZiFMoWhe+rbQRUwVF7h733GiwknlqWSiN
sgkoF2oexfemij6ocGJFsHYK2M85nC1mf6TuTQMKiaEC7i1l8OHP0HhwjB5uS+DWo6IoSrzOVvDQ
jPyJrGIQoBCAivD2na9r4vgZMFbo80n2i5CA2cWlCZtk1QZhD/3j4zSCRMuTKz+lWMqL5UWi72qv
bMbxtYxrvqjLjZOAkU6jiNaEW2id6EavrQPfi5nWuPkWNyvYbpkqKg6tUAg+S5FzlY9hwnRs83Qa
DtvAkhiZkOvG/ozqtqDtdUYjV/uVSJxN+Z2ofDCESd61rDAvE4/BUY1vtVSUGou3IUkr85n+RvQ0
Zfcsa5FzKnJzfgrjyxDpcupaxV/1vCYM1OsKUwrzjTG5pYVfkEFPOKdYVtipX0K8+vpfZqbIa2ql
Gmj0KE4r5UCjjQOC6mITzUOeSBseJu75ZzDGKsB4O6UuPsYxw5XzmCDk32RNPU1XhCm3YXbtVMdh
krtmVxa5P5CPplKGfHbtq5UUU1NNbXtnBJGq1J2/to4lKmQnwOPYvw+j6OZw1E9xQBzmI4XTQhD4
jcPFf7tDoB+bRhcKnuI8R+r7wG8XMqX4Cbl9lgwZ7QKKCVuh2+5+D94USPeOE0PAMXeygNwZT1C+
JT07LEg1Aa1fvH9s2IX55cyWDw+oQ+/76X1kezAP8v/KW6oJ0Yrbd2zLX0r3PWRi9bgpvBHcI3+w
Yx/NjUZ0W1TrBI66V9MJORecjOvEw4vNumj+VDz6PpND7z4v9fvCWYPEth6RmVYxTrl5UoAGQv0B
WbPTkOKNKr6t9uCX01tNFG2/q/zhJi6P0qWioYGHqFDQAY5V+Tt3kdQs8qla4+5tVH500otTP4WO
bb70ucMxTqlqUj8J8iurpb21F8Fy5BWVLft2XTkTpGiwb+0CsNH1HAiftV4CaoutFHyAIw6m/x5q
EVPIW1y81OlRa2Rlmz0B5pzAxsWcIswTLlk1odUeE1pj/RWMTbvF9X6/UmyZCDJMLYzFyKjwYvGK
64lZVcpqSfhJLA8YNaKCn8gx1aqowFsnUjmqTjSm9OsQe2S6UWQxQk6Ukx5wt/7zIdRtt1busZf1
8vnYdGuESs7gANVyUFuhLBLJfCATeGCZ/5D96uANhUgkQ/xlheVOBdxXHlxiSKVgfna+nuls2qx8
35TznmDFHyiSBwA0uGh38fhm2rnj3CT2ocz0CrLdOrprOh/NciA0kdtOc1MnHuYitVtLamcpnuqQ
bJ9OUD+6qrP7r6QJjatbiLkbkw/6BB2EPMSPbWVDfpJCDLiKre1a8hif4qjaRZi6t7bkHeuPPer9
PwmkNoJUrwHkIyRSOmiihShOTJB3kcN0Sz05HNMxUSrSadneX+SLrUH6DmCBQ8eCh5dVKAB8Ty46
LU1AEYGjCfsVBPupUjHne6DLhkejIRYmthIJUX4A4DPDtkPc1o2T4G5Ay3+81t/w/zCQBqefsYKM
JlebqeU7ec7yPUxo4OW03MRw6+AIAkmY0YUgqGdjTSib3dTMLrcA/OfFnQIqMxwLG6HfaxR3Eer4
RNPUf5hQNUGC/AWk5gsNQXX1C8WuAUimcELtTVt3yLcV2MvkubFJKv79ugbawye794vU1/ZC6Ngc
/3ia+Ci5smQvJiWxVuVlI2PecACdXozch6KtmMFn3JJYxYMd6xpuEkkfCc1fim3pxZj1t7kmymY2
GQfRwLlsA+DEGQvsm2wfrUcQ7HUWbZmauZ/OyMob3oQaO5jWowpwiOHoH7qEs0TztoAz2S5Hb4eK
M1pUIpBvVb5LLVcqNTp+sBw45K8HFtHYjxR+ZIZt7Z0GTxBWrLEZrnufIf/FJTpaGS1HRhKxM6pz
n+xqB2W8CI0q6IOkuD0mJ/qO3mcXI2NYE40Apced5UY3CTVLK9IjghA7SGlAzSkdZIlZ6edn3S78
ebQWtZbYdcGGBP6sskpt3oqlDOqMQK9+OucDDFDHPcMKSV9xxZmAS1At/Ao84cvD/7TumweC5yLU
NzD+z94hjN3aA6XUYIRZbmqwIXOC4QcunkAUw8YqEKeQvEE7Yit77jY4a4TpsPuQeUZQ/OPJYhkf
BcfauNP3lAEuki0zz5ulhCchrbZPIDtyze7hUxUCxFwcRYwPfCbEgvNWWVjX/fprtrsEXsEcjxIj
WsGJNCqJtK1p7Xc3kFPusslsO2yZjYpb6jeFNyE9RA6z1rcB/YxpBxSSMhdlKwgN1i6Famn1p+nA
27ygUZ/DN9DTkkBepkNi0d/PoxJy7rA7ZdOqsG+PZRedTcPPcNrY4mWEdDmnYloq3kGpohqqxA7L
gAZibsM7yrCY9CSCFbs2Lt7X5qlKsPGj9i2/f26GIPihaaGSCnms8tXtsCzaOyghC1At0hkaBCa3
N0ZP+7DimNZGVUzNwb3FqCEYE2+d8ubIgd0KYDhehjEq8uLkz4aucAiPu0zX6LZV95oOtLrnVGtw
OH/8+CAjhjM6+UD+FMoXkWi7GbAuNhob/KsLHwzLJy8f9TJxusaVsGugU3Apr26qK/UadPQiFg9Z
bWPvvgRM6mUySWH0TLXQmGikIt06Nkuq8OXMOs2js2IIxN9ODr+/RVknT6Ig5yNQ8QJNw/tD25T3
+W44uA+5LJHButDXiKLffSDBgJY5LwM3nNo8qmTBV7i/1ZF0vjONOqdu5IUJLLcql4OTGI15jp5w
3+mKhMNshVkFQahVlZjhreMN/QtjR1shANLAiGheUea8ZHUwlVxQ9mKJBTnwND3sNY7EGbwJDIBZ
i6X6DHB3qJmVQ3V7viuLmwnIdKa9p69PX6oRI2eyWqajtZK1CXzjbGQ6mcMPfKMat2qldmQYeWFo
TpgnRSJ0A/QWaM2d0DbjCfJD/IxUCn9LeewoCjqukHa12At4sxf3xw1+xkalucM33T5iG0xiv6Kv
D4vcru+mWnq5PmuXldEHg8VhxVWUxe9/keO1PTB1f9qUGDg0NkhLkNCuDSSW4AXslztIoQeb7yp+
XnLLsLo/ViMzgibCFiIQ6gKHX/a4yHZ1QgykylJXUjrCuD+rX9EvWXclVLU4A24kFOqk12Y4eVhq
oiJMn4UnOl0aNPHHqY4aeD+3s8kcOz3MWuhXTjY/cGEa1bXKcdByzHSCq8PKnbMwyJC51OT7Ffc6
1urmH1ubb9Z9cr8x2/ju0AHEQwgloIQ+MdddVjGKMiTfrR29S7jsKUCIHQp1t05jo582P3hhdPIY
6OyZDtH1Jd9wcMyP8ABT11XQbOdgckbJh61ptdyEiZQ0er4iPb6xaPRi/mLuZGwhuyYaEEm8lZfE
/q2/H1JO0wGz6uh8REUwE4np4u9B/wCpvXzWc4ynOtA1YxQefXLj4pjk4X8JDMH+wrClocFmXLAZ
QWuw9nobkO25sqg1oL8dqLfqkgx9d3NcQb7gurcu1sUxUZcF3g+jNL8Ar0hSzxx17DnIOyNRVLVe
afP30bhlCTr8mCLoNMIAfp7+hptKN0vHoH6j1Mf5h7k7F7PKjpMIKw3XxMfZj7rYxkVQfeLNqU57
KnKaCZucpYt+ngx7zZ2W5A+lIbajuc3W6sdEEsoXpRGA6hefMMkPeA3NlzemWOiLIAelJyFSjvlr
fVZl5jKZE7i1ib8tkegoIlD62zTAYCkbhwGoZWD0PXjmvUoOSALaY87IPVQZWHUExHbvHGz58MdY
nnla4WQ92CwmBfsd9UD6eKKk6w/6xC/eeqJfbbArkwiC4AxqY/fCW76Anr8BTAlfNEgftj62xYQY
BDUicNmvCUAEVA6DWzuEOMTZ9xpNciOhqwwMXLxaTKP4Jyyf8Sf9Vw/q1S2TekwohxLy/mvaX1hT
Q7+sllvLN2EElmTHNMim3VuAjmsX1Of1HlXsryuRLRGXx5yAKCo0TSfgkWrndMgvxbxsmuYLT7tr
ed8AP8qzGQOG8pveSlPdlyrcsQIVj8PKu/1CdcdI9Cv6HXqQ5qJetc5CwAMH1qey807VAquICrl+
hzv3X0QENz8TSoE0i5Hb4wIhtrZ8bN1X41ZY0laoUEWjjtbOF/01Bxpap+L4M7Wor067Hb6y+klH
pJ2rCFEAbfsEFvv3nbFTGAtxCqrbHRGjyWknpwYyuaOGS5zM3YMs4udqY8lUhsrnYPBp2mhtI3qi
apBnOW5Refr8CAU/AkBTn2zjVJ1hPuAmR+ZmB+9jPY9XSFwO21RURLGacR35UHHwrDr5udb9h/sM
vM65PD8J+LQcsJ+1U2JS4dJRIdQcquPCFx7noWU5tND98XWODNOfhwI56f65965l+JpjTCpqe8bE
BVwXoahMBQoQQ/yhxCQkD7aTikZm3gvysytR/mJSDnid8Gbn3iZ1PmFPSaPUdGG2Bl3NydvVxUM1
z5VRpzJ15+2L8xEcmM6CKOSJFrrd8OT8cMJDmNuZx2VnCKDaDSnh/vTjpffT/JlanniNkbz4soDG
IS+Pt33wNaimVsqP335zeU/SL7ZueQhtq7P14qTwYA0hdapRwrVFi84Nt48Ap0VkMGWC5ktcCmQ3
PKPmZ12V0yO8dQFRjpqVdZDGm5AQhkm7uhP30nmik7PAu7YtMHBltkyzxJF7r1ORi55hcUUvgzBZ
vEbT9pzp3tbhog+qnRi6AvouEC/mVTacc3Yzuf7D1xJ4CM0ImKwil6bgvxld61ovUb1bnB6dymgp
loWbO6rCQP837UkZmJJjEy7PffMlvp7etQuo0DpLEojMJUXCqe3190gL7e4UCSfQcemUImWbSl5w
zbU6pjJZ0EOyNWL1zdCNiROI2RtgPlFEPogUhij1cjoWHs//mfG5l/OakO7krKBR6Hhl4IutvYqp
2qzM+XTylpi3ziqPTeVQ+KOLb7R6wafq2xJa2oIg0zIM003grHStX37HmI1+cW3YUoVTPoF1dCXD
cLUIlj2I+T71KrUjgS4pa2C2CQlAuHedEqhedosG/y/gzzmoleCgTF+aSyR0tAk0lTwqUD6Z5Knc
9jK6/kgMctnBqINCFjiAAI2Dtd5A631AS12ZbrSS6KiBaxqZmQ5MxdjwXXrHUQkbuCyvL5cKlEiK
rt9P3Re4TnCnD9vuHCTJKhBaoHOc+/+PWnkR1qzaBRvHt5G36MZz3ttVWzWvdE/y08B8mp7nD0QO
LJyvb5zcB81rehEm3Flk44eKazCrbmb9vyMF9qK+GHyAKHZZZGajRgm3xiH1Fra7lSEWdpTQZYIV
P7wHSWEoIt/xaCER1InTNaLIE47z0KFjD2Gl608wPgR2pG2XT2A4EdzDr9qUxil1mZvTwEPTEPhG
wHhhjazTJO9rZ92mQ/O3PqD3TZojXNjcwUV55IodIXulfsEi8WPHe0rHShiDBruVoDdDQgUkTYsj
Z5TxznZ9So1PN7HQwDtAn/hpyHtwvZiVrXtcjYZe/VEBGSzk+avxRS9sHo7TGZGO4yRW+yN+FhI6
QeLqVjYqIUn/8PTajWDyrCd5Y6QXp1qoqEVnYxosJpXSTHCEOgvTliEsXhyLjHFPW/3+q8ATo/rn
3YSUzPQyaqi7RVa8e1yp1lp+ueSfmBeqPMyK0HgLz+0zrFITO/jS565JwwU56yv7FpFfefvvsy4d
BYBGmjXzPVxejxxz1pdtlmihbIRUDOu/EFfJeB/Cit3qdfmRccq3V6gd/ZHWG05bkyerVb0FDyJS
Lmi0gxZV9JnJpLjrML6bSs67sSIzZznk/cmxLFhvqBwfOcsdbnU07Vxxgr4b4R9oKnvvhmWuHXzh
Ib38zD6sPMckrEWc7mCcTk550au81sez6gGOp/TNW3fU1u2gs0J80fO8GzB2gxQ3O7BeKwrZxq4x
Nd7LsmyWFQytjbzFyTbw7CPLprcI/acQHIJpnKpMdXxP6qNWZPy3af3H7VkuVtWD+5Lzcd1RT8gx
O45uyt9Cy8QoZNatVmNy+aDJj3KNhBCUt5cuOWTvc5c9rSzArhUcdHGmip9hvyIn2fbGzFtMObQF
0YvKqaxYrdqeb487AhafFvingppBJ5r9DFYR2msXAyWRTgZnktRdH4497YOYW5yMiRWJTifyC932
TdOaISu1c+iGVqB9FzbkiwnJUbyVz5K37nFVNUoaIphUMEPGCwgLGXjpLQpZV194yIzxmSo5Loc1
cbA/XjZhn3MMdC1DaFVLsqzq6FFNPFjWqneBfPfahzvDzWmZNqVMLDzfPfeIgHf96JgpL8cGf6j7
YXBB8I96vg/YQCCn0OZYqq2mMDL4PZejAsIbk/L6fDamlL6pSHalnzahPiD86VT7BYPq0PffcBSP
WtV9y4OtPCv798+yfl+G/clXR0vVG4ViZdALjIN1jm3xPM/dIcyyG+QfI9h1Y3mr3ts4XclUAf6A
P2NC6ixW26iRMyCj+EpGrv19sBukOwD+wQixe1DNlnWfNowVO8RPKMyvsiIGZNfq2laYpE+dOXbx
xRtx9+JnGGpf1nfmnvgBt5V+L2VvmxzaQ3UaNGwm9i7iqT1GiorG5PgeO3J5b79a6OH8+qbThIsU
JSvnDSEuDqu7/H4wGpc2QFWoKqPU9mIQGxKKK3xT1DfcMB2yudeQKGlQdxwa4Mw4hU4EuEQaBsl7
UsH1Qm+yb5EgnId0Ky9rq4Bv7ubt+17303Qq2tDgnhCUUUsHvg6qAV8tWsHXBWKmqLUrF9y3d6c6
fE4LHnRmZ+4pBR1TVswF4MhTE1RiSaMcHXSL4vC58qYlMZhQxIv1dR/iocunT/ONiXA5Hr7H/pIA
eej6TIYLfX5YjdvVogz2z5Wgk00LFqKCeQwuVEJ+TrcBGCKxvA7dUEBhnShhl41wx3MTCZRl4ken
q6Gec+5ZuNDTo1Wi+lWzIu6KsV4oUvBSI8lEHWK/mhkF1pEg03hsOKbIdTPc+Y7dFD3VdMeB5JvQ
stfpwZWxgJnlNFbV1jt/oaOgrBgvauhzawVpREYdTsMlKkfbtbTOpaSmJsTtr+5qEk2wxJQk/TeU
n7Q8sZnXP1TOpwoCR0K6nkpX2xZC1TkgQBNJu2iiQg4qtn2qQB9sQ1220rhQ0XPHDF0XLZXsbvDP
zj9nLTjQsMeLLM5HHZE4Iivb6PMmlJg1wUdzCrO4Pzx8pRztzY8ZAZi3FAd9QuBAJfg3goDmoq1P
xq0Y+ajzHBgPWs6uYlRFQ4dZmpls4wXOKTgcY99Q3In8B2LqwU0V7S7Tl/I3eLvuK+bcqfYceI9j
spBHTQWSPu/Rj6gqxLilFAKoN1ONywNq4ATXP6Bk9YoFKRcx+Env/dA/E1bHztR6lM8u+EzCFPZh
kMJCnlkY/G3VZUSThHtDRvWV3bmSAOKhZMJjbnSMyQZcb5anwVRKrDo98ecUzI1vYTPA9RO/Txfu
YA90DPb5ja3fp0mTRdEoU5c6c3eF4WlnNGznTSRywPTpMw+IGbrWNDU3ms2fH4rG1LRTEBS22+Vs
ALny0nFGyGxyjxi0XS4bj6HTqraNRxO360+8wEAA1x3SqAajUpTIkzbNbFktyDsYnFi/h/H3hR2l
THrptqZoDzzy3puGVs0bwkiew+7YeSQK1CJfd9rnBYV+OvGjoX/hZRRevCeI2GLJZPMu0hlCuvh8
aWHSNdS9ZkdTPISWpcy3fxhSTiS4JJoTSUh8Awnl4twcU2oQmX8PRNS6sa4pNCgSUOO/46hJAYXg
rDG9xAPCZsZVvBHSuMDpNML7yMGoBHVlSg9M2+vuApZCP/UD66Ufdavk5rt+f6ACIW86uuqvf0f9
VADi8eB5adN5r0poa/UeynxqkNwZc4JwllNkT8A+VqEc3y/pvWFGseu7WlLSVpv+8ZwY0yqAywmR
FjBni6ijPgcmmdK4S1GnD7D9jciDBsSBtL93MseOnqffYnyDcOIa9K+yT1n1bjDooF1uS+6d0MSe
dUq9uXP6xI3voGggdo5UZi6BznQG3/uM15dIIMjprBro2nlj7Siq3yYfbZoxvpMvJaH6YoGR8kEI
RoaXC+v16k2jwki8VADkGrk/9jQ2HpTRAztmEfEeZ9hn2NJGvzUL85CsZk3vxVosNM4pZjr8RLbM
7gyyJg/Nd9a3VDEB6MM30yeQAVFxWHmK22ynq/OujqOGiFe66B4mSETZth9X0AHVb0J7QH8a9bYP
yYnLHBWbomUHnyQNSvuesWytTHoklPlkGSXtzsR63U1jnWaOyYa3+JZQi/7J1p4Abmq9fApOMD0R
w44+3xIDHV+1vNNpziG+J0x143NEQm3jvK/FF82w665kotIsZrqGiZ609InZRmsUFz5pH6aOBHXO
XSMjPff9OpQO2HJDdU5jpRK00262+noudgP93pA0pGuQdgELKPKB1tEuTrdq3FwUAuZ46c9QbSvl
epM7FUzbCWA7m5xFFn6DhDxF9twqAJPcI0L9n5xxko2zbNtDGsryz3q3GdW1DU3SP7zdL4Oq8Zn4
4R0JL9rCQng2CdIXr9leMn5f0qNkiDTZo89sgiobaoyNgDOE/0BqzZE1eoOKiRZdwcqhLLye6p/v
hdHdcx0+cYe7joSpaDM81Nc3xkdab/+D1rN38sJ4MO6eKhM+SINwvYhNTzNMfN/UftIFyyOI6GiR
7n6YuPhevthGzUc2qQHI4ZSy8Ym17adfjpp1QXLs0iNgt2DqoUvIN7o3YgQ3F2QiXWrGNB9UlWlS
HjfqzYV9smlrLaGIQo4xn0+z2dFgSuZEfJMJfnpBLHdHtQb6HCug1D/kXVNtGI42Adb55lZoK1Iu
Wfu/btMQnAJtRDu6xgpzkken8FHL1VeAio2MSiUXBggWWwd/MrY/LV6PNYwz1292qWuGCswpMFFX
BcXLF8g+Ngwz1/VbG07rG7A04dAdjaD6sIuhvqXtpZmziqgo4Y58YjghQttPSfkpCH6vJPiWNrcH
6YQ8+sLU3Da5Tvgy2BCXBd6eTyJhCtJnuAScxd1FJX7H4fTr/MkRd+katVMFAax8ppnIzOmcCgGE
UcpvKjF/bncTC/immzdg34tHddUOShjed0zdKH3ekFYdjyebdU5zhk9D9S/qrHqUfUh5iL7P7l4v
0xdh1oazbknu3+NySGrAoiYImI5sH++z4qyhT54DO8dtSkflURxreR+K1H5lGxCUj7xYQKLnORCw
kPIPGJYTSsiW607LRYx3vwOHRPPmFMjTI+Vt4w34cZzniwsxtbOlSAD4vsuJKTzN9r/USw8MvstX
00l2BGL2b0awbvvQugLX8xDWkR7VcK3grVmJikNU/qWX2yTu7NCDr+Z4bgKHsBOhAI3+HdKSYFCX
YkhHjruM4etv/t3toOYz/ZqG4le6/rXbbKbGgr0bMjITo2MlA7wTiblo2BqsJjXM1wpvIARW9Pud
b18WmoCwHJO2YPb1miNi3tNYwT5qAG/Vo+zjr305iQFwexqQqJHyNb0mSzETqjCjGqLwzCUP7tSz
1IrKhxrtJirJJX/OOhYEtkp4yGlnbA+gi5sFHsUlLkD+J6A17CbkdtCFZ1ULslancyguaC193Dtk
D/EtdcruWHKk9AJuKdmUR8XP9LMTHuwoKYSUQSeSXeet8cdvP5XWyDw/2Xnvi3q1Y+Cf3M+6ZSEs
jLhbPcevTjFJW6iEMBiyf7u8Cl4t2VdKVj9lXSqussd3msv1x6gwo+pA5PB7pKSORg6rUtSCwwTL
VF+xs3bQ+ivSNC/f42svyd0UPLhZ9vZU25KdZLMP/fhkSeKSbS4ylDoFkT/cOJDBGIYRmJTSFNYe
AFPGLSrA1oFPoyA4UfEiump+42tu6W6zExPk0kZp0sqGHbemAf6Osl1yKWOceyMx4WROeCIxTi2a
KRE/QKzGvZi6t3QPQS30yW312aNRWrRosqsFNJs5dmqh33qemI+Z0LPN/2msKbAbHkQuKIEvW8Nl
iy3piGK+EafoZRKxOu/zJUZLx+GNYSFXuayg6ptYKqyD64rCeUyTUNKpPLXAlYHKT9J2QstgxaqX
FAsH6YWbDzpvCJtdf5VYRLq2RvmOGuvLaWKZyncF3L3aKYN1egtO52YSlS0dAUMX0UfCy9hCavVW
hryU5pi31LhVCIg8V96C1GDsP8ot0DNNa+2ITyocw+za9pokfx3ChZ4wTuVNa69Fl9ARV2fOdYej
yixY6eq9PU/bTAEPgypRQCZuIGs1zohy+iEEkt1w63hQsupXVpSt2mTLIXWGaAY2hkEPOtwVUJZr
rhgwzYRUaXlaQPDcEJ94WmVio68flpgMcJ3u+Rg7I49ahe/COwkT8zgwZJj3soqOL77HSBfg9DKj
fzv1nqS6SxnY3mWVWdh3U424PpXMce5WtZ1BfToKhurfI+0XjqK+G7vbsHAiDaRxHKej86UsxpUn
sLEAEX2zjeQKLueVB57g4GaC7TFd/fbW3AI85Fst1FbupAq08vRavrces9f+4LzftKzKvnDb0eVx
z1o+1j7WxxbxmYFNnYwh1J1VE/Y1+7PF/qNd8JtF2KrTZPl7qR8MarGiIT9oFUbHJYjb5h65OKu9
WSJo2T0qFbxw4xnLmlPnSoJMEfMbcIjiN77fFOv3IqhXEmolE6fbbxs3qS9yOPLGEy3sVvHB+dRY
HLs4qlbd01WVXT8fFctk3afPB24ltD916o1zxmIVsG5HxLW6pGjiP4qmWqKFaF8h6HVePilg0vjz
Xk2QIgABmdmxmPXyjHvftE96Fz+iGhHhZYtwKY3zWjWoY8PW8fOGT62uFiJssBbAfeQD0iZfCtGG
grX2UP9foCarobjE2kC96P9QaN7ncaGnX0RN2zaoyhifr4BSfukqBDDRkRZPO/fzKscrQwC67dTH
0mWEluG9bW73pgNi4RjbHBHYAfZvmn3zu6oHqcaK6dQDvcUkruI91Zxt5HIL+L7NhhcpSDBpfbwW
Z3np4s/SYociY9vvsrGMwcbiB/TYoN4QDMH+pclXAIWUj2DvvrGNpo+VadzQGfeICsy1F4cMMlGg
3y/6Lt7t2w1JfT6J+N14Wq2TQzZWo6DlptoPNrV7RhwxKzclXcDQNMn5/dMym8j7BnmfaS70wEkw
1W56dP1q/idTrk12sWpagwRzKH8S7TxMNsBLNtN4vXPzLSNmCS3wb88qZDVTIiPQ7m8dASCkchP3
7rkZgsyjV7sMCziU3j1WvqvcOubMNPgg4Ma0BFzTPodUHk3KhmJ194sWFrsXMSqYrZDuctkkowUE
XOismJEbW9f0dvqniw7Q9GHlki3TJUxXAzqcaOxH6agcykbSUzrBsTMc/AoJhH7WXynO+5dEv6i/
NlJnVqeK+drzaGloxX06mSciaPcYauYZhT7s7inkr3KfNmjGRqqcQU/VYTtOHkiQG66GA5CmhBpJ
PaUChwu0EOO8sraMHvLQpPR1vImubJaMViMKEUKY6qqKthBJbaMjaWpbzF9PvuLZVY+1U2hU93Qr
zCLFh0XPbsdiPwrE46urTCVpdGDpT25p8iyA2XTT5AJlF+vdQUlQKzMd6fzUm69246jOAhnnK86p
G7jKh+epm1gnMVk9aBrVL2dwwHLTZpnK0EWPy6aKPQQ5v21S9izidTn8tdHw5JtDfENnW0fRzszc
QeDcg5nlYZvVpWdzJzMV9jA/pMHq6G2pZz7bsCWUFE2zoRoKukJC6pUtNLt5QS5dImuzz77OB1jO
BAvaUZE1iS+5gfVdS+E1v10Xa89vUS5ETzQPUsvt9TvCcXo9jsGtwHBzeaLRpOlQfdp0TW0THitk
muB/hem/8RzftfA8ZdYFxOfg3X4ZwCAJjuSfGWkrl74YMl+TynjBIxYETywLjrcjcQjpKPXD09e1
Fol1qUjb9v7YJuOTeG21HoHmDCq8eg3387ah+h5E7Ebhti7lh8UB0w0fXXutAoqk6Y9wOB7iD7Yr
115ZGVICmt0+r1y3uewfnSQH7ZChnv8uTBV2lr+KphpaMs0huXVNKqcUaAupKh8dmjnkVfjZb1+G
fT6TTQellt3VaVhjBcO58mzlzhH6ZJ1oLJ8LfNpLDSaOHEeBkcW4wDKp+pVw7d7XC1yUW/vlUdsz
VldMO5i+Dryzbkc54aWFAPiJvF4wFTpZ5XNd+1FQ6bxf+bn3F6gzE7cb9ULgnJsq4vsurRjG7PN9
PJNIAVtq0Li3Qr/nmqDd4rv7B43ur4g6gNboBx2HpP2QyhpFb54QnLJPkEeB3aAuLd/V3wicluf0
0/1z0ukZT0J0yP0w06F0/+KOcjFWcG8UyaxIfljargZ/iFfoehJlufJwLLeIwSf7PFqjpP0V69Yw
bPGlWqd35GeW0QDUPsujL11LuBBc70xNrDUpe0KswNHcwejJ35CqGo8VTlP81xr10jSbySbLVZ7W
Xc8TYcQJ6cCNfo9QWwiIGTOEcPOxkhLz2w9gWotyD9RfQIK7Db64/fdlThHOMr/iB52fEyTdjFWf
w3HUDFFXxJmgc+qpyqw+lWr+Itg0mSe6bqASzmea7ieTeIyfdlUjGJip5t0oPnHZoqvwSfTwnNms
0yGezpYpShV2JJxw8J3Cb3ZqcIcMF6ssEA9VSFrhLksnWvcH8g6s95pfdqvPp0/nE/XBlYwE0Eze
ujHOSHtTOPMfFXYg4b6neWq8N/EyAXavCJNuXxvSLr5YDNizMIsNDVnKZdUeuC2GD6aVbkNM5lsL
KVlAE+fDntlKbYtdIlFN/s3BxkvdOapuURlFFYg7DIRW2z5VHMUejYUGRMmuwCvR5iIXY7og1ENO
usu/x6L1OpSLcs9bqSDyBletbHmESgiGJ2hI4M3b06ZEbxB5Yx+uh5ZKYDIJwO6I/7oYpKZ6XQuw
bWH8yOs/yNY69BNO/mSA6tpp9WhoFsCeBslvqRaXQjSHkiigrAUEwl+KIMuCog34rS3Jx8uHRBs0
hTa2Nt0Lw6k/hZtx26efYgJxlta1yIP8D3nbZlEDW04suvznULjUMoDVfP+Qz2EtFpbSSzNKattP
6Io6MYosLpxj90VqJ3XfYQmF7DFuC/T4cpfFrt3SxSJskl1v9C7XJ7MV3oLhoSUV33kJGiBslp37
F6UKwM5PM+Lx8sNfSXIS0ukC4M+mDremQMJLBphDR9UExnJ766zziPwsN0ea8WnnCUA/wq918ha/
8TbEKK6riV9zmMB1GFk4eyjYoTuc7WJEs/OWget420HE7fn1Cuqm6hUKr/Csfd+W+m8MBXmarzMF
kSMJjdKaX/lnGYjN7cgkUCtTxALGzghtxHXsXfnXhwkJ9BVtUrxfsA43yYTbcz+mHwOXxe5/Qndy
fHyznLl6096DFqu6AS0JPMmuItOsGAy70jpRLbOQ5PA37suXIAT46xWTOGCHCso30aRM/tpi4SRM
X0pIlsM3c4EehglY7GE2sm63uQPh7idV4kWqZj9367NOqs1NL9DGt4fe/1vjuqosmlX1WsHtp9cC
EFc29gxGMqgdkpoK6myoz06jeI907NGC+KvlZmCwkYAZLp6VTV0tJndF1aiDEIYXiX5XB3qbldqB
EY4fksKCOY3myzy1UrcStcesG3zcsB1m0504F6lPOOYQtI7avReOpleztsu47oC6yl8N8OCnT10/
AVJtfg28S39dtsE1v62A3L/rH/IFbYp2LfcVM0gjvG7fl7/P4ggiJoBcrZt/ZjNaj/0mwbJO//3f
GvORsiZzxS8SBXjbZD/vgTxiEhgtaeauwqWjZhgMWvrbNmAw/bKQhGqe68x7oCmscTm11yWPvEaI
b5F/mlFGmY+HW8d9VwRoEuq/ko770lH5ao5IE/H5f+9Sy4nlNaoN0ehHcuY1FExMSmE3O074EFBs
htR63fKNL2dv/q2d8YG17G1wduTJrWzn4/3uAhjXSCkcMoEsTcKXYWKTu8WfFGgqRFGPK8Wl0CNy
JZe1+RtXzYjkVB4kHxnDzz07nfSlmEw2WKBG75DmcKOStVN9xaYQuBg145+PtNTQIk0cgrJ3MUOJ
AZF8UJQjc706WlqTujdSY3wP2zuN5Krdg08JfBC61YZKwBzo9rkkGn5SjYqazlcvIJDmcHqZE5qm
b5fRxZ4b6mL9RUvCHoaE9FuadB8M7V3iIaVAOxvsHEG0UrNEoBhbebT+VngHE6YeMA+1kAG5hDuT
AkNAMT1OgIba5pc00gm+cEgJuvv813DgnCsIE7wcWhHBY6b8R+Mslt9R6WhLy2FZOILuIK0XiJ2Y
WetGPFxP75sf2Bmw0FplMcbql+Vop8PRxOHHCrvCROrHjwFlIb9fFFnXh2jCtSAGF2HCl0A1XHZl
Refg9hSbi//+sKFGzzeaK8+fejESSHuU5HXI8wMSe+ErHDyIZJnOkRsDYTv7Bi69LEcl0G4Fhsoq
KkhJ9Oz0umecCmpU49RW3GaNK4kSXG73a++ISW8AWzgruGx+vcowyMdSfukqMxp4hLC66M/dfqry
4aD+gJ9KrpBfxRhirJGzBpocM740+hsJOJnp9i/OQt6gFOcgOEHTX7mCtxYjusD9w/+QRPQ+Xr1D
RqNfsezPrSneyh6If3T2NMRJchYIR6mzChDTeAjASdpLDyOoCS7XUIvZZbmOkFHWpeEyTLcZSAuN
j7t6BjxkW3dhGZln7XCDqLpk3Lp62hfOPmK7VrVwQQQqyvOdhLmGLW4nU/Hx1Vlo61aBhYaJGjK3
2aRjDp07kpLeM7iR8uyxxoTfduLSadrjLrMe0hiWi/8uMjC592Wi1fCG3VCqu0OR16mClkGpKIfV
zei9K8+ixLCFj9z6HkdJllI9rMvg6EXH94mzWeIga51GUNOh2ZIVlR0PO+PylLf0C7lwfGKr/gcL
r7XNpJQhGnsAnnA74mAOBul5fIrPLb7XQMVhp0ESLXiSoFEvJSwiXmCU/hQHabh9zJmKXsB3ozkL
UxTkdoSyeF9GLtX4Ndlpr3oM+EeDHf5H9brcMhGtIoCVO7BCRJNKujFeMaSFuKAS/hm+9qUgOTOu
7ymI3dKDHZl+tG5JwjifIF2y8s34aaseYvnvU0JJK6Iuc0B6hyXHNBJ6Q0FFEJoP2AF7Pc6CqcBT
gilxrDu0f2SmAJJA27sq7zB+nMX51SwmYnY7Ct55Fipv3vV9rzljCwltIICQJ1Yixpc5pi5LgZ7B
M2p9GkDQVks5SL5sI3OWzBmJp7xLPRcBwEVkKth+3y5+faFNlgFzM/q7ncza0FPJ7hkg4lWDMJu1
7C33u4LM0gr/ewv1IWwk5Wo7eMqZhQoEwcLDGe4plSL52rhrosroAEZ2emszq7ugYcz9URj3a1rk
vEI7yiR/xG505fdSDBmnqnNGJslf3Wyfiuye9lLVjTshzvYxCxKBk4il2zt0scm+1N0l/69EWarD
6fjzfs73xccbSsLoE4tNJ4A8w2DxX4TZ8RAty5+/shwRfXn+9NnwkUJsz3jYkcF5NxuIwKLp9ocw
eMZtoGGFbG/4IrbVEfljhRli4DHXnT2tGk1XbgK0dabkVkF/AtpsEkFZKCh9jWWZZYuemlS6oWqD
A5IAVwJaTAsnj6G0001gtoNJxCaJ+d9ul04H39rI+D2itsJfJzB6J7m/4ra0Orith/gUxIdsaerQ
j1HKbvsBGkTu/LC3QQyvpAXIPP5hCOnUx5DgKwzBlu27xEzkhM9Ea+aZJQhoVQ3MaZJX32Ho80qt
vu1YZhgUdj+IMsfN+qzpbT6NmTisDdY+GWrvQAUadwZkEDBlvtgNJli7qwyFx2MlAISuxhNCA7yl
KLCGuMr9wP/jT//8SZS+JFjMrwJdeEf4SnvBjNtAKGKuZqnvrOY1LtUgjjg6XFOnjMof/Fe14fP1
IBJjfB+y1bdlD3Pq/n4Po3ViwmPCvz2XB7AfYcfV5iFE+PT//QKAdwq7JKcIxQasBQc/seSGLDzw
fsDh0VseLkmuGIDLRQnt1b2Jb5ZsL02W0USgnZfhmwKtRrl7UHFgbqMTBwe7xSPCQQjDT47sxqS6
/gB74q2uxZkd2hSbv+/yK5WagA6SesFZk3KgxlZi6ezUR0LHNBZfZlJScWpQqSR1JOg0fOe0hB03
jhYsEc5wwtwt3RMM/fnVwAm0J7w0G3wagblv/XXxfYqM7FnXkrEWptECPGPg75im+/mTZodtuCdl
5Vqa4QHotRW+XU9673VcOJWzVjG1oowNN8lK8/e4Rw6FkUzC4f7hVOeKm4OzbIM7bUwA/Ou7sRUo
jB0/dHNfR+/rFNLPWxV0M6WKFjy+652GlW9GRRH7H9oVlgE15v7Wf1rF0QGK9vcW+4XGouUNTqf5
lSBTD1ds58EutZ3ZdTLY071BLomXDd2154XjsFWbk56hvKhEIlQdoAUq09R09nUajo4N249SW7fB
W2nTFwGWdG3hopTJruUso214kFHUDeZoO2jNgkj0sw2AfW2w4nRILoH9bxdp13gnt/bQVxttWTHG
MhlVsDxwNZLau8tLdNVYp+gjB23FVKE5WyYDsNLNhORtQih9qo48wtdDRxnA6fUrd5wBCciYv6kN
8kiF0dGNQIFCJL4nUIEKSiETkR3P+wHcfzFC0CWfEukkseTblUA7PVjJtPRy4XWClldslfzA8sLM
TLpCMXbIwdagxeJ2kU0wyN0c886Y83iRqK5YO1VFMuM85AGi0y9ZyO1P8IQ0F5vr28mewA3tqcUU
ZuzaVDyTJanSF2csVcZd/NL47u4WzF2jSRtV3Xkk92P2u4VcaU3SYSKQS9p6kGEhIpdkbXkZ1dQU
YvXdIV/Gsu5WAG3s86QFWbQLHYebrtJ4BLUN7c47qewFlMnAfNCUSnKr6ZDWXMLjp4/qW72C2Oit
HPTn5PHFv4yQ8cVBl/wrHqU5j4eCXQKDiCflQdFzO6TANuy2SykGmHs3FJtoRDf/+rhSCRoeBhUL
5ydqEXNXKxbCI5usAK/hGeOCpkgtH0xxNXDB9wb2+sTZQzTQDDgERAefFeH8nWUpvMikb29oVdEi
ElUdRAB5eHQM9rKbbqvHJxyv3V4e8mFWnK6FnRhCSRG5aL/oDYX+lsZpI001k4QieFRcV52qkN8h
ZGRDIwNzxJ4X/xctoswGw7mMlJPzADEhIXW1DUE4A2PMUvV+/yWNuzXxR1PmAn+d14mYNtT6MXxK
MhxQnW1N7NhiBfAPRoowKtVgFUY3g33CbQnLM8ZWxhsAirn+uS7g1BC44Xv88BBi+mWHYiciGH9k
9LePlCn7WTRxhRLHTpFUpYw6yWAUnO9RyeBLpiXINm1nrI2iCZI7G4FNWDFT3MOpje2+ZSYf8CWR
BUfby3FwKdEm29nXUj+iUO+EJMVZIalaYxmfZTXaH6/FUagfNg/PUCEH7tuDpD9u9J3SrB5OSkQP
Izmn8hj0GUajhvYrXplqvwCsyEKE77dY8iHohPhLpFpZRyXeZb17s7lpH2J4ntjaqt4+jb/S/Zu4
bdaYwFjgTgRS50qec+LbY9CczGV1EbnNI4gOM+YleDwkSDLWyL/G45iRSTdNm8EYfNnAVbNUVzp0
BfP3awuj7b8Shad8BWD4IGcX+OV4pH7QrVVRtDh2Cr4K8GAdP4GrZCKsgRVHMcrOwxD5KHod840T
YLtJBA8U3XuCP+jAYeu7beImFEJIfOZZPRQhBpHAiwA9Vh0VfSwHM9TPNIcN0Rtmd0IfkIB7jSIF
dsOGxeOrcKc7M7QPHKkumbMh1ItQTiG+IZDJj16ToAdeU6JXkjUHMknP9HyWc385Z8hheXnsmUX6
RCKHLmJG9tNp1hfNOek5WR3NYOHOZTkG/e4kfq8S8k/vQDC5N0NZWmT87b9QLVyzCVo7VGUqCJBW
ke7VhO7U0ipzGuzOKRIFf9yJDGNwqYHYiaAGO5wGiTvMRhDjt6qPPNXKXRyY43JhG4zsthej4veN
faNrOuX+uFWNGJUFJ7SaECJ36CU4gn92S3scJf65bpjV/xZceUvKLYETDW0Z06kwXOE124AGfSyU
VGl05vKCQy5yzkzuzo7JJeWkPwbfRcTSyveXCaqZ/gieOr9hEkOT37UOw9EgXAvSUbf6m4JvG1u0
6nCDluvKQ9d2ORHCCDDCUzdWE/298klC26lKFKOHZVq2TqGPXk+YBSTYk8MEl7I+KobPBcx4RJSE
i/rx78Uef3MS8n+oB2NnEFl/KznH2G44j8lprfuFNqyWypNCM8pgw6utOlhlEjEFWK+cpIhWhH1I
So/3TN+HM8SUhfSYzzWG1NOgROC9unfEqY1sctA/qF6e7+kCr7WTajeJtXeB03I6qikp3Z5gtDyE
KqOwUSNSeAJo+FneKi37ax7wuAIbmvLRNDgifdwSbB1G88EEKbebV+qQ1ZJgpfNtAjUicMbVekgj
g0+x99W66eDATgUUBalyg01OuYnaxe+wEBwgT3CSOwNSqZwffivgxzKUaPQqjQPoDSnTSFDCtjlC
vYsP/n+s9S0lAflPJmco3FeNsBpCD9+FgQcgxec9XmVcVWhhZoasKTlA9tGUjpJzMp2+QAWauDkO
TBdWjRyOAg1KddPAtWUphzNwjjT5bNbXzGhVqQrVaFuhMPMYPpmlb+t1WotMc7BQx823xvDWnXUl
LFs4aSXKRrni5UXtqRv+BgAdhiMNbaEQUi6y5QgHmcbMkn3lNyViA0Pl2R81lUF65dbfMgzthf3F
hPXmGdGqRnIxoDyFkSY2+eTXuq6Ak0TWt5FXApfuVShbrrvhFiPPPR/fmhux6QMDRAaUqbcF9W+k
pk1+kYvPhFkg2pLJXmVHgDQXtKE6szrBCdYiBfVrGM9NUmR4sBb40AlDyQtYXE5NeBQrFOHcpIzO
gL+mP/pgV63j2R9jxq3HPkuvV8DuUnighQF6jHmZ44OtLpggnDzCfeseZrqxpvifji9H9Qvjxz45
I/o/ATPvWP3heKKa0dJIHWgVtx9/q/KIGNbgfSMSujixPHa7cRDslK4NZgYSIzBZxzq2IRVu+2PK
RaQj1D6RQDwhECuwvKyF2R29182TmaaJxRzLvblR7aYqiMwgfaIB/mExJG+1ts17eCvAQ4ylVjgD
T4yAeUXIcZ/e1LvB0b1K8orcG4tJrdhA6jLqjKYul1Bt8qflSviPmuhzNbrvJL7v7AD1DgMwG6m+
OtcMMACgdXNUpErVWG6RVtczCBNVnTppXxXdTE9ORYj7mq7ee67wwD25VkH3t9OgbP4mJHTb6OHt
eU1ms4hVv2V6QHVepNQIDGkHTAf5/cxJ/FxThXjm3rk6DD6yDiSa+4Qz4FZoRcKuB30/FJEVfZEQ
ZRMYvXnxGzYEYNrMMMrxgdwWI+WzUnNu9gXtu+XH6H9G7nhqbPejyUDmqyrIS1H+mavokeuadpHH
94M1pO2m7L+aQ2q6/EGMVw9mn4BVC7Eh6eN54MWGpDcbZd8a9l22COtxRh9iT+KwUf7XOn+EkIic
Xk9OnZKLp9W9DknuGPG7IyoYvAI5nrwz1cgaBJhsMnZfS9zAb/u+Hsp8ttXAR5Ie1ZZQGZBi5IPQ
8JXlxG7vPnVqg/IxSURhEA9oUGtK+KjpNaTlf69acEO3NMj0chiGF70QX3rBhRNctg50mLhk8/Lw
iuxOKA5gGRT9RKmeQDLNc7OiNvo58si79jIuK/cBjJtHJn0UTzUw7jhPbLGPxJFVkbgw80mGFEL/
8TQrWgOMdaqV/N1Y+5LFHyoa0aLo7Qy8yzZOYwLX/06tMkb9GInc3LAXkswkIt0kA85lnvvZLiCy
F2q4REIbbgw3stXzisH31QOUYkkRFholqujvO54T9xTIYExC8Wroa1DZO8IaGc6hvug5LjZQvtuO
6ayKm4wvF/leqHHcdGrVzrMPWj4dqigmmzH7tZbNYC3FZEQxGOnym3DB91ADYCsAXqaIbwBXywTA
3GOmLlAb8OceAVQwHA2ogXCt75G57xtH0XebmU+oLmpzsJVY6kTZYXjXt54ZQiSn48J/5i67zEQp
dzTZcokPD91QLmMuuDrHRou/Lro1Icx4U9ifTTrUwcfcROj//GPsCZWtHXeXi4yNyPpP8vLX+F5m
R9cu5ZXt19x7O0Z8Vudu3YebGbjeKRh6Yg2hk1G/aSAHsxZ0gr1qSFPdgHPZqTv1/9vaOnd4J85f
GrQAEkyK2zzAZ91VCm1NcWJbZ6u61nygnu0X633L/L/ht9ECtAO94WS7p7tjcOLJaNrwdOJkQy7A
SpnWagf9LzNqTkqNTqr9zLNMz6wV0+4wuFy02yo5gCAA0hjCx+m304Ny4EsFsHqfVZBE984d5vUg
SjBWv25If9zI58E8EzftxInBllrPB+GlwnCGlP7YXqB1LaeHHT4HFRKFAOgWZxx0p48Zo8lyWZDm
VfbWvJBYhmtXK0IOv21KZg+5iBCbF/RUlxztgUTmh9TX4FNIfsre4b4WASzWoejH07sEQluNf360
fRzqE11cZkf3JhnO6UqkqNgfIk+QRKa2ue7LqmbfocvJxy6dzumAnXGhq+C9vPi8q7EWmFvNYj28
1WvUnWywphfiklzbEPk5js+o71/vsdeVhFN8YVCRoyL6td25ZV8tc0L9AL1gi408V500TD2O4ICu
QJy+F2wBmznh/VFVeE4tg95xwXpRZEvLxs2kiXNWPzyFueJkkCoMOcd/51YWqNTCaI/JqOqjd9V8
lV1gBYBUKNRNn+Wj6Fl795c30OKez+a2ysE6W+gJ9tafnV5x8uROblwBDMEy6KeqS8z1jfAt+T75
Fwinq4HeqvmcYsy1HAmorBrZUpw4sRU2Xvw6lHqmHylXXs4kZTfK/L7182PWVT7zA91EzojNSxXD
Oq4eZolduOGHq5t8tWWZaGldE6+HIT4kD7gDPUS2e52fpb8HuPKzXXof9pLXCk8Py8aAJM+VPSO8
IdiggaVlgOojFIKr5QtpVFkclgJI83CUH6KO1C+zOtNzoDy6eLYS8pJawmCCLiGNmXL1ksXlsQAV
fy7odvMhaT8fcNqr2Y1sezrQArYsPr0SX4akdTeETPzSSBgVRnnNjadk15Po+5+w5jFWClET0S0S
qPjpmNkANc3NC8KUmO0W1vFzrzyXwQoRoLE4aqongfbIWt84Lr2V47+Fwh0gnqsqGlCaMFP6RxzA
5V+mfDnbiPshAPV1KzgewfDWDvyifE4GtKgY/yMY9E9aomfKyT/cB5IsVd1qH+bM5cD7sgFi3wqA
SvWovq9+3tiicTyCwNmQJMQFBtDforFdfguxoVb7iPAfbr8vQOOSpdPzerC4IluRGDUqq6ISoY4f
HrGFhuC1wFHHZANLiW1+p5M0hD+EC53rgnQblOo/gCrfUrc+gErA4al16k86XWSMysm13Qlb/yw9
wuLb8iXFOQlCnN9wGlzM4WzUkXfx0+v47YLw7mTeJtyK8gAxh8Zc22ayuydroRuTo+0DUDmBEP9k
uUzqoM+5eDyJOZyePK7F5Fe+anaBJ6IabUnnWOUinF4WUd45wO+7byI2JQbT5hTEZDKgbSXLDI4j
x8bgtRLQ8+bADNl3gpCpYGfNn4WxSHAdym5J+oquuyPV2DcEid7Gy8UPyD8qGGGoJpxWI03sBopv
5VJyoJ1e0QcbZCn5O2lGp7uAvGOh6BwW9NwpBhC8vN9XOBkrWhB/lUW6yF9Rl4ZwaW1Nh2NQq5iL
JlgFKtumZB/BY2fmib6G3M4em1JmyrCN2NkByOHgwE1PXZDvmnToHV9QVsvb6HAxSJ2E8jTUOBJ+
18UC8VV5Ofi3T8jTyFpACrXKafYf2br43KJZpqN/dOKzzeuXJTKlWvpebMU6V4pLeN6xpu0/095F
SKDgOGFlxkZNS/FoUIvusoEPS/ZcVEbUtEQD/Vr/dqvThraQgHE8ZZlNDFDzsMVHqDoZK7uF1c/O
mBs0nE3DsZgYo+JHAADuka8PyT8FJVTJphry12/HX+xBqSXjIWGwRdjaqjiEuFRtlELtqeUReLD8
+1hUcj/Ybehs/cVaBn2VcxfxaDYnUWOk5sN4wda8oAcFcuE34nPil1i6vT4rHh/isa/vYllYKSWR
VXwg44mpx0rgQbYDb8i3MPxHbC/yMjrM+7zZkWLz0VptTg92E+jXwc/hAoi4Oy8+H6vWcRk06wkQ
D2gzdJoMgRIZrBwGCWRcmIRPAWpuHworESoFIgu5fFvffPuHtbyjn0oNrZSO6/QBb76etkkl3fTq
O3IqJYN9URV/iMA8/a4Q4BQpNWQf3xXfwvLMycXVWgM5opggj1+s9u2OTbdmXkLK0ICwdUDNXsW7
3R574eaOoki57RoxEzyMSkhnDym60j4RJnFVM+5N7NM2vthdpPCIq+x6ZsDBD58VykaI2GezmZ6j
5/o8Tu0hvp8/NUzCKZR8Rc7ap9aH/vrvxfPVNchA29FhAKit+ngI5oNx6IT2vGCe3y7hYYzHNKzI
lbpQbN+raIlwbTHjduMXCTOzSAo5pF4eRZV/MgMLpDDRVgnGVAoChCoDadQp0zq4wt0pWO4M0FIX
ydt2MH6/9zJGGreSwFg18tBZtGz+7WOwnwHzJuH9husK8qpuw4C8fey8JhrjGwaszpO5rAwBdrqE
/NRVird0ljn9Aumx8/Z40xFt0ilwrzCznGZxoFZ/cw2K8hnWBs/wW77k1kntb8NLG/6IIfNB7jQd
6wh8WXTHKGBk+uva8NiEc/v39gtU+GvesrBSZ3OXB3vIpXuLkr/4FnAaHezF/DcLS5B2SkbGN02u
4m+iTcKkq6UtBlxrNStR41Usx0vd+L6hzCVHACGnJV1+XOGjyuUjBQ/iLsKYduLSd/HhbMUby9cK
NzoeewAyzM1IUZXbHbQx6+schMXpUJzco/4PExb6OxqyZRlcHkxZkepKfcr908UXSZ8fyQh7whNo
T1+rIvqMgmVaPPEq4BOr7IQTnidAUjmwb+k/c5oWIkBcE4O3PXeAmZpoVuYPp4+Pyf0HSUo/1X95
a9ciDsz15YqlY7O6d4YeqN8ULBauIdlQGxnKwd5YoLzLPcf9zDMDUvdLsKrwmjB55ccpa8Ka2QZb
gqUNf12h8gMTDQX05tXx6ugpjSYUXTCEaIgv3MAJSJv5Xdpsaqi8Y+vI3PegbfrC58h8BV9C/19M
sVQ2zERa4yy4mT8T1ozZKF4tLFdIYQU39EY4tGKjnS4HgzS2hWv0lXEIDpfDDcY+L9lVxdUq2q2T
7L7n8jdTYuKkw1NjrE5DAZHBS0TtWwTTYAJcnjEXwrIacb/aVbvc7qjb7FqI1ci/txoyhl2xiAIb
m9jnKdzIVBByvttoN9BXc2OH7IlwRdXFUwrPkC2IN/ug3+B2LwYBeRSfhHt06XlTwMHOBTU9jv4W
mCASNhU1KcS/KiW2gQD6oMI30Hs6ZnijAzhOy7LAPhTxWa8RGKqr67PY/ZYALq/ZXc4UYFCxkBKI
9G9cDntaPjGmBmuHIvsS0nizbRHZNGvtkyBMTf5yA8kH7QjsFcnt2Cgx7U65x5Yqa9HdytQKhM9v
5wQrnwYWOub5zET9YrdA2iYXr3QWRdpUgAhAVW6UHo0TY29oMhsHf/nF9LAsl3J4O8lu26/eDzM6
FxxsirIlWmJrGs+Wo2ZHpCZFsxPqtcw2DMcX6i3DYp3CZRfc4VlCiOd1mWdk4lvE7znZ0SMGfhvc
bLPXkYrEqHw3vec/UnWGdApexg3CxY+WD09WBh8KUK94jG2nkTlXVnKWLCfBSp14OAu2XhEj97l6
Wa3QikJDRjJhEKA0XC/Ew44P0a7NI9oLMWGw/8eCo4436fdxi+LIl1TKAe8ntSXjo8cUuROJPST1
ALtOTr4ftnk+8DcfL2BhwLJYn7WllszpCWGrWLOp4ciTqMkKlmoblbAxjvbbxMMFeixJlEypC9Ck
eUfjrdzb/vhZiw0YVvbwTpfD7Pt2XziB0HWuOSRSmfm8LLPHXxC85v2q5wfddHbP3V0hKyOWRsZJ
QljKfdfl5bbtdxF+3h8s/SHVn/LsH7QY95I6dDQF45ELLwMczauV31shnjPbbbWV7aqj+h53Bdhw
mrGja/lZHr661XnTbDHijzsixO/jpG3i43r9lQzbCUhPMm4danylLPFPvZ3mDF6XGT5jzxGm08RO
mcB+mhAwTkSg0tp2aZcix/vnb9VnnK+gKo+Y1iWvJvoruDjANfgA6aR+p7gn5j0hQhJnaSPaWPUB
u4y731BQLmfltYMnOj5FN77iCC1XSKhEP+WwH3S3sSKDBaxIRR4AAmI+if9DVMbtRy32GDG6TQp4
KtgNzidZR9zLQoYyek7t9OCRxDiRnsceICaqNFKdwmN9Mt8wwUukZTZ2j2YMezE0FIT5wrTCBq0C
cgulnE131VSNXgHTWgLKb2IKH9ZDkf4QpopFvccZFgxnK2pFOxAg6ZaOJ1pMq5djx3hGovjoUMso
UZF3//asDVQ0rZ2CgpwwsVWw3oPEdkFzjvR8qwDXtPKfPn+mhebn1qZqu0uSSojFgtt+V9XPlgDg
q+tEc1F6caE6tSIDx/X+9JVtR8BacHEayTd61c66jxMPZ5Lt/bcWB1gWncfbD+hpEN+jIm7w8aZL
kDZZ9JcEcEwBHUJDyZFJLpg80/m4CVkR0Vqao7X1drjLGrpgfWjWUsxV7LXFX+fD2Cm/CbmXzGiA
ZzKa3HG6Ab09bdTo2QifwXGXpjERn9DNtY9H+JBIdmWq1Wqvsdha/0tvJs3G7glrSopX6hc05Crg
SrtYBwWLHuNLAod3hvLmFe3xJZpnJG5xaF+uWermoeY4QKZpQqmC1WAiYiVuaE+HBaQdKJb3jN+h
+FvloxdMeJlhvHJKAhLZCEVPrzOSdeeqDssxRONbbk8mm5i3z1/Ax3Duw5nSencRmrEci1m+/4qX
PitUSdGQL+wOskB0uus0sdUi87NUCX6FoXMJcVbwmj+GsoSb36ReevgLRU4x1Y7TiG7Cz1Z1KgNL
9OGwFnZbAXniTLfn7CWf0STg3zalmnHIaLTE+32/BXYwd+KiqWGtplTH2W62Ab/oK9miHoy1TPOu
2kyWGKMJIAKn2XR/7KfbArvV6kVz/FvELt1r9JAwVUECytfNC5DixQWO+yJQJJJZ4ACc9Da5DVmA
EAFTGSaoOC84GhBWbjedmEQ4j7xELSUL5VBPRVhV40S+JrJPJvL0cD0G7V8YRpyrNK9gtcH+mg2T
ppqt2a0aTyKt3yYmhYHsXH4x3oBnbR1oGr/MJspj2nGS75SyfkMq7JPGdsKzhNuoMGW5MBk1SS1g
vy/fwU8D9sM3dQjBlN5s6lHDo7f4reKVYWwWzPJUj9fy0yDwBX++H3FipUXVaCWG7M2mTLlWVdPb
AlCK3QPetOfPte/Rsxm/T4WCgpVOx+v8xsjSTzZFMtcn7akUHRfUzrAmCajDkJFblwKUWage+5Ge
A/M40HVncZCj6R/s0xpxgfLkbE7rZH/4B4s6yldd9MJHIZQD6Ft53e9kfBtTgOxiIPI5/FtLQ/Z4
wn0F2gla7DSFnBeVJwyPhZn8Ix5jdeu3JH4PbnKERAphgugc1VsHsnf68xRUZ9Xi/OnUFpl4V7Ky
hTYiiPfyZy7KbuNkw/hX7YW4hx+DXwF9HJoiaiDqYjlR+asL/oRM8NoDiDUHS1+kDbo7nvS5iPWi
rbI9iUf39ti4MvNe8X3U75urDJ7WMPGc8SQgMEW6UYfl2DI0zcigQCrYPR/oLzfqknldGaUD0Def
jE71a1wLZtpVC/3gkQ/42AvRm8xxkMqvTFqsfz4ik7oqZE4X3gjQacRLcU7UG2sNqQeWWnyqRiUd
nHtv1W5nGYcTZ6l0UobIfdM+JaruxQYOGA466omD+sLOL0bH+sUwKmr3vrLQ+pRSWvXtLPE4ymw6
GV9y3MnoXn0qabcfp5S6a/oxz5iuZ7oG/MmuOmcayxMBkmIKA4hnleYbTdWabuIgcd/NuSdkMWE7
Gk49MwPTI7t4whLPl/0FKHwbCBck0Nv6Q8FxoeXcrtH3VaTvT4aio8p1nO0oPS26gPpZvEiE+Gz2
5KCYYpxkBncNyKROgh4TRPjcNSe++cfKrmHtpRq9P9+X3rA+5XUxS1hE5HRvePITyxXh1aH8Aafb
J8rGo2JJmpOSX0pNWVIHw6oD7cPNAq4p+SkyRsSoTug0vVSjxRNjs9odfSEqtWUgiH4xB9XKeZQr
lSDvKzYtploEmYijR7YFJGfO1Hmo13UEFIHLcpjJy20kSsLNYxY/3ctYXnddlySKmEnzgmGF6Y0+
zokfb/KUm5+3Z39TuSWqARKyRbr1EX4RvCL60DxmbPULrMlk+1oWZ63LmAVrqp12GjO4DwOSlO/r
dtmAFFwOU2q6lquIJRwElrXet8hl6FDmxkOnytMJb/0cmg7zJLJ85gRkbnG5qj6sizBskRlJDapI
hAuo8XawQSTeaj0MSpuF/hf9Zb/ViZSwTo/Vn4yWews+aSgngJjrWpwJoPDYDZyyOJ2mED/KPlKn
mb8XqYq62/y0clGHnWZD8D42fc/B++FYffoATgqXL2vDThzLR69j4RzDjge5fGhumwvKIIz6I2Jg
GT1gBkF94yidYTTMf+5VXJqEAVv/NveGxQW2Mllm3AMTrH2zgd33gI0Nh9h5pRlA/dL15VGyQ8AY
Df2ok36Tlo5rFwpi3nvIpxq5ac/6AsCVbd/UVaYUmgdia2oW7GWfYksArhNo3hZfNZMfotazXJSm
pkPYifQ9YldPWocFs0f6OBvhWstDnQxwLpCTb8JW4FsH5SKetA3qtu3RtICNjYXv3uNAtcvDZnh1
AtEZeysoU98tgDYRwZmCqVlNpaIfc9udpZ2pJqwKdrlnyl91pEosjChKeUMwTIhpD29tmDF49gHy
vjfDkPyIgg9zgHS40fYO1bQfF1GGLvWbVz1BI99s7cQpmgIERDVV82t0mI7bVKBPdPq2yxqr9vpw
cBBvrA0C6q8mgHoTarJS6w9QemPFTJva0EndfbzLyvTC/6A518VtTAK7d4/3kjZDAUf9xFJ6lW3e
mQL6UDfdzNcIT+B4eJkEIcnvvX/s9viN6ZOneOoYhWcGuUBvKH5k6sd6D4S5M0u1ypU2stjoJth2
gHHFW0HP/ahGwu4HS8dcoqF+vMQslXcKENve8s93livLvShXCUKmyBaDr6+XZhDbMSR6FQGu10fU
HAp76sXwEq4kIuV1t9M4FBbqxxjbaZyXtWz3tCIPlhvoJhXCkGLe1LePMDnWqR/NVZAN1f94Cq4L
SKFryb4zv2HTWD3mTWgy/p0ktzYIDQ/NTCmA3n/XfFrpsPxoY1CAYaSiljStVygVRNnYrQV20mFs
i3tTYjPkUxtUT1QMQ3w5krxdDoFaByoaIWhs7AwMUrjy6syWBqiSgw672FewKL8B995NGe5VCakD
AZyjXF02CdWWdp9DYKw/5KFbTUenuntVw4Ba2RyBe/8un4NYhtS4+9yiKC71i0jUBTrIVHHB7NNO
qqmZIHSMaZcVXBLwUduVIVEv0TVFLzvBykxm3xUE9IIsbBJXbs76VClLSYwaL/Mb61wTb5KPAh4A
I/NkD81foIAFf/m7Uv+WV7eJKZoZ2RK/FeqV5h4yxBqMu3SJfgjyK670wL4G7mF3Lo6ajq8uDoJx
00XxbBZaXBqpkJrEHrT0XBbqHftM1hjcJ8nQuAZD8O0N00l5x6MA3SxT6KttTxdgTYJEz+wiziS+
s1EnqJcpAQ7NKdUwH/fwG/7IH635A2FkNbG4v23LbU+uL295CPagvlO/GpjnBBrrrnUqZHk2OQ8x
Pa7i6CWMNOZFUZTWjwTTPdb1k3BMCTP6oT4E8ofJodmbv5SJ8lX1y/g0OasJ9/OVqafzCnTLSYZK
4ilnMrZm7yJEKXES2BwZlNodHrIHNTBO21nDXRVDBRAHcXYx4arPSICtOhySOBWmmxJ0GVrhKh0X
y6Vb2E/l2Ou0r5T7DbM9Jsc7TKnUn6mT5Fo60LU5dBXmSIO4kgU5nVTDr2ljnE7SMuk+BhFToiZy
WivWICvMgbSWHcwz0kP+XLfr56EUyO6B7QCvvZ5F6Qiax2yIiOI8Ua5wvj5RvO0fB/K/VFuQwf5l
pB/hLHzWP/3GK2JWMTn4AJtOJhMq/vym5ec5fZEPToLdoPxS5MtS1cY3GUIvEn2pD7gBZrlUgDP8
bo3ob7vyOERA9/m/kktbI3vGgoz1hUIkv2S1rh2DYjbwxtH6EDMpDCI1wOKlO5vpPpEhWp0aAU37
8Cs8Veb8dSzkECYBWaHGyiIoYJfuMak0qb2SBKMbI96kYCg6EHl4apGy3YPMIxCZ/qUXbRJgieDk
YNFZ7AjnrNLsifSYFCaSF3AWo9hEL5tUug8uDz3y0vSB3t1wdKfXBy0Zoykcf1K4x6F9CzEcW4be
iGN/IMkLVyzRk9hSi2Lk7IcSKeLzw1DK4ZDaqwS5sIqIiHndJnoBIPzOa0h4v5Nd0sImA/OMkNtU
7MR72us2ZHvbqMCZVrbvMMy6r/d1WHHkjgM9wI1zVzZ9A10isl/M9uzI9mdhjTKe12Py099wKCtU
8PFxKLplhVbmOf86cqoYK2pW25i1USl8ybwgKP565azwxcm6CPLGwNcd8FXx9hXqAkc7i1b+P5oK
iAQW8wPdbkkaNuSbrdtk9hBNtbEOKd96i8/AsMwLp3grF2/a9K6h7FlVPKpCkqUfWzkuBid779zp
n3GTaxMkKS4pTamkeM+1nZ5XosVQ79qWCeBXwIVBlD6X0RtiSTFG6jb/4M1nywEN2c+MxGx1UgCg
TW9mz3z35cChiNYFZO9cchArXDny2iUW5EpCx+fA3UFUz658cXvRWpY3I2ptRlnUIDJnAd8BjI63
sao0kb9Vrt9wIEMRD0MLXyd97HtSBwmX47jTpiyGKwQ5cqUdhR9Zvdf/0I7kVOeA5lQmV6a35+7B
IMEgDi9cHbbQt6A48nRU5bQ/DiNwSTjVKB0n9hGesX58M0BZSe5aA11APJxxacqUKFzokDm1oNaC
f22oShrtSqRw4Jfrzl8dUqNRgJwN4s4c1fw49d6WapkFEuUI1vzNJ47HRLGw1TZt+e+EmaZsgEzf
SVMZuCh9T1GbmPQjlsfL6kDGUObSx2+AVc95J3cNJR3sLemovyI1WrWHY7El5GL6ANqtyG1Beunm
M5qhORyLOJZSWc1eCnn1NReBPXk6OKlBgd4evGI+NrOasjYw1ovyWRRAxyk9xGhom4k+EADfEQjV
garHJhIMQrhPWreDbBj3kSZWjrNwan5gp6EL8aRIiQ/AQbG1Ql5ILAVUFpinyHPHuIUa8ds2JsIS
IoiXIEZzrZSFo2Y5Dk0bEbLa4KcXegp7rm5ZP9IdNTUJ/bkDPblI3ZYjxBqdKsUk+EnIh1hXwRJf
7coqmJrSmPloWDOc9Fnxxr3DcNZOK+1Wwb7xSxMO4hcL/00rFRcKezup73U6giKVTRUxnbf4kMy0
ZWdCVgvLuVMguwuGrc5beAoLAWk+5attVVpMequcoqkyE70N4io+2ei0mBzSxh0c0BDgOThhxSQd
NStm/lhcXngX6ujAJ/bjmteUGw0bMQqrF+2n9a7iUpR9erwuU4RxDU77N2BJzb1cvFPWc4H4073v
vDrM71JxFrPEaU3I76IVUAe2iDk2k9gMPEGmaJ53A/9AKg5sqgzHGwFEK/yCTibXqcVrGRQzNnXb
t19Pu4u2yVTXNtAHlThS2wCbBjFfOHtP/cvnzANzTcCHSZAeVzQDGWgpqgu7GFw2OeeJXTb13gOQ
mf1FypLG8rXIdYvtMRvGZUlI8JAyM1MZR2TaQknbMBqAszwkv7757GDVFOJmaEeNfGQL+WLvXzJ4
II12HHugfweXdXAEY4YM16gXOwzfPGJvKUr+/cWYT+x9ugrDMXCXdZIP4uDndlddPh402gDfz4+H
OuiyuNad1+jwrk1Aqk96PqDLoCmndeUSWRvWwdsBXGpHXlQ5RbQgxdEIo8QeuXzsGwb3s/jxmiHw
hZzCotj74moZ4V7NvciIeV9YuoqiaIopKIkGk1vURdamQBZ3ka42n9iji/akMmE4/QLIQR72oCVH
RTrLfsUz/1SWXlcj3V+KfFjt3QQo5QDo/1Z0V7w1HQky2pkOg0OlaP9ARxJAiDi/6rLLKJFLr3Gj
sJRbQpw+iv4KLIyDAALk4tVxs8vGd2YQjWRLL2WNdaKaLpgkDLVujzQBT0o/VEJ0saEcPOQ61Nyv
KiiU5nIxxeZWxkjA2zqaBsODanwG5M9+uM73NFPQPUWSXGoPBZiOO0zYE148luvH7lhpg2qOxaWK
TV+gH5M+pgf4n704o9nGuQraLxyU+LRk27EU1ri0AC4KaYjSRUMfWRtOFjNMMa4uu9nTPIm/2lO6
pGLPSPqNi0LpP4/XMj6u6FHRy9srUORb2pTazafNL/Jf5MJU5WYQmdYTZeoVrnLRiv7RZesyxIJ/
YW1LQnOoVEbr139A0yTD0UfufuYw/EmrQ/8Q0uV2d9lrtRGAFEC7Z0XEUjelkpgVO7TYaeF5LDNL
jnp5Tv+U44WGkcgm4ZBN2tSgbzWMjZrWVWoWPrvoiPU9h03smjEtoO9Nu9ARaYACptlh7MLfcwOv
Pztd13Qy67LjUmHH+VAHGQaK8LcNkVXXCaYjSt+JgMG/ZauyVz2/p7kECAP7WjAIN31GxyHSk/3e
VSiaJGdfAwyVDLEhH+b/issxRgG0wPHetvoTZHAPAvPfqXfKdAocbi0gxO8V6snPXPeU9OvHi8Fk
iS2rUokQvCSFwhLoDRwYprmN7lIrL/rRXcPPG5RFEtT7+J/WdrrUSACU4Iqw9mQidj/kzkRgKo+m
R7OYsxf+FmS5RBj+cxfiaN83f3+vd3sNQ1kXwR0os8hajJUkGWNE9vDld3uDnANADZKpWJ6jGfS0
efMDB7fqNpynVhiN1jkyDK/E30NNsegx4xx4hpaJr32/6FSs9hIZ5/UCoJVYALum2DbZCm6xIVS1
t002/zF4AtVLB3InCAM0z+o4j0lPSwdgUkLP5Yi2famqAh7Ebt/CME+N/sMaIZKurLGS1xgmr7T1
107KsdyeSJ4lN4pg/TBZSt5I5VcEB43X+x5xpiRAoWhEfgtOvAYrIYi1ngOZFRHGYUsa1ekzeu5h
nOZps/jIn8aPvJHEQlhVSxN2vdGAXPhrzHthRHlHOov8qOWszSUvdbqYl/9X9S1FpgcQUrlIvI4u
fP0glpuYwgV2DryrStdepK4QJKhX7Tej
`protect end_protected
