`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
PMgDwTv025B/YeylYZGbmxtvX/ioIU2nnCoNdr0sODQ35Lk9hPw+IGhw3hfnyGom5HBsE+4jLndl
9+alL4rk9w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
d8A9jmgbHGUrgdW9r0mG2z7gcVnjMYF5vFvL+sXJ0arh13/0VCpUY1zK+nmxqXy//XVofATvnF1M
KGZ0u2w9s0+4AXCMkwF7z+tRyLmfufbvY9j0bu2Fy8BpL4dL0pgSDmvlIsJ22vfZKll/ztx8oRKC
p42B6s/m0WGnsPf5lM0=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
coVPPXqglGz6mew7NCODD2UA80vDDtxircBCJALlgA/l0WySuPVhAhYpOFcItSOMmh4KWaq1F0qn
B0kgpw4n2MB0dye/VK4bMRqup81rlfOBTFyMRIlv3DWjrc79bh9htvw7rgDmuzHif0VAJnHoaJM8
nLS+56cDpvXl36t2pckud6UUaUry+ltDqHkh2Ye+Y0oBJDtQVmjcveUAtiigfWnd/pJ4pwYyrwM1
EfeTfNYvJhGmSlFQ3YcOtJfjqQ04mVXmnouFQW5uwDYClE2WcOPJPHjz+lc6jvfOngdAPPQ62SxD
j9JC/yZTHDprpYUTG6rB5B0ylQvzjxq74szrDA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
OB7AzV6ri55/pOp+MhfYmh0CETeYYlkTjQd495yrZFbSdYar0PzCYClb/a4HIV4RnR3Jq/SUBH92
Ku/Gw0UHCduw4Ugj+lgEU7vG37pq8G4G2yJFxTDfYbvpoVzS4NAm131JzmQiZsTZFZeVYnbGeIZV
BM5kBFTqal9+2A5wbWY=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KRTL9wGGYX9nZ+wFLgO7RDw1ThsgNfuYZWgrwImdYe0VIBW7HBFSGzX0W7hycMD1M+hW3/+muq5a
9LSgGeCB+beVafe2MEvmOrZF246icb6k0+29n9rKtXEzZ1IZa3kGiTWktQuSCjq5TyD9B9VscKd1
/tW+eKAulFD81RMboZgsWw6Fl6/ciGdGIL/E4h6X0Y1seXWfd4uCBHN6oj7ua7bTeO+ovYVtfLkM
5Avr8ApwbhmfQiByVUjkqHp/K4XVvo5SkioJwiyt7Tck/0edEv32L4yUJUrzokkieBJfddnuOSf/
N7zQ1SJyaLL9WPs6vKBdKFzXYkT0VhvpA9SmqQ==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Jfjc365FdC/xUaX7kFURmyzVCZ6MsV6NiO2ygH18eEniLggrSsIhWG0nn+ArZJ+zpsE8uxL1UP9K
PHHckCOZE32v/jD0Az34bHRsn3e87DdjpmJOjc1MArn1Hwa+dXwi10gZZgY1POmd1gvQGFnWlVkO
k2By6C/tNWVDG6YXMXmCteoryJrsJUhZgl39McDuHHpRm2Js8lHAFJ5bbIU1OJZReppc8PbI8Guw
CAG/vk0e+iZYZoIXXJUvs+94FUdaF7wOpXoF2GDT/cKmEiKdfn97cxkfVoUmjHvNhnVZSYZ0UjKr
KUZivnIfoFedTX3Sgo/ABhf5Dek3f/TtTn5Y9w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 168544)
`protect data_block
yF5/qmktyuwhKPJVWT8TA0BtC2m/kRnBEJzFqwgTCq6WZe2s1DK2v0F50NkEQj+2f42DOz19GA4t
Lrwgr3tubHFXVfMdIJmHohy7BJuz/0EIj4j10DA/PbHWh5eaLKxhzQTnJZtlysQsYi99Py9io/qs
8wMwCnRrlJAWN8/ydR9+DCIPLTu/QKZYID2OlhH+Lz3Q1jezceDlTKbGELaVljehdQncsw+zjAH4
S2SLsohwZXx5v4rqRFHSCeLk8ywBCkb0ZnEHz2IN57fDm/0pZQ5MwCrC/31yul2CH35HG1kSdN8a
kZriLehm0FoHVs4VBf+6lxwtTkLspuOSpCb9KcUfTP15IToCeBmLhwl6tisyMjygO90F1xS5n7Rr
xTv85iJgEQFwQvzCbU6E5PmUdTxgohnCn4TNCnaflCJHlAfVUSv1qevcpKMiKbG+S/gJd24ovYoe
dWppRiE/DZg/bVwXBI/tgyMVfAiLdm34a7rWvqdBiB8kEyTtEX6EWWP5VTyAwDLMFUmywY7VS1Nh
oCAGrbVrVs85uYEDa230i+3lGmg1+7WSYDU7Wr4fxMOxRnyrBOrMeSxK8HoTZXvkxKug7tmr1kzp
K2k2G82CwQD+av0RFC4M9d309Kjt/QoOLN64BX4wnHX4feKK7VxUG87Ch4UlbzrbBQmA2IdjZZA4
KGSw+dL702g/0aUifeh7IMeKBqYv+Ea0i0wFLi3fXXCgRkra3X9iTG/DNCyzPWjCBnCx35blVtfS
DH9zOzmr9+ftOi7Ng34m4hDyKJ/ovmY7FnqM9hUavEFXlZ0MKTDGp53GPc6+kIJca+heAKbVXdgK
ZU8XHh61fODtB0TNvwMlFkpp+7xmr2+Omqhg7g8sryaZ0FpbLEUlHBgMaDaxE/CL1Dfuqps+6Ltd
bNadOs6ySh4EORZ93zRfLXC40Gkhjlni15Zw42Qd6PKAr/BCUwVwxrFAdV086PfGspjEwjuDK+z7
7Blrzz/fZ+h4NYFHvKXaNJnf9wyCOjMRvgOIEk5oR2OKJ0ircrEXbY1+RymxbBtkHhjGQvs23bTc
YI1IZB/0CTVWzNvkJBRiiH6kHG8o+AJfavretmDquhHWAurHj7tiJjoEzGE6XEbC5C3LfNDAVXkr
vHZm1MT7jJodFcg9PPabU2IvoCmLHjgtZnlviImJMi/VllUpNZ8pzE1mLHsnIUikkNgmPetg3Cqe
HudGNUxakXkV8qWObI9NTbJFSV6uNlSwB9j/GfE3tmDvSYisiphgtzTxmhDC1baRJlEYUZlU+qL3
fNEHmyN4egxZXgQ2qod7fbC4RB6P9icmfoKkV/l8Zwgz86krBCoCptTNgHwtg9nGsb5Dgx5FURsU
YEKKQvFdk6qmT6CjePOxsJLrIElfue682b20AOwJipFIbAWOBFq3+U8ejTlVSWaNsnYrkGfitoKz
BUTm+yg1q0T3iFxKRR0z0p/+rCGhvOuFSJ0lhGIeaKxw0+gFYuA11dhmrpzw2gKmMkuQ63pkWTz1
oWfajHWlLvTaa8ms9/X7DB6qwy2iPJNkhECcHILEZrItdK22LLIvTuvWaZSdcnDVWBoO+PFQ9rLs
sLogdWjaLabzTDZlMUCO0+Nscmm05cy1ms/CAC+RiFhkbTPOBb5Wka7uAJ70UIYdqmLM1CrCoEUy
b3rP0dYSrXGSoOq6aVpIsDK9RjPK6ti8J8UZGg9hy5UiC2uiNc6+M3svXnWuhebRXAaFesBrET7B
mpjjQoFrmTnhtlwLlNoglVQgtsbBxAnBIfUWH2HXymvcFGir7An+3vftAMlS/NX65iIdaJdCM7v5
p60rm9Szo1P7aJ5jR8rYqhUEo8gGoEKPyhF5qNVciHCi8FHFh2WBhDPuIsz6enUKKKRZd2HdgOsU
1ShtnxxjJOhzTshk1s1IS157vsd823x4N6iXOE2YDnImPHKUNMVTHSrs3kJL6pDCqjyfCryga2s8
U7lp4wGYkk2WgdNKvm+A2Qi1It757PUzcRX0Ajx7SKoalUB7ujxRdmQOiV1Qr5e3Wm3sKs272Z0S
JkhwPYSEJgX3yPSOW/VkNB58xN6+DGzNIPItsrzD8gsvU6rCBpWZWl1BIGzL1AkFNpo1MQrN0HY7
OlO/HFlnLGlO/JZPiNRp7unxOu/2C43bdiVkDXkim/8rxob6P0HJkpJnKCHOtss8wI3CVREE3mfm
yDK1g0qMsPIN+BfYPYsLli/Gh0Hw0OKcR1fj/MuNqiSf/5AWWxR5LS6WnYOxP0+bY4uRJZs/resI
SjhAezTxJuXHVrqALb95CbTzVeFXw46l1ODnFXTBk825vdUDNTVwN9nqm9LWiotTtBGJWxLDJbjA
jtmqeN/I8bVxqXoBPvqrQfpX4kfONmx1StkDPr8YdOlJZrhoXE1X8uhN6L+SILi9xxA/ZZ/f6Mka
EwyWVpygm7AF/U4ReaJ21mcdV83eMYYl1VYTqp5ok3I9CP9Vhmep9i2gNmMFxUF6ibwR3clX3Lpb
oVpTYUfV2kz3besFcXfqXj8Lp7HoFQFCoFFj6jld+IWUTj1VCrhVo2ZoPmh5mjP/jlgkXfd3u4Hg
Xj3kS7MXCEN3eXWxI+v1K6biWPNur4m23u6nJ2yM3mVmGnK78L8c1CJbIOA9Yethl1JELBepmzkj
aELDCFr+KydedYeBWcZmBAbnyUkbPEaaKjY6VbSwlaUC52S/3DIfiduwTsqPHfZpAhPdQQMsbK/m
QdaTmFarlcRRb/PM8TRmt0Y3g/HJyUNU+76fOilvwWDYpcZmaQFT1xJ8LihVzVGvT4JlPZhz+nOw
SGD6Ldsb09rRiP824AaBhRrLqsq5/kwyYrK16LYId/cg14Nt+2qqx2TXtcL5TgYKwpykefNwiqIN
xkh0XMX4z0kuBgPL+y6ZqLxbgRXBz1ThQgsofENFLtaaUSCgiMdUYiG7ejQcR1rqEANsfTJu+Woj
e+2M7YoaAWPRx7uO5AEw9MvLlLHND8C4lEQIXOBzwW9mtj13ntslwCb2yt7AHEZ5u3giq0Y1qljj
FOgsMLVd8Lv5Oi1VFKP+g9yyjAFle0O+5C8ijsto5ZgUF6AUXG1Kh2/h0MQk2ivhEGUPy9cdXTdG
pqJ4hNYpDg8TdX9piOo/xRXVs9yLdaqEeNoEpTCraOVrGr+WL2vHnU+fdvSZUJLNg4730sVwbdLW
Wb6z4Pe4HBvSXt4tB8v0kUjQeFjqxEUDb3asz0RhgBHk91kANzmAucwytV5qsrNyQsrZjTHFKC1M
hUasLuBa0pyt36JlPPy+A1KA+qLWnoOqWM52vdAtb0xO5iRX0MytfNpN00j2t7DN1tumFk2T99zC
hxhtrtfa2Y8NHqK56tfYqaIO4RXkoUbgY8mjDt19HcGxt3Vmdul/curSBCgEZwyZz4pTZqPEo2dB
FOTqaW5T3Q2Cpg7DBUhBCHDZumsnm0T44wDC62r0JhV0ppJiLxQLylr+hdNxVo/2Xv1T2l90uR7J
+jvANDzqglv4sUu4g2S/xlUS0+8ZCKPr2K/JrxsKtzzlHTi7HECvMHBIcXViftJXkQ15PB6MNMIX
4b8TATcVpxV6CqaAaPQwJ7jmcn1MclxI5Z/l/BcXZIoG3GNJ0QFHWYwuf/E9rMfWvLdmu+DW5lL0
Mo6YLXsXM42fgqDwT7RoQ3Rw9Xe0e3+XJ60LjdYd9NwC1ll/N4NxKGoXqedVyjRBvXCj9c/FgRVp
nqRSIZJqET1n9Ik4b1O4THof8xgjFCV5WID7wZKo83tbeSdQ/EQPgQNGY3tFAE5+bu5dMmGgguyz
yWXzHL2bBRueU0iylF47cZtWT2sxNU/gIIj9nQD8DLGeCsWCC9THhgK9tuTuyKFXAQcFyFedD+Ue
JU+B7ZiPvAgxBnPOwCJ5UHyEYThQiZbp5WsAExuYRhrQRYcn+4k0k7myk9K+V/v+a3QAi4wPLUon
APkW/eBXoTzXmXw8xuwQMB/uuE9ye7JEqQSqOBwJ8dtQy8ihB8g+MHZb1CJJ+sTd8/2jtoW7JnwX
NKuOQYPEIPcDfU+/5vLW32Ngo6HKkR5Rk4hKD36b1AXV2h19kEnxecWTfUHorw4E8tiT1V9MdCfd
T690ULzlVP5q9+ja314+IBwuhmbsbZguOlnc7yK1rn0cx+2mSFaw03poaYTeJJU1RaWgrVTM9w3a
38t4z/UPDyd0y4dwAe4pKEQoM7VPrelK1oPZoz2T5zadNhL/VB1J+SsZmSi30FhHOSxDbDKKrMNl
UK7ahW2HsO0GOOCIEpxeBHUMg/8TemdrdgHaDviNysWzmyMNj5J1mIyTUejy2w1QVk+X5A+OwShn
NwNIoGPr53/ShvmuZJ3CUfOfCtkaStcZtejp+OaJC1zVeNkudO7reSaO9QOZJUtGdMjlFyWSjEED
lFAXLjh2oBtofdlu186lTSfrQsWfihg5d1R1zL11yvfPSHbnmqKh9oalrMDwuIYZ3cT0fYiApi8y
nzTjRU6INXYuhulcyKSfoz4MSqBKqNIMEA84YA3YNuMjnNbCD9i/kBxkLfkAMgaqbRiP4wyU5jGq
rGP9QKHPd1J8j0v3kupcZlYqCvp97tJO3ImNUx2JGV3xkTaNHINOR/JLPmwc0aglzhfqmiblss1H
zGaarOPvGU1s8Gjp+7ZXiFvD5shelkZTfe6IuoYy7yVEdphFagF5TPme8jky7RrrlrFzVs2PFjtY
v7Qw6K8GZtNIa8l2vcppNkoXILrxiQR8BFJDC5tICRJ9A4tTa93HhH/00si3X75U3uO9DEfYoOt5
p3tHX2BvSf1FaYVw7wDAEQJ93zZdNWYS7SflfO04FumkEdqvpgpSfshcJP4A27f/hkXvTbf6RPuB
/vR1vBt55hWFXKjZYRDXTVsNYP2vPHaSmoWhQwOFSaiIJX1/vEO6g61aM/hD6CHREUsUBKTIY/G2
f8rZtJWYHBF94E6gVBFbxjwi7Wue+B9t04GconFkeupd5aVu9pMvHjn4qL9ZwvNrtiKKDuqPf5e3
Gzb0poc3rBEvNmzeDADBVJIKKlybLwEH0Q6ZTetiW3nPDFy1Sv6RbTFLUV4NIXnxwiahGdRde9qv
ca0Hq63gS98VGQBrEu6Dd+vju1G9zDYH7Xk7O+cQJA3WQNRFf3qumVn78fl9LH1T2w2kI1iBd0SN
JJcjSAZLCykL6HCx4waO1kjj75jkC6WRush0wv4S2aZc282hGVSt6LnkIa6JXIod0FFNPuqqbd5F
Zd7Lc+TLnQgCXU6GLxN5T0vDIjM1cOI9bgnyxDnEcdO6ILE+Dup/xEnf26UX1BTs2CuDkBBxcsKb
Iusvut4NOptMmL4VzIO1qCEq20+RsPaDeJa1jfeWnCpDx/NNJgP9YTtNswbjhg+LbIfLzkolBjhW
yvf0dQj2v3m71n/VSwgvnWZ7y9Mqrilqz6KL2d3IO84T0xKloHiuRiJCx7vX2/eixNgwUzm6mute
th03A/ZGDkdxCKzQMiFdvGZuEXiPWPn8LUhj8SOsPlDc91sk+cZACzEDoL/8YLTEry+3RkV+qIaa
RoMSIbJgv3WkqxfJHESbFoWIN055LRUGrdTCi6dOweG9QmrqEYw9oUav36RI/VZFx/snkuM+jmPl
7f9epnFLorkVV3w31UxMryuQdQMAcJt8FXja9c6KV7wLmnxOO3nRlhge8MOr/0Vu37U9H5XTVCgR
ZJ2G+NXC2d2O+EfI9gV9hiW1m2uptLJJrAND3kRZOE4qpu7HpetcwHcFHa/VeS7qWe/5ot+aHUy7
LHyfRbIOfYWGXO4KvZtm1w6wjpun96rITH09FIWHvLA+vGRsG98UCFyByPDcZY0RtclGnwxHoTmE
neptmaulINcD7jHVx8VkCid2zxzt0K/XnB6m1Wk8dL4UcvqU+aF15cCXtTMPwaYW7p1StzBmQrsR
dBBGaMkk4nagBfSMltgOznHNtRKiYfrDX3PUU/dllzP2DFyvwk9AjvIycTn8AfD9fQVppuOfMV+x
rUIShAtKVo5L9cDJhQij5vXl8E61WsFgOoDUa1MifNOm0F2xU4TMAajOBJgdKjTUw+G7He5GaAnz
joDfTkSb0qy3Xsmr67g5qptAUosQkDCXMG8vLlJLIBwv/L56s9ZijhS/v79oKaejWVsFfOBy5lCZ
Mo/FnegOxNx4Q40I71cpxxFuSgjpgFeK2slTtI014P5fOq8AqrLZKL4FauOFc25OuRa/Ve4Ratrj
d4wBOzMPTLTyrmozH7O7BT3CdGJPztLiOgmO0qWiuq0l6433nbsRPtVknzc0Zmyo+pLp5Yzxc2Vs
eCRllV64TMD2aDvUWZvSMACojXUgQ5awIrEeYX6uAFf67Tq/TgC2/P9CuaHOoexkXEYTLr8yiGHC
TZf+A/DUJ6etviNO9xcDEVl+CAsQeKjkT9dzodyKfkfRrNaxJFFRoZQIt6efwZC72OX53LaNYvNg
mUXbMVEdX0cBViJuF4nh1ExVPX8qxQ7+Xa3vbrssfTxL+Ld2Gl2F65i7NtGrZsO4t+1cewPCbD8O
v68kO4fi8dzwTs6EzWtCEpJwtjG846SF0If0TzxChZ3rgN/Dn+7x21b/aWwp5m8BvjSElf78i//n
IB2FERLBWvSDXInryia6Yb3dSQd/zx/YycUsizyPGWBh6uQVqwEJ0oVLs2K3SQoCBw+kKljmdzjX
papzHPiPtRyLsLloAg8QiBRPXlCx8y66STUWypcl/9QImGrTzZfW8pgMA8wJDfdVSZv0Xq7Vp8M8
KaH3fpz//wlsXLE6JGPatW52S8B0fmwlVj18lazgKU04yoZwCVOiM6Y3Zs+IHVdFXZduRJIKBkdZ
Q9Z4UnKhSjKuNp4a9RqB088kwg0KhBUgPVzx2n5dXdQMNoWJnKStf8NKhWteR9GhgBSgYxHXEtOT
W1bF1vnlXmNmS5cnfNiUIZKrtAC2pf+3jmZWwpmdb6IQJjHE5k6YpWUd7agMQ0VI6RiBCQqjTBhQ
zbuvY6P6XyZtuGAZcNIBcc2GSerj7ffnW1vv+XXmhqwSmG7M1zoM3OfnZfW0eRv+LorFG/9rkJQs
9+v+LRoMqHPrjs2vthvO37VVhm/1z8tzxlLzWzn6FbGKtQmAtEJTNDTLYHwd+vNoOX5og+OYhbTw
WVq4exL261T7oEvxT56ykCIqevznb7ukBCm8Lp5aOUYyG5ZNDxwwJtI3bMtz/zdEeWJ7Ro9f6+rE
KIdBl4bwvlFeQn+Lc+ire6Ednd4E4VWb02rGcPDgjTAuHQMgn5yZ3hBEqKwzDt2s2A0/C+fx4ORK
KZH1KL+xaElycrOBJsFcVK5LW/gxY28B0pRVVmEBjD3fi7KHcfluX3+Cwgq3nR+LOLLMBOMrvnEB
+SkMNCET6DyjZ+lZjiJHaABDfTAX3hN2VhyhmXZz24KKVS+o9XIF4iUcyety+2GS3rlNjzxZLi7q
ucvtekaUybbHfWhDzbTAQ82Sw6tW+jI5NSu61yxUzGclxVX9xFthve3OXRvJTrYqEh2uZ2yJLOPX
yhyYkTpu9OwYX/IGDBIcN/dDDPq0Srqt8RoLI3wSaXAb6zbYV2pLN3oz3lwJ7AffT522iHI9vryb
GCVwCqDrH8sOFRZjDfH5/JbrI2MyvhNBFduvnIP9MtGrjaByq1ehGioiBfz8cg4/+vnylWKx9GQg
lE6fKnNew7x39Qq5yG3QjaSRjbltBo3tab2L0bgRKRFJOVh4ZBjy5LSNG1anIEpSPzlK5+OVNlTQ
eXfDOOkH0y+UxGJ14OYEqksFDafSKowAxkRqKNMK9CMnTfI0M5a58d5iDkG7bAbB7/y5Zm1hQpFA
PMg+LrS7H8OscrIJwsxY1dmU2Nc4Tc4gtwVUce0UdFW/eR7lQ1mUE1J5n4RD1uu1RDNLTrbIGx+8
AYFDN2INDCKyfXBcsWkv/48UqZk22osPFx4bRwhvxfV6qdfm8lRQmEKZ6G1ayMuxvK69agohVvdM
WuSj6pUz9fhJMjzBv0qQj/4sANgWkOWBcSXM39c7IdpNBU8o1ewlUltHk/rV7lMB1R7TS+zixXB8
uqjuc0hjMSyKXFQ6xtwjaCIh5FXBdKYICnh+igTmznnLjj6MNrse6o0os6hDUysrPmgIG2EtRQKu
hFBWpYWvYgrUkNHMIRKB5c8aY+kLq0i8oyfx9mHPMGJEonQncALo7rhq1HCVAtMF5IybNKZ1IX8Y
COUpE1eG2AstMCDjWxNEA5cqSA20eSa++3kSegopGZU9otKDEIN6wBBoEHPSK5zpmN2BXBYpAKR/
anuYVsB1VpdhJOJUD73QiDkUkuODUko345EagBDqfFY+CM1gNrPauZE5ojvaGtOGasUNHBU6JweS
fvOnRgj7YhTIrabrMJDGXb0m6EGU7stNfNwCmVyfJXl1nEQfX/MtXTr0tM8vcRp9FGIGhtwRSV75
3fPhnCJJRa9xAH8+KTeo4jeMZzjzvrvFOPadvdWssbyAEMn/5QtVJr+xeeaSlSCGuY9t7FtE3tUJ
gfXzO/KALw9HqK3X/giTHbQyHJnHh70GrwCFoH6KN2m3qAaw56bwL9Iv+dONL3yTKAjXrdmE3aVs
1lA/me7hz2z+1N2EkBHLPasRWtIKVI82riSeALYYvv+ESBMS7BOFAp+wqMqqHGsX9N6toz2Vweyr
4HGdD8Esvz1ZZAbr7Jpa2aodk8uTp7eG0MYjDRWUvw8jVgIysBmsmmJIZh2Ju7JX5trZFU4cQ9/P
rWs9AWJt4fkoWPIeV72IvQcan//dIkJoS8Hysvr3JP8VVx56Jd2NeiQ7+w2G4ndGRU61PIBhO4XT
l0Dxouv0sRVusptDOGzQT3KirGoidq3KDC5oYX+Saw9bR8c/jjgPgw7dWD6BW0c2XfRBDE6nGWcS
8y4kkz1vifzbVF3Yt1xwhSefQMonzDo/8jsEBMnK8XkMN3wLevMClB3bLKf9QSjAhghgpSABO0AY
FXwK5lVcFtoOAAlfwZK0KHIPRg+RBm3SCaNV+/4loGlXdGLWcfBXrVs5S6biDYKMtMYmPHnCRh1W
iM3QYkxesttdPYqLy4/dL0dj90xPItuju/P3PlPF7FRQNYTDo69Zv/Co2PaJucYCaUPtHU4aey2v
wai2sTti4WuiJecDoa2BFfeEsDczTF7YFhYh6q/JOIvu4zsQZ2e5oT2XAq7RJa4ImvUda4BUwxLa
nemu9v+4KF8yDi+hyXN1LJ/Rh4DHr/S0irY9fWKDgXCcDVdRkrwOQimIv3W5zpCoV3vsIpzvK5lt
5xZTF2cYGtMh8vjlK7bLK+guTY/yECqblyiTwGS+vkHuMJr47lsfOXysugTBnpvJKEyBWEwUPoc7
GatTqlzJ32yMLaF6AI+4anU7TAwMH7Ae0AOaSrZ/C+J87SUtgU/HgujT14Sdyj2oy7SBUy46Caul
l4T9odeOsfioUqmmVpsHcgAQzFcX/SgukRP7cUrF8nVRUMu6NHpUk54jZnjR6yJqaH71Yg+rMAQS
ywqbLdBFUSBYZfJBJ3nOM21eRUB2sV1yp7CszF95RHNVAY6GDNmefKQrk7WhPipqqJbsbhvOOcTz
wuoD3EYsaHvAAVdiEpKtLKF73uJkyZd3KMNlXbUt3bDEdW0+Tp3rdxCsf1dEhywUzSwQ2lzyXEb2
6HkSQZT0yxsgjP8jNKBHxyxvPt5utDKi4DcLux2/O+M+GZZbTrSH1CEZh2RMUM72KYoKsGjyqL+W
7qsd6c8Q26hgmMMe9BWU8r/DdEfXH2pShGn+qphRCgdCvZwwUHAqD7q9ALA0zVcb4sZ1i0VICr+i
z2oy/6BrAKP4bI5K3p7uE5YKUSVJDiWemneAQ8dckGsSpBeVy12zxe9DxYHzLU0iYtUSVgWRP4Vk
cep5e84lyeNweKk5DxzSPJjWSbw/eAW1kdL3ZsTf058odUd8Ey2QgRxAl4clf/LwuIwLcgiK11/2
Ub/c+5JVCzitLGGGWDcb75pCBdUz8+6wmBosTloYFguvDkXClTL1bSg5pFdRfipb5s64py6HEhPO
SsYY/Ygrz+mgw/psdynGRKnuqtF0dW9lIqzpft+SbWE8TEqx0G4EwMMnW5xDCZ56WuBud9f3gCGf
Wub40iMFGh9YplP6plIivtCm6h/flGOhH2itlICgoBOHmqOUznLb6HybE98XTgSgZyQbjMp849+0
1rtDM2asByWi708GqXK0M7nY6iZkYUxQK8RbYxJxTyev63AEuKGhVwM6VyNgnZClohtL4VIU1yYX
ynf/zbFp3kLwWVF2WoIgdXeYIPriPo0PrfChOS1JL4PPR9H07ReqVgkmI5tS4T5ErZ5BEeIsFRqV
wXVK+2NnJpQ7vF9HpS62lwLWUhDzhd77KrdyYveIhO7NvNoPfowwcjxonDgNNTckJzUTZBxtsn3v
s2+MIz1+EJ2lGXBolYR08Udwo971xmM/OJq46uA6RviC/eVzUE5XBWqdompHGItPYt/E/Qx39Pbh
s7zHNDPgc8JUgxEQ5YrMpKX3EroWlNxpawYgJKzRInDddgZMdbatr8go6BiL2je9+TIRwd3sAfgU
Ni70hmOwBbrFACwW3upa4fBB+vnuyZItV0lszQQ77jIMriAmVbd+qEZLDeuCN/7ACggRjr1FPsBM
l9LWJwMdebest+TJgqMqEHQNXrAbWIOk5EX58glKGbnm7DG/Z1ZPY1uIwAnm8bFsHalXOkLf294N
Hd3WGAzkzgexmmkdnW+OmAKfElcBMOxGjXMh/LF9EWtubeVuUU0PjVgjPC03WHakk6c0lXadIJ3u
U7EybRfnpr+pz0mK8d/avsWx2TXGz/Sq0SAqzDKrAG5Ru80hZn79tbl7ciCF4ENfz+pwuFriWSnV
874zNCk2WXUlI03Cx1BZQHs6JaKXvt84sF8N0TA8M0hS9bejxvlCta16oC6GxqK73LHR6eCc6Ho6
M8TDWekiXbFTt3gEY/elepKuTQVo5g+8Y2t2DtNibTa8XL0RWB0YTbJi7yHoTCnQZlv5Fzdo7RKk
j/+lWlp0+I2iCqZ5XhJDIW8+sy/gLSrZBIf7ALglSIXNnf0E0YAF+94W3qyD6pAEsoSwm8uuVMM2
JoY19Rbwnwm/K719qRczuI2rKjEkZ4wuDU0mxZjfW/x3wUlHwXfMqyNdV0zSZ/OV/yjk6078e/X+
t7iFJcyKDcri5Z2iYQFmQta4XNJi1qcW8Spcwb2OpFm/50fXjxX04cgyFQPEF+Hqx551NXACsIYh
puFQGuCpd5wd7YLBbh13CH2aBuGML9RoA9RW6flOvKtLCi5jONhn3abzX5GpbwlRN3koaHeowN+y
Z4dz6oXS1b7qx+42ZVEd1VdU0RRvXKrrs+8ptjFWL0Q1xo9fvWFzyFg71tKFO0xn2V8O13LFusLk
V0mN8sKTeIBcbAX52ald09uCDXUEVJXK4fTEJUJri3bZMLUe4qreLEINMnCJeTUIm2vCAh55dieH
Rqjw0bHDWpUYYORk21a/cyCzZeeMLZpLuwtCb1OZK0dDzV4FlhYfJxV5oclJpkVFMbvnf4gJhjTB
AT8GyGdlKPBqlnDkgBCy1MSdaE8/dsTWpUXRXQahuGq0YAr7R8EAhTHLberX97e1Nf3ej7rHK7te
g0SdpfO0d5tKiuIPoWQBJJuxYzLOCBzahJpsIzbk9x+ImS4krViWqIvh4jyKlycer/3fObgoOjbY
ROLUluWm1Xx51zmB5zA/U5Z77TLjaEXwxzqn8xXYhS417VGh8Ye9oCGzb/pmKz1oFzMZRVX9QgqQ
8HI/g3PMdyM/Igxmcou4l87ussrvPFQOX9nFL5nm4ctxNzdXtgPoq6ZR2YZE7cm8fRgbGtyyrXIw
lpOdbm5MCuh6notCe1qgAfngCZqEmSnACKb0GE9KZRrnbyER/S39bmAUPq5XPV5OGYDpwq0fW4mU
xU6FCYgIGkmKLgv/xcS6G/coV00KISmKc/IYgDc1IgPvtYXR03THiv2EM0neNuYefa+U++zPJirs
4w/OXYm/bvGMnybn9idIjIIsU9ojcH4ULror8rP82LzDKobI7DYFTnfXDM3KL9rBYvCBukCxyLoe
NgsVrhpUb4RhfcjpNvlnn3OLDhUHa75t5oxHXLCMBM4k+psMJNCo8nyppLDWDksiIhbYRAJq/tHh
s8jv+iSYqt4zU9gJdsJ2pGkqPwbJ7OZet9NfmuVTyUyWpICmnmO2Dd6ypAaVdcZ0wgaA0VuI7SxF
LZ57Ts8kVJUCd+OS6BhAljCzZowIcZataGnYN82imCBn/BxYk/VAqVaSCHSkINciaJhlfXPjlSMj
ZZeynoQJOC93y2Cz7303TUBCryCx16Kg61sgWY0eU9RJD3XcMfu1k0PZUgmm/BpB8QHWyx1VF/+V
NNTh7iEeXc6xQswFriR3s4rKZRus1saZ+Jl3kjuvNfJJ3epFBDWHEpA4eGGzV1Q+wh7Sa+nm2ToN
3Yfv888KeVsHzXAd+IVkZFfvA8wuowv2lsPPT0mo5ONBsGaBNRcVlA0coApW00Zl3tr5CdTSWPW3
FABMIbPux/QolAD91sB1Orspm9JubW5F5nXh6MhoUd5n7X1uwWVs0GYIAQYSTA6ssg7GQoKclWNA
wX9NtwmgC23S9SIogI62bCO2kpzRoj+HQ6fzX85SaPHcoPMHcm+ht6SqortKwzLmvKx3glujVCSs
5YAdY22F1cc6paF/611dEsvZTFDOjlPBS0HosoXozym5mFZyRaSZW5qABFibIzo+KDlQevxMDx0k
Za4MYKvHOMh7eB1EBFYdgvSuMQ7kunCtGFApcxB7rNB054UkKB1o7KzJczaynYkgtSOeZuHNJTfg
XiB40gAA00Fid62KW7+NuH68Nld8Dm5yVBlqVlI/O5I51PmQz+Y/nynkeSdVbPmNqz2l8lB10AVq
GY+ONhIwhziSekJZAHGkujiO/HE7qzl557/2YvncIYZwjO2lG8RKZZIg1eUg0pB3WyJIE08NlKmR
CMSw5w65iw4fvoUH01WDHqjaMTBs+GKo6QVpjoi9OnNlbgRo9Ahsosf9odEiy54y+m6Sb5rFB+n/
eJJz3HgXPq+VIggtIlVY04M9QxUABV13IthDi0aId5nSg5hgz2NwNw971580b/nYbzAikP9K7Y0C
JvBJ7o74/iGDSpgHbdUQy+jxfoq775SIsJmIilXYNGi9kcUHNnUhO+cQFOA9zpHvfDWGsRZgsuK9
BjueTKP0YFPGcewe9M572YYWTNaxwyJZYdc+IisOSgein9sJeHz7sbSBjyP4eoYgriFmtL5SId2E
Re7hdlgiBZ8KxsO78DnP3Rz2ZGB3T2U//tktAdqZYfLb+zu5MXWnfOukBkL9gIZ2xzianvwtmOeE
cJMqW8KiQ9Q02nlAlWriwDKuu/em4kDRVrD4Mizv8EqT2anFkk+6Is7JuDEBGQoG0figTE5hmKvU
0/vG6i45kIQFNCebq2gcQnDldlmDIgzsUpHeJxV6JGqqaVT36kDlJoR9RcmbZamSB3sUuBbA4uKM
rsJVHvooi8q5lDIgJbmxbowMWmsXww738zSRm0kXb0xe39JzUItPfzuTmWv/KpPHav/J+KCM2kNh
qsVsKUlCyYhdTIv8s0k9yjMmeo1qtwxDLl4ddWem6ON+2Gdt54O5HuBDBe7RhkGBxesXNMBvM00P
77Lg34MKJxTuh4Ce2WfNIDz3p+I3rqtlFXGaBEpDYNslvy05/x6z2kigigtmtFGTecmxKWG2PGXy
0VBd174lt/eN10KwcsqCLrfy2rm1a2Q2lRMOYe8DMM6vwKjrxUmSmoHhPuKjVFc7PrCRpGoygnJT
OGLbGuCKMj035/cYKT/wWpKvlnmzSU4B7x7H013g7BG95s4UN2iiubhvL0N6AttatqhXtIm+M1mV
sSrbVmHu8jkO8XeLSzlsAxqeX1TqKAdOWJUMoNHtyTNumvVIyuoWNq3T4+hy46zc1CuPV1rF3fcb
nt31+bwbXIXws9R0h9Gl0NvjxokXNAqGNjZDupb+t2ntxcAPsVMQstKMkCSVvEM0RQQbPgnOMyDB
laUU/AEyVsXK+8PQbgiQi4cnjdVXIQwfEu6YcLpaQ0rN3c7Qw0NfZl6XkwAerWD2zm/mYIWDvdRc
HO7YtW5mVT3P1o4grIe6rB33+8qwqfA4NXXODw2LWEZ9mEfbyvpbT1FOCvC6bCsQCnBJuQ/XcSGV
mu68PiTG9RDYeeSobJdk5M0SOh08WKv5ZrAuo5M4xVpdqlMk3pu8oTwPAIp9cMRPlZ+S5HF47bJv
If/HbrCFbc92P9rQRkxUu2bWk5tE7OFFi/WtkFu5kT/bo+W2+vp2klEoldvJkEMCvpYIeaeGLflB
7veJpXby2iCozvBroikahbJQW0FEkhd+eVsBm3PE8HSljeou7rI2ohmFEidmXo8+nQaAPl2P3nRB
3kgKtVTYH5YpETYdG30mm4/E0HA/OWfs+uivB3Up2HYr9tWLYZr++8LJwVnF1zlwOCek8ACk9jgf
UR6TMem7Nnotz+FJmwsVfxhgOYPClW9/NNCvxeEZBIVwL8UnGm3azUR6gxSVTi88OG2phx5E6T3D
4x8TlopBAHbcQp+zVQGWJaV4l8VsH6WzT1+hZ6dvuQ+tz5IZkOGxWASuEof33TdfP64r0zwMltTb
VzXeNQrrnMUa2TsvYNCC/IfPMBuCA75hAcq8G2PJy0DIhVMneVjOGUgpsqH/ZYAES7g1o+2F1NFR
sLx5AhRt9VXu7IMY/9B0QiCuC4pAyzohyC08vstPFLKn7tBjGjnoLm30pr4tA3GUC5OGZsyDRcX7
Yjlt2ANETDVmYWEADxNqT0aVHT98l1uZNTf1zXhq8KtqeOvf4NvedBM9p03xn3c5PYqmBKDU+Kcv
DZyToiP32CkfegdirRPWkLz0A75TGosS4/Ml8pdLf98C161rJ9WWoH5GTJxCeQyUn6FbnT/JEBVy
nvNU+qe7XQEXNOkBVZcb3SW3fVFxZ+Pq7ENdqzvG27d4ZuYPiwij2AjyTWvtG/aKZevPK6LTIx6r
5Y3poH8krIaFD5eeTxkH2lEJT5QJ8NC7pIdrHmXvPipaM6ZlRRHAokbpLra/Su1cwh86UoiXemXq
GQ78DIHiK2PQPgVD4LVV5n8XPeT+3FTNZd4RfYyVZsFxVMdQ+eQr3G/HRhoSsrLvRC4BqB9vJErg
88MwkDx0BDQ9vUQUoPy41+OSGmX/UflhEz0f58bKB8U2dQErA9DgMg5l2Njcn2sqgo7/OMC/afdm
dYR4VLRfti1ZvsBV9VkJrycKgNPRYrjNBCWBYEPZJqQoMcfgnhc5DRcz5Oc7tAbDgYN2nTf753Rs
ppBvdq48IRFuAc6F4XvLVyBnDcoziE3YZoxt/lBAB1Rp6IKaks7EO5uTJyRCKmyR+4ZALaHL1EVk
OqPcaRQkrW+PtTXOo/v1QXYSU/btETtX3/lMODBQ9g/I9cq2/3/xTVmCR3j+Juu+RE4ruy9+BuwF
4UB8FD/zQpnUn+zm/sPGcK+tvU2HK6lgdGQlTNscCQR3YE5lk5nfupCx1waH4GulqOM6D2pqi85X
n91dZ9I+EuLTh7BI27VrmZl9iM0RNa1O8F8ae3CZ2/YS4h8gSacSxDW//GL30JEeI4rxUWOOQ9SQ
FGeYvrbv+1/panaKhtxHCXjartSl43mSZvEWTVPRxvFYfrt2MdYOsikLJjEmGRNijqU1X99M92ov
mOI+++WkuoCy8ueAV0aV98zGWxXcAhMKWq1R3jHbaWLCOQtrZ8ZlI2t+NcDqrDQluLgSdw2U0XOr
Rzzla8ymMPP33/cgWx6qhpn1UObog+1lxOZBTSfitqv32Vp6NYYNJ8aMiHpH2tEsJOCrv+VyrQzj
msCVGlCPQYC6nkjiois3HhtHb056C8crf+iuoyx5lLky7ttrlsutCsvDb1NVBs0L5r/TPCB9grZ9
3EQtWI1Fct8yGP+NawXWcrMyrcnfQIHfKLz3IZ432765G+eVSaEOSnngMQ03gPakdyceDjhbhA5t
fJX1fmo6RVOO8JgVBf3TZsZglt2UP7EoybLD20VV1cKz3l8zlMgRZi3dBu+XXmCUjmYjzNPP5OTI
eeXTNm3LGFIN3DEt3CRyOi3mMEe8jfuev0Q17/GG7IuchaC/6fQT1e2StEdinHkiHXzH+0Os44eU
+11W2vffzTIiO0o0FSMq2XRIOr0M/G1Kp0dxX/ytIwo2cKejTPyZhu1BOPNtwwwiYik/zEzC5mld
+AkLMHeWbm/hUSqb+Cb8v40GbOtYwL20Y08Xac+dQkz8dE1Dw5myv9Cmozs033vw+ldVvK1KLMsV
UBM5zGp84nFOT0wWinql1LGIWv/meNh+IijWOdJ+05EdbqiChgVonkFIKiSmzak74n7WtSsRDVqS
DM+QisCSwe/ioK8xhl0EMZxp78lBxGfA5DggrDpE4jbpf1SW1IBpJgX1oR377py56qr52LDuFNj4
95CvuEwsTcL6rZ4x8D3+Sja67NeMsWcw0koh3+S9vhjDFOA0gtdYU9C+x8XHKvW3xIfopwplLN5S
prYOI5UPyXZslJUNSW+8cKVXettmWG47gz1Wvfoiiy/1KbTIGBvWTu1tHQBF96TF/lo6w2xSYwDy
dOoYE2xvuqEOp2IXFgFvsrDSHb5GnFt8eKrcn/q8E6r776S3jpRaxDu87cdsr9aJIE0ZV0ZoKKjf
M0q7LU2Lg6Z1goRSEFRtUPXz+bGMIgBp7yArYuYS4skDfaXsKF+yYBMM53obqkVUblBym+nQEcE+
K3k++AB+rzx+9es0up73MEnz6dkugtqwEC7Z/imd5ZM+EYSTesHQtTL0fjqtdO9xaBe2wWHd5VeU
D8dmmTTZbDyk+wfCWliAEwiL/4Oe+Z0MExHRf8DFUpeVERfjGA4rSAcIxjYtJfqGh1Ogwc6WI52R
u9B3klKSplKlNumFweT4az8cnTuxIc2XECqb9/qXLj+v3VrNuFhcMpX8fbDjBZhnYJE0ezq61YT8
DcyLGFvaL1kfp4R3P6M+tYh0YTekRKAIx75SLyZzCM31Kdvyh9e8snlVr8woffkuFN2Dqu2qao2R
uEFgfQXzDbG8foTMwv6u9mOJumYJNuy3E5WMn58Iuc3nXZUo8kvN8p84GBsfFNKzjq9ss792XqvF
dT51fGvfa7UxsEbFno6jzW7EjCCdMptemWgqRgUikFxsbajOB7nx/cxzUALuh3VUuKOinDV1x4y9
8blRGjXGtoOfmoIGg8ovZeoGC9s6KsdKRDrbe2szk5mrzUr/9gTq9LVs/0mznLwFMOHDwB9gBSNE
E3vjexlxvSeFKbpO1BDlKQtYcMvzyy/Vdk+KPsJbwsyxvOXusr8BIAVhIMaSktbKJMSraa8dsO+Q
zbB5Mu6/PTXp9eCDKoldJ/LZWCqtW8qsZ+AC45Yc6wNfdufnBB073Vom7egA+sK1UFJ8XNvrWqJM
J4GnFjYHgXKh7+ddCEY9Lo3ECnwdj5y4DdhbeBHgmKlXLM44wbUx1gUCdWypypnrSL0wghTpyQ6k
Hja/tIP8yceKYp8ga3pRQyevovVLqXOXUVQvGyuCjkOkr3w/+0b3G+epN6GkLbUNmZy2MX0gyPfQ
lk6mctflYN+bIdpGXH/v04UCyPHU2ihaEFjsu96IBGqOBHlvDqpVQSoaDD5QUidqBtQLmqz+IBbU
BbnocKuREJzfkcJXcKbSYcCde3Ro93QJdAD7rbIMFveZRaf+KsUh9PqbGqgTNQmqKzUKyl3OgeFU
IQllnQL1lTLSjp/TLJSyS5BQe8pv5LauSPBuL+4jIvVM79SVAuAVGjoOwpbODcdU7yikLz85s+YK
HhYB8AnBbyXtPonk9CVyymEVlBfs06Z3e5zecxrteZINzmy2tyiZJ0jePtDBe6tkm3MolJQHzfEC
6CLuM3MEcTGmaD4f3Zeccr3kAEAOuw+Dt0HNXE42Iyy4kUcf5+5gHWmwsuVIlyrCzqDas6wNxCB2
tYRudIpD1RtqlXvUKSBviz8p0++xtYfvQv6elLyvny3yKFxGZ0tBAe/z25xE3sld2FaO+dPPDULP
PlqG8pFUce6OOahSq1IONYv6MqSktLmOpuTJS6lu6o3sfj+YFH3v8WedmOwRMq8/prYa0C1jX+U4
grSRPblwVqXLcNYIb5J4j0b2iGwfBhNBhi+bc+B/bQXwgREyiJgvM2drPdi7imzwVSuyz2Foo1wY
mc4XzGCeGQDRHmjEGQCeZ7iH2MvopBP2TJN4sU/1UHz+zzKMm79/zuM78i/SNPxn6j9+f+cIbCDW
mo1hotKFy64O2Jegv4wxHiR8U7osEXW0nD3Lgr10ugIwpLL1ceAqaXfY836w0FgRdoRhdvz/LJ5p
o/IJTWuqLYfg4HGUgui5/yYq5mINuBWrd49K+VnyPbTovu9F+63UeuJxvQDoo5rZ7Vf5YNb63eWb
Ux+CxWxsLe6re9yTvuDLd7iVyn08VJ9lqxuVn77uon2osL540GzFttVArtpP7aPEHUPSVvyEV53C
GGOosalSh7KfTpl3g7OhpMFzFh4tjRu7NSI2HEHS8YPO0Z13d2bzMwgPVW+nQXYcF9/3/bCaaqhR
uQnSgrDJrZmhqASBf76TO23646tBBqtBkqkGDNY0YBjdBaj5f040DhwNnpQcwqAUgxMPtwqIcFg3
dXCWWEZSFDHnqgNpeGZawHnrVsy3IVPjzXoZASk+eal/oNGMhyxY4nbCTbdu7YdTmvE+JLh5zH6v
cemTbKfhG+UkydQbLZyB3EYRa8DpRA0GB+/ux9musL+qtaYDnU6N1fwctEyqiyYuBDtYjmZ0/ku3
0k1EkbHCHlG7ylPzZdnMGKzz8L96m6EiWtAA1m8dbPoJi28Qxh5eWezVBXN0+f8KMnleTLUZslSu
9gY3UKHWW6LPCJz253chPrOaV95ONm9zCH6lWfLzHc1w1r7JICuSf4UWOiDBhnUvXRnWT8i6EHEi
k9dcBv9HKhau0gpasAAGpytNSGEjLugrJWbYmut2JnaYhmruRHgjoI+7Yp8Qx5JyXQYsPMLvL5vo
y9tBoJQlMlYbPcAOs6FjWPF8eJvqI53m5/pnoEQlysyCdB+zazUdSXEM8xUbRbnC0EAuXNFcqb7t
FsFntVyUm2XElIpWsYR9RhyBk0s8qJP7wXV/CN9gLKiBinDqHCd61PG8FknyH/okf+hLIVjqKJjl
FcPgVGbWm9uhjJ27cVvGRFFJWOs2yrFFArTs4x6z0iT5bB0kQLA54NoAHWWYmjQNC8YOl/vQlwAA
QqFTDHkdPtiJfQGQxmPMWXk3JdnWd3Fm3RjCFA7h/p/0FpTNMVjWcKs8EqcFcurU+Dd74H18X1f9
sLiuC5BR5cc4PLYV/79f9gcYOOqFOfQwBS1ci2JtQr2pfpR/bavas9Xbv17ovjL09JpItXTZrdiv
RYGAHo4IE+WDindtWdsn2gzt3Wgdc+ORqtA+n/xpnbSkUi+DC6Yb6Oe+LMK+0mP9mrgYTrmgz/47
/aHwuiaoriwAgYmTnovR2lSheYVV8Vd7aTvWO7E+72N+Rv+xC4k+Jnd7gMOqdXFdZEQULtWeB6T2
/kobtqEiNqr5pxHdYS6cI3xr0xLbbmffKjLYYuhYu19YOSH35ufkZSAjdw+x0Ow9OqLctUXfsCne
96A1a+tfPtwsGx7esXbfB5xZh7vkuc8hWMzGa2XRnCzUMw8ScrffZJ+7xgcLohb0X/Y2BW4EHOcn
6jyIrKVuKMiuJ/iMK4UPaeeOoTOcnGmpDl59QgWBpoxjZidNmjz+1gt7xI+wWfiVvpIw7Q/M2rPe
JdR9lWA2nZI2tw4tHHRJx0S77AXjbrhHXPsR0+fsjumqcp06cfBSaMm0KW2yO+UtBfLaQroeiM1A
06VZyyZpCgVKvRWVwTKuVuj7cr5utQ6/apzdmqo6r+YFPWMOS6h9wWb2N0HVV5PUbiwOoYjBaf9H
MN2EgRt5iiaXSjiCNG8aPF7ylUMwIfL5nAYCTVLx47qHsRPsPI1807JfiA2ZxlCcDqaeyh0txFoG
fUnOR1tnvyESclnlIndYU7KB8RIVtGdWU3imSMkj5oDxmNU6R2ZvFVthywuFa8hGhmXVySuVX33u
5eV7d9MKk1jZuH+78hYxE7cdmm28LKJz0NCXOrk3eAUJcW+rFN4kb/Kpf1Zkvy3Gzly7rHVYRiBv
WnyyE97dwqnps8WsiYaxNkwBkcGDE7dFrG/QRXp04mjhqJgygIiOnopAIzJCtVKjbm+2Rr/pFhGb
LDZ24EcVQtNc4vuks4k+Wx2T2D+fgQcNmABOI+nKIFfl9XT990J7qD+0MFmNtYnY8OvbEnkdfXMx
SRDIFziZsIUvZvFNb6PUnNbetXtnsFSHJ6eJ3Mk8TAtaz/aDnkkBdYUn/ZupDxnS91iJwuuLfK2x
JI53XS9rzTPKHIcphdDmnb3cJWArWZCNvVRKesc7AdqUV7+vMVCHx+X9EtVoT0eZMduc+az5l0k/
ZrSbMIaMtUZA3GAKDlp51jBXuF+pADtZ4vPqRfcpODwLqzYInVb4l+LzCBlXbehfSnwei4FxmefY
9FrE0/fqRjVHYciJX6iwmSeBgscHZJNQBLZ2zd+KylFcaXK4Qhsk6cOaCm2bu439nT9l/ba39kEs
UBlOpRsNkGy8kx1Ae9H9rRt4+SX6WTNCpetiSBIzTgUQeADNNAqVrniqG52bmlRctq3a9J61PiWP
AmLS0M4MxHcyJh/TfA/9SwJY8J38Ifmf33fhuzKRZARtQElobQESfXWUxCRo5HS5SCQXTX4TxgJB
UNZdkinUq/S1iSVta5wF5AhUk4LlZQp4X+0EslDL9N+Ko7W60eN43C7MIJbrWzflk3AjqP2I3PNB
Qln4/JAd8e5P0A/X5/NgUXnnpM3BIMpGP32UAJ7woBV0k8UQmNOso5tWZUei1m3Bua6Hl1y3CVwc
5N1GmGXxtIpmyJfZxkpDShJV/FgcWEj7loUAA8PrEsdN91rIEpoQC1NYtFMCrmbexqWmpsM/eHey
TMzA1DIWFde09qAq/yp90DvrkXexd0VORmcoD92xOZZVLp7PPsNmgrYqXQJbfOyvnqy9HMFMyGzQ
OUIyGk+nv5RQbQHiWTxg5LmHB3Sof4k9SpY5CSKZvSTdtjJYXbnctJSzHz5jxn1cLeejOttRbdKO
sjIkyrRJ6l7p/F474DDe+e8tTu54kAbVXTEWGd+JV02udzFE+ntHzFLJR0hjg6/Xh3qb+axZn6yj
paZP3ldXzEI3yGOlH3by4pFU5zHgSPE6Kn8ucY9CjKLGHTCfNI5MAPBVjq7hEKY/1OHh0qkhIE8x
thbqpDPmfgm0e55p7hKk9i4oUClNWRGTwdICNIXLoBQuhVfuWiRvrIXvq08y3PUUEDyOfJbxNwi1
MPeY3eBNPiSp0N622NYs6oynzyIpIHE4yvpQicw/84Pd6yI8TCrNvTM8Pfzi981CO/0i9brGvab/
YKFmaycgLrd8okIlTHXf0k1WMIRo6eAJAnC4vwMQA50j0iBbO1hHIfTsfNCAYUXTuiqwoZoTqlA5
Ir8mBw5M74R54KDEiw+Esv+Ut2msKh3dirrrT/NUG/5/tZXUOuUjFrU73dpA7sIqJKr4qVk1A0lF
XGLMEIQlETrtyQ2Souif9loWykxeJ4ah1Ya9RgpCZyhizxG0VN1vEl5gfls9ZE7NUwwhjLmXsIWv
TRP8FPfKmWfORTV/e508B5zneIc0p4gA5rRh414iJNNEWeO68dqbEBBD9xnB+6zj4gtuUp41HWDb
POH+dtp8Cea0tF+Hw5+FhlKUH3ZDXZ+YaWA3NfkG7gTO/dI4aYgf8NRglQe1+DAetie4IvsmniB/
EDzM9z5UUSUGpkspl8rpbDoaKXGXSmMruGUregKsznvBJYRHKzZ71kC1CtEPW3BJFbRUCl1NXzND
qoBS+6Fwmjgl3Tkt2+KSfHBWxd3tjG7W3iIGrr4EjCP1nittgM5pKICnlAVl1KZkIKyKhDfzZs8b
RczhTZFQAHXO6GscvLf/nMtz+xS/sFC6pb7rYW5OKqk/NdO99TPzFdvJu161ZgSyaB/5GsUdtUpE
2CbLNaXkj2e2FlPFPf3IsFZDhy4EydyrQqODDSvbxlYF0Lxoi2HBWxnPsbDUJK0z/ZvMZ5uYRQLJ
rPjYjljAQi3vKULJ/zVW8nrnz91z10pp6PYOnshu4/TiaSdemmgz+0dlnirz07fre/7FJDli1neq
m80PSzAHb36F5lSJJqKRghaFqXtgZnqyqEdstb1KvSYVUJlqdzbGknZ5fEVG5k3SoaJRUtb6sQTy
B/L1qW6+T/vI1jlolNatV1UbuS6Jx+Bk2nGupurtIlSnY2bg/j+ZeyMSLlDtuo37R8oMXWrWIvJP
7/pCopQzLZD/hmBFEqqMFRrjtwBUhNgpzTS+gluXjTyEXwcT/v/Hweu6QFbOp87NZuqOj2eCe8Vn
gVAZhxM2PMQDTeyqZStEXsRPYE8vcHlR8Q9yi4gRp39rQ/qrtl7Oc1BXsePgqhwXJCGW4rTtnTFS
0Ko9HfKVzkMYcR1MsokxPVwQcnITFvIvZXSq2kEOLmIFioKYjmzsHJcd06IiqHkd7Te3KcT4u/TY
vEXYk2zqm1wahwKClAlHjWxu/kPyVJWJB/d1AVlR3pPiybt69nBnm76QX+HspmsBFXWA8bbggLli
iACaju5Qsm6yqBj6trNw7r19xcY0tcT1kJQXKPY/G665oARmo9P4W5ka/XhdSveCrqXJb5rLIzY4
R5RyYD+12NPdnPcqFo5LCdE5F3cmwh/M1L87iGyuWV6RBgzQKer3SELDKbcjEDWFBxM/2utRbRuB
CN/G/vmZANil2Mp3lHkT4fWAw6nhpHU6AbCHQeNwGon2g0KuCqwkrYOGdqw9pR5CsTJr4Fih+dlr
xeXtWHMJEKCODcYjFiXwK4753BTBwuaGDJH+nS1Ii+2OxgmpKdTef3v+EkaCaFbNBYzqozxAikSc
M+ARBnfxdEEd7lUKEz+IxSJVtIb92lyfILdjckD9P6BY45Jxhi7jXiPj1+Z3jX1yUJvWoxiC3Vuk
919hzzx+ZSfEGG1ccgJDN/ypvgLGQolvAX+BXImZ8luGB1ShbzSKfcArptLtwtynPfyE5BsCXJFh
vgk/Oc4Jpkv9YeiACthJ4olv6RtJNmluFdWtgodGcgrrUfCnk4KAh2En4PaRTP4OhsY74Uyv5arG
UNVO7kVjJLsSMQ1E7ZyRCbz1A0Trn73Keh34y2P38InrOt1zctpWTJ6CyLL9n2Ji8ythA983MYbU
SkNtXHc8CkhA/l2/Nt3o+U1S4aV1uNu3s3Zn8jIB9GxJ0SZy/lL4K4O/VCZWr7WCHpy6urZbJDYS
QVuOEZUTeD8qeFZld5PJ5gZZlJyjpkDsjE1z7h2IKeu2JC5z634a4vhGLgKUZ4iJyeRcc3UMFeXg
eboJpFjlHaq44zPJZsgjIllXaXCjPOQomZMT7tU5o8sSgtwLP+AX8iIwq3+Em/8TaSDwgHKl3L7Q
BWbuRL3gXllMyODW3C3VpPfdIUcfvd5TDsld/QFgKH46GRi9Kh57b8Mm/vB+HuaI72XNwfeH345D
SflUDav42/TCCM4LEf0uBALTU5hiE8DVrcoD31TLNfqKZOjGMKvG6KfUmvHRT/tjZnWiaTzZ9MI+
dBYKC6nP0bz31zDBdI27hEXt/aaLoA57cnxt5XQ0y2xIDb/eNDqLRMoGcaaC7Gv+L1/17CY/7elY
AT5EDUdu5/jWpV0WoH/ptXPVl1UDd8+4SNYyrTgRB2UGMijab0oil6703KkDY+LrutnAT0F3w2j9
hT6SK+OnCPrMoOV9whSdSBW7EedTu3z5BGMZii8aZIQny7z+fHYpPPRK2I5DL5oFbQ0DL7bWh1rk
GtOpjCjXqvxS9+Cr+YM9DCbm1XM5t7RWF5TuZBz9fcfjohpkIDnuHUUdDYY1XG35AoV0u4tBvQEc
W53GdTDpmdWBTbEjWWLXENLhurfhbJC5ZrQ8mEaoHoc6LZTAUibQYRc0H1Fs9Nzw4P1pL0QY0tXR
cbKBvxAlI6u356gb8bkrTb5gP5gDHViB8V72OLuo0RIkQULG74ByjT5Fxo9n1VOmTSBOaiWk/dmM
EMK49xAR441H/6ebhhNYDNK0ocy+3q/IdG0DPqy3PIpxN0vXJ1xanVayfbtJVeYhNrqNwYZXcvrp
JlkNHiLxFnT9S1pBXSndXuIacA0uTsBKPJbS6RmUpQweah+97GCkp+n5E4vKwgUi6MPo+kUfaAWn
uD23YMJY68d94UoblgPxU7FlastuiUmJD3tZ04rswXYidHFhrp7KZ7TqknjVmnKBFLLctUMWM91e
Qp8HSvQlMOOFo7ZNmcC3rbzgmOuviBFx5BSB7bCxekI2H8974/EMCJOAWKKK3fF47Ktzksk6L2Js
0c9iHahTzdzDz5WdJvtha6ukLmDoEK6gQe6lqVluKFJ/6WjAfZFAz8wmt/jxxyjvJifcN3/oy063
YdekmbvSuipl47VsJ+VPHsLzaqkysan3wKJ0kKJQJhS53t44VbQoYMNr9y/Tb2qNodMFlTP+u61f
D+u/OyEVqd5C8a/1BuQc9R8eDqwoGAmzgHqjq6aYJdv7HmeTz3xLHxYEbOL2tdlBkJUOeeTLI2D7
L13/x+yHiXsss25OB0fLKJViOC+CRVergVJsjxwRCemsbirRpYmqb8YPot4mqawtQgi5pY0dGzqw
rqFqEmsGy72hgHQlAJL4gbEUaHrCZ1CmoSArGQyYMz58bX8toz8e6IiBwfIJaZcSVppNSbF7mGFR
XhQzshdroi9owaGgnViNgD2/9Ur/7gOHnF0FOUuStK8ATamjgYxu5yM7EppbpJEeA79soQOKu2ac
cPyj9w3/21XWYXum8/QXErcj3nEQlNb+kv3k+CwSrLvmOeHYT4tjOUZlS+wfzeDuHUDZOVazl+Jw
YwS5KSDZdK3DZ4L2uHypmbfsR6B8gJnHIcVoUc1GtyZP8VvF3FW7K+Udp3Nw2hrTNtxCSOqoOGzo
hovP/ZsSn0T3m1ZDlWKQOCBM4GUN2OFnbtOiCOtXmFuKiq+DYG3LgZA0xwDjYfRRrwMWJ4XXG16l
FzwXtzHKydB08qBcQrZUsiRJZTiXu+xlyiFrPBYPYMAGApVK/JUqLrLB6/eRpvRKW12dF7jzQV67
0+00omGi2AmwZ8Lc69sZ0Mr+AQmsJGdmwCCzu559oSPsuKwMLnf9HP2LZ5ee5nMvibg0/Xxoj/Oc
3LHMAZlT5quCCEtPfDRFqRITEECJVeJ1O2Mynfd5rTdazgtmuBd3ePTrxTUoEW5cOR3WU6Z/x1V9
jH1GDGLSX60iLmODZPGqoKeTVNXim6KMmV2AxEweXnn34SaerZ6wq1O9DvSyKgs0TjQYiqlYmJVc
SafSrDAUDCS/EVXYCQKvzvAUomaVomO/JUMpqI4RcQ3dEvlKXWLrCkvGCbkwMxfUYRZQRIAQpr3V
Sh3szKyCo1aW8zpgMYhunaH9tkGbNAt5SMCDwxCCnQOdTsDMnjhu+kvQHibrBnZAze3mldKOsHNF
en8UViBmFzvd7wUntrMNcZ+h85eYEHtA6fXqQF+lmi0UDgL1JeGYLm212KdHTq/KottIpFbf2yBT
bFGs2+ibtxVbiqMW0MqBH1Lxa+qKtA9hNNEoYa2sUKXoi1O+6Itr69gKGVhWWr3a3myJfGaBDhRw
1lJWXbfUwlD5w9cr71dXWdSJyi5vfkeOvs/LE8OFv3AymI85UeuwZuKMBsdN6zdXD9ql5+CCKtH7
BQ28Lxx3ctrhG0K3Hss+YWgAsqAopiAafeyF1BCavkWCPZAGXKwMqAQOD4uARX1X1lkgFUxZ92e+
sa7jzeP2jZAvYSnuuupD7gTx89MtN23PS8Ma01cy3xltUU2oXIpebKOrBF8vpI4IzBXxvSXc1+BB
jJNO8wHz7njlhxU2HKWtWjIpfSUA490oBbIFBG+k402buN40vno/Zmz5a97p6VszqIO5nGx4c1n5
QqXmjNronPM41GZ1EFOZdPbGDbgE60J56YSg6gVvnHqazO0qCQX6rfu8PGhOpqQrAjDlC2/OSYa9
Il9YhBen23tKtYNkSdPtZXRT+rsRVEMYM3jzipCL3gI3Rl+ckSC2yfh3VtkG4m1wPrv4Ya3h7W9i
A2Zf+fdhiMfiOxJBqdU3y4v/wqXvKVMJ1a111Wuhd90/qAQBZSA+8gPCO6OpxpR1PvT3Ofb8RePV
OBklkZtkboz8YSvVdJVlaFuM0DVRQOUVskxJYMxSslKk8v5V/No/yY2xfjUzUG9bvaZDgO5Q8vAq
AkWaJYs+tSxPELvRuQt+MyPuo2jEK9MBQuS508ELjmn4oBNBfPRcPiQit7l+KgiTum3/B1iCj9mR
kX1m7kJeQE2WKxz9dl2kY+ZDjKyrzYEmZ8yRCRUQBgHwnmdI7RH79bP2wmsmj5lOi9n6kU6j/cqs
zMEBYwb35C0HQiq8vFzTrrj4vv8LH3/c9KCPVyLXs1HdvxpoDB80lRekGx7KOHsaD4b0Ez1+xLQA
riEn6i/gi6SAHeI07r59062wFF9l0Eb7n5MDpOabFJzoLcOgWoUMq+lSR383TZNqm7XjXeC4iGqe
9syy5gJdHVLr4/tPb6niPX7G+vpoeCX68Iw/H2CP9Sxapgfm/kz5NVP+A52vAtOCILJwIkMQ9rYk
oADv0KQnRzXd/C8pxeKrqmu7aS1ruNpwDzBo7dVh25O2SCvLuMfk14jtvPhewNZgcfsXzkGbaFGn
tuQ7AqpFtV5MgjgXSyvlruAwO1LIjyVZrxH5ImAybCSc6uSHJK1M+dfzOXlHTdmvU/hjuz0F3EpK
voUh3V6z6OpvIl8sb+xB3oyV96dw7gNn+gBGZkn3WNrocwd4B1KOqNcWObCxHGaDQMSAP2NGLaha
OtSHCRw+qtBLoTu1l63/OMdT7XPuBNBVZeh7X/abY6kz5vACfE2DF23vbHBk7TVbLOltgdid8Pl1
z7LU5CTt4218jyHFUGmO+g0IgNSIQ4+5+8OItVUcunpjy7UEn/Ey0M8O6WeK2ck1eG/dUZYk84Uy
b6q/tNQXyIPhofRewzWxiGOvvC3HTaYhsQlEUB+ij3EBeiBKDdS9E3DBTXa2MhF+Z4DaLR0wFmOv
Nog4I3oQIxnt7vjKITDT+LilyxAbdSOdQ3XKt0iszZu+3L8/uDnGwfNxViLKIFJKvt9Ubfid8eWO
16VgnYvugfH3a52LB+fvBjN1ktf2CUOFttDYxRgvb4M9E7wOn9UuQtaH4rlpXoxohVNpVs2bDG2e
iQz7M7rXYydNkbBDIN6uRDt4roTD4rPUNTE3gxuOxJdDbgP2uAgYkMjeEO9SZHWSCaFCNltT5wiv
L6v1yvP7N38kercqd1BEkFJaKSwZ9t/nyzE+VQByHdAfaGmiD5JE+zxD4jHER1jAd7NFPBqsJL0i
ZjSEASjPuYX2IwGFNxZ/1xjQEEOAPMHaZ4zppM5CtYx9EIHatPnOXKDaqe+SjGdwFVe4Svkce6oA
VtDEzlZnhLWTJFbxNUdRWLXzhPkyPjqO6VgDbDPlsbZiCBpCHG5cXptUkkE5kRfIRwdhD8xkmTeH
l3Z+2VySxVTYPMeXWmgkfTleW+B50NP6BN/caf4fLpVBwcECEAdvsL9ZDgECIPq+pFP3/jC733ry
gmdsBGMZK6AI6bFighiX6YqGZXoHQXOZ2wnxpkQnC33KZn6BjscXe5195JnbNpw0+1Mw8yPBIKrH
VGvQOQLqwyQCcpZBv3wuwrRjepoYFn1jOkP7gEjos24Neo4ipegghKTe9MVoZPK85on2l190V93q
bAUJSCSTRUnLUpezdIbty1qtB0zrt9hrFOs4wZviZrqG3Smp6PSvPiiL5RsS6ayJ/Ni4LXPyckVq
3RPOnSbqqwkDgtCRoxhvfNxgfIjnko29IN16wB1rpf3Wjd9jFh4tUOSmCTtvKNq0tlqTNyhaxRPM
xg9uU+1B4y7sq21WoTO4xsouRGExIkNndmARdhDeLh2yMUPAN+QxZHFEUHASUbhBIVvnyvDFH09i
xhG8EXnHvvWccTc3NavZKB8U1T3ZMPQVpPTRF60NPL7ra9urBKyaSdwA28FNWxU6WFPovkJ7PHu4
/6NAXegOHDSd3h/zM/oiHxMdR4RrU6p8nfkk0UmWvXSvy+L31I8IUKGxnqbrk2a7bgCRdDw4cZmc
fzZdt60+4jkg44ZPFYvtkz3ZnpNqqDSAqOkUb3xMMZW2O8NMeBxaU6Sr2834UFHP3RRG/e3D+iOb
o5/J+7Cd6bn/1ACewhFZBV0+bjsOHTWLvTgoYtZ4lLJPggBxN0pCgoxl59BILy4U/pF2RWczlhAg
OIOhX9LhYdL54gnnVtvCj5xtOhjfUECA7Gy2J9iDhbliUYBGJk4jDwIJpfbb2hsvZQa85gXdidy8
UhTRkEVK+0gKcmCQ4nWPzHEDgmJOKusHH4f3fWdheIREh27rmK/RJlZeN4TkdKQDM43E+u+u1Ysf
s0nQra20yLLURkEmDh9LrGLYQFAHmeup6AuU+yOZVz0BkMpOcoKn7ae+xyTgOeM69qgHLIH9ccv5
5BlnfQNqWR3Vw63atZyvbAdl040qODM0hE0hhq132G9hAIKWKPaVQJXdDWqkzj5tFuxtQifvZYZy
1Mpn03NDyYqObNdK4dJQbUTHfGmekEXF3Mzkat383nkLWZssx2F07K2irOoIV1Me4yFpdqJCQEj7
bqradBPnbomz0fuTlloxQtcaQEflU4cNposdPaluUtI+nEjo5qGBBOCBvbfm3l5/s+0YVMmUPEyy
HQccTjHeT5WJkRaDGRG60gNOKDHm9NdaxSSbPNRRdgZT025jLC6UOX/Nl0IbXKaGXs09BTtMoac1
iDz/ei8eykaXwVNF0jU/WADyXe/97fQqF6DtPVUJv6Z8AuXMo6q6Lg5Pdx7o9na8g3ukdGoGPvUJ
fBFRV6a9WYEX447dF2xYplxfkEhDZuqpAmCal32OVFvWkHXA7dnpjko7CFOSfDz4WV8sVai7LJgD
m7eIJwSdNMOPlO6avzxupWAVg582cWRwSe2xcX44LVXvFBd1h5Ub7R6WAFBMnBIVTmazwTtFIKGj
3aC7E6aoWarFtfS24DkxQD24cf6PRk9Um/B+EsvdkazX0sHDkYU/hYB0hQBkE9iAjt8kw+dgQoUY
fnKQMZycHlEZvPNQzfVQfNd2ccFCb8f07LkNY7c2GYICQPt/gvs8XRkDj/ps8nG0XZNhvkLsg38O
mgSDW170F8VCCgTUSapWX43nDe29tuo4BA6WkGAWs3tlF/f/cnu23rK4YlAIx7yrygZge5Ii+PEU
Pjg84wYsig92MVKy4tT2gmA+cNxiqmk9R0w29bzjjjxE6ntKO2nky2oxPQXO6en9ch9dx/dIhvd9
wm3gXH2erM17GjeRYR1JKip9uS+klZF7BpRot4T025BCm038q9w4te4WL/IV5AaYQJ4CtM8tx8Mu
LGgNCjxs5uvudB8eImFCUfhr9RkxIW76dkrWtd8WhDFd9UjCTTVfy5U2Su+jKv4U0/f8qsU2gP/o
UMQ9iCWLCJaLLX/CgUH2IVKg2TpjOaeYnvcGP+5+JnZLwP83hKaz5NXeQ92wqLk+gHwxYzl17nZv
giZgBJ7pUSZFaosYXEfHD+rwEGZGQmiYlG7eTkdeUs3eeWm0NTBvpuOcqRfkRJK5RUlMAQRjleQf
Jl4jtcHKwYskFmgm27hNsPn2eZZeCDj6h1x+KngV+6hdLnfxt01Botc7uEVxK5/qYc6p9q1h8gsp
tpDelrb8cv4NOCGlW5mW9i+A4O4eqsodRK1++982IN9eFwYnTZSsdaALDKBEY1mQIPQ4qiCx87Mu
K8Vx1W6iyioQ6O+gJkClM6PMH2POKlXxI2wkqYcFkwyjkvulinJJ1mjkxdyco4s1r4DoljfNUIZQ
JyyKz4bjiXyPWIKhRkFS+ws+KJnsri6Hoxo0sAJtiXvo7P2n6QBOlLbBXmjaVAQ5dClxFmNpKwRD
XCW3leGsfL8smMJs5moUCbL8NpRMUw1jivq36vHgBqQxm3n+gktyGrbJH7FEpDRjSrASpyquTNF6
LbJXnWsUKipe/IkZOPdKyYI2L8UyOv8H1W0G8CKt3TtG4R6JEINURW6DEwN8GsHgXlnJpTOpxpzI
U/7u5aU/+AENCOZbt34sPN88iBtI2Pxq6xHwnb+VYTp+gTBogaaqvRlZgVtoHESXLGSYZgiL/1m2
/EaLcUhX57FAWXneARyLrPoiAk5hhPWof1nXy3KY+S1wtmuo0uDUbBCqHo5J+3KNMFvU/5qon6Ex
eEpgd+/cyFpnck1kJ51CMt7bBYhFID5yy2lj0KAWz9B+0JAce6h8dDlTvmgVXC3N3AYWIL04qbY1
v8XJqiJeaiHZEIMFoFEE/KrLD5omQvPGD9qntURqNdzFOpiEcGw9eSNrSv+NipNlbse++HC3sP+x
wkubcR1u0gROHTNIbwH41+Z1Quo9QtkUyi37S7qiuY/nNJ2AboA9ryRKN/237et2cD3ai8esJaf4
4L9e3yVZWhefGsvoze+de/eOq4pdBNzzHP1QAgPw9rEz/cpezP+XLGrWHTlLdKJMYHARp0SJ4AlO
euCnbO3DtjkxT09JvUU7BHS0TKd+oMmcs/1b24d/6H79Sw3uLO0sU0hpMuMyJ+53qcy4am7X8pXx
/R0CqG/KJ+Bfp5yQlomIHFG5sa7yVgIibdbrsCsN3zPmvm9z17rJTzqBZfcvAFomPuXRnRpyG3rc
7RYwU7yCyzk7NqrEhim1XtqEvtTXGO7F+bSyoWdYJWTnzug7X2MnXqaMnhCEw3OZTB/btMdQVvsp
t+rHVa+TaOCyMiCdB9dA53Gb4AvaiJ2BRlQQMfH8ypwS3siFGGvmZzvXMQriMAKGuO2E6EJ/1zUR
PYUcLC53Vw/6hjGeJwCJdH4eaJyGPo2xUKew2s1WYSDvVin2pCHvX1sUiggds06/eByxVGWoFLyQ
l5ruXfe35fyG9pBSA4CKAjMWurpDETMd0IPivVIzMcQ+y97Q1sL/v12UIJL8B6bxWXXxU0XXx0dr
UJwZPvN0HO2RYyjNH8DUCryzynj53BLdSEC6fpKHQ3DKNNLo4E12+oLwFmSibomrjHbfkRrz4r0j
h1+pKD3uGIvaYNcX9xnyerh5+MOlZTCJRmLTRaeJsMjL5rMUgTBwZ0iPOXGgDTBgAktobBUYnP6r
0Wz0QbujoC8GUT1U4cX8e4RE5x2lpzlKuJoH7e9Bwsvo9+Ml4pevnwagG8kfn6XxJPSGeFQdDLtj
JTvE9KuxREI386A2inDYILULv/Mzvm4K/seZAxI7HCL5Wf2TDa0NekLpzS9Dtnoc2im4s7wEv/uy
N/1eN/C4TfNneKktIJ1xhktGhRu+H0a14Fg3hmP6dYgD6itg2S37Dw443RssS2J50ReRMhKTJ+WN
8Xw7wGs2XOTcq7n1h4McE/Qu34JkmLF2QVvfAMLVk9uXQnJk9E3Uqgvae1eWmXdhBItQ8e/P4TuJ
ZDHwtEOVkUGqRCwa/Kal3lmu5+jFvm/fINqhGXALgtNkY6HHolVp7T9ixhGtkcaOyI+eSKjCHgzx
exumRQxesLC58zxxZNcEsIc4nR72PnvQ6OZSS2dqXngqw0XYV8u6h3ID1pswnfNZu9B/vLUmVkI6
t5GmMEQkLfEQLPO9vlRxpbvq7MlcRIvpAguY0CDYij8bdXRPx+eJdFJBZQ9vqbKwOFECs4+bASG4
+UWeQsAvNGQ+1CxrNHdw7mv+SK12XOnRYPjOGThiX9ao2ZKl7JY3UhiKQFAdG51w0mFIU1UUUGxb
eRVk8yG5fS6E36/mPaguRzivg0fAkLM5LisyW/fGiRLc2eYK4Xo3s2OcPTp1Wr6A0akUkyYGuDX/
Kw5/vSv5YGeRQ4QFamWkY3Toeokbt1QO62s8sgKfh4XCgUYLhilZtnSjA8xFx0yKr/iGD8DoaQCs
9MVBE5hPMybOImoBxbEVJvwbITnwzOfbJQNeFnvNIldUIeUy2DDEIKOGLU753//wa208ysFsgNaz
OtoJBrWVlIMGoDDwflXPuchLSlYfGMfnKPCr+8J+yIrm6rP3BYg1x5yVTtC2lN++rDFVxd4trc3F
nD4f2gs3QUDs2R8DpIQP3zIoVj01qfyVvBlMv35sxJkiABt5eEPbbGIxhKXDRDT8mttoQBtawSSs
QeeFU52kY8WrN3A2PAWpSx7Z569X0OA4D4CHe0p11X6x9a3lYoN5uOOs4G7rNG+qOScDtE+JyJ9O
3aplRxotX1JMnLSI2bLfD9k4qg/VJCf6xPizlnKUFbuewJdp3MPwNzbcFkfDeK/hhcul7h0wDQsl
3xEg/WdUDxpdma+RB0Sp/t7clE8tMdWXq925NNez5wa7i+dUAHFdBsTh52u84sZ1UoDxKao/vhZo
yY7OMnqb8oWtULcsyjx+BuCIACu5nnwRXyoFg2nc+1wOpT4O7XMoXCF6SmPPsTJt56jUD4LOW2Zi
CT2XFH78LkE+WlQmOAH1wdrc/OxCz0QR4tUzTW9c0Uy73AGOY1eXyzDH0U1zEWLEoEEQdAYtlijd
z5Hc9CQztn+C573RbE1eVX2HO3yD3tvuLmHoqX+zNjKWUqkokCL+4CKG/eqzGwQ+x0utzGAJojp7
KBIIdfQG+TdoTLVTU0pN4oRJkIaLStuJ9mQzpR+6l1sOO88Z4vbPJ9hssBosx8Z/Q0mB92lKUnk3
yY/7VjTjVL43976EOLpp+E/vcDn++3j1KIgwov3XHXPjBy8G19h/oCAQEj1EmIavDVoGSpryfWZH
0lHuycY4ehAIVnABFXh1WQP/KinimZC0NtSbvhRAig+B/yVIJ1Z4Dn1PQEy3wcgG1gXysx6E6m77
pwnOA5ilTW/PCUqbVH3GAuFw5koaYXkp0v5ebnXc7queZuv/BIe1YZ5IOuss7reQHa5hK5qs3sOH
wLSqbypn9Mw6yQysYXb8R1gG4YecK8w8vM4J2o89olSlrgOXLAWz92yZS+Bp1hl30y+LMGGW95Th
r/OIfKeyPh98DL9DjReWMYaZjgYkIPwwOhtV4peO6S/lrqO5t3KRdcRE/7pyQjP32m5MookqlRns
W6jCWVszIlmwQ69ZBs8doqquioBPIQxo98bAjixnyI1KX6/Gq0LCN1nJ1KV1X57K+Ve24CsEhV/U
pbcdfKp5HUpMm6ADpWaehNu6rFORQIWVVYAeWleADgevq52JFOOzqVMVIzHpIoI1y7PVfzF+XMRM
jw0gukigfBTl8c4Chtao21SH2gft/+fAFrb+/Vw1YEh8gyZk1X9cjNU3C85ZYFzH+cpiS+HKNf/Z
lg2KKzBXBqttdDkTNWnuGMIhjfop2ntSOQeZjgvsYLnFoaMQU9iJNPMZ9Lz0lqmAMOkvSnBN8Y7S
NPyqyhNpust8swF8SQ7fiQ2qwgGGhxU0XuDKo+VIFNvf3FU56lkjyebtYND/EjOP4/3DcITt1P4w
/vk7+2efyEC2+FFKoSMLQcfW7iEVA60e+MMtXzQB2rHNRxON7jS5qbnkT8GZ5UInVZCNBvFGX2W3
IGzqKwWvHCUDyoarb79CraAr4Jhu5GXwwfU1+ylRzcx+4IMOmIMBzrVtgrxIhBT5O6+EyUgNhDCN
LwQSB3Gay9KEeUESauT8Osd7nJEfWl1ozThY5thmcJJ/qSV1HX4xEgLhtsDnNPPiBJm6p3OpiMTV
KkYDKBqXrn6DbWN/fTy362HGzizmW1K2BmiKpV56Y2Yq90PCTeUTGHHKGycgnIQiq+hdLM96Xo+a
MhihBOvfc7NPIJiUbYhoDQdqcwDOtr0+LKGRlJr8AZdmm0HJB3GsxJ9jELDNYJFPPfiWJyZvCFJj
YD12kZBBlVi0egSWyDE+cP8TD+M27aB7oYEG/mVw+OC3xlLCQv1Dk2ZfHH4/YgrhAZ26F1lrn/cm
JFI2BGRjs4+l8db3G2TREaz+CkOR7gBfWq675MiFeaxg8sBmpw54OhNimbDGA7Zhl5zheR0LRK+a
MXjwB5GrTkcDLu+9DTBVG+9eT4gaasWnUJS9O2/k0+3SSeIw7zWPRkStAIl/vIJ8NKihsBvx+H7h
9GTXtPIHP+ZIvO8bJAZAU8ZTU7F0KNxXIoRm0vQvHqCcOSchoTfiSewbDfWvvIeVKh/eKaZn+b7F
CQC/cQPwzoA8avK3/efNp9zNY3hedOy/sZV+XT9EmyqcomWmGFoir3WOSA0Ycx6zkGzZVoLql4lZ
AQb5UwFG3CZuCX8QPxskex4LVRfb73vw+ODn1RwiE3VQ0H5Rl8fvpri83rGUjBtEQEaGUjBPYs5S
uzBOU0X148PzMpTKnNrZ1xfe+Ag4YbBnt8OXHYkToGAi89sIyskdCJGy02v2ztsq0zE7J4uT0fVV
SdNF57eqxsdR2j4VNt1+EUnVNQYH41vITbBp2zF+ht8PzFasAD/xKHLqv4c5JJ4YVFvPwwZL2PlH
EwvjGCobVDSxySPE2WhWlnifn3YZBecxcwvv3jrLdBuFKHpuNhmOHDVW8HdKkzl4GvECAnSp43zj
CoEwbjuDfqTOovyMk3LgSOpRXsM4XeZ7p0u4RTtlyJ2/TrNtViUq+MCwyESbMohyokjTpO0Qy5GV
QVR4ja8vxVciNrngsTyKEvZ4qrkGPODqLXQS80Es+o/SV+HJaZiTmqHaFBRTyDbZZGGG5BEHHxqP
bvlGWSXrXSTh6srHw5NjsgEkyOuyVvgR29QrQzZdSwo3bKS0kwT4H95StE+sa4cl0MbgJzWLk7s5
rADfsffIDlf4R3+hRJKPu0WqvF87jKsAV9DPLOA5Q9R8F993kDFw2BukZ8CAFkBEHUEiCWj9DUtV
SoiiafUBOojWSO0hAe7/qE20BTHn8Lt9bpSc6vmmWNVeNWHUIyTQMJDNMVpWTaqDWEt/QG5v7nUT
8rmOsmc6zuq3Qscy/oUA3RMYwcbJQ12xj6Ji/09I8uMLrSpz0FMoQWRUrpPSdxqaOBelEPfOFlJI
DeKA8MoYwCQWaXqByFTB5C1EhlfhXFsIUMeXsRBgnV32m2L78Vkifwae3qTHgd3w403+gGDyWqLF
TpPSa4vCur2K5+DA57RTqir/r2U5q1TGSiJ0BeW7D9hNupbpKXA5N8Z7nensCQWIwRWenP6dlC7N
wZiLVjmJqHc9ftfxHTBGpaVtx9JRRupxS6NX0gJuycEaA/X92pwfSwxFtGu8YdEVyX++VJRYKHJf
iKfSnJQZxJZ7JJX6AhmlWaQaxdZ344R8iGta/Hp0OxyXhDxfxSR/1sqoBN0nmbABdNiJJ1j0Exd7
vTMj5u4d3G0rgnJprRK9QCc8rmNBlipv2JIQfVVsUTW+HjYokVltArLkaNdOS/4F8wKqF3MfzXeQ
5vp4zeeB7oYc4JG31CUxTyVCumQ2CDQRIQ0x5oMQ7AKFLehEy8bAO+JByiBsjAt7LjuszTxDpKKu
MwggtY+VibT0p0mQTXZ33Qyv4+jjZSbK305PmQWI+y3y7BuwtEg7gnI5tmLpxqw0Utn4NJz6KL1n
b8HbiVjqq2M8XMWbHvSpoEk7/nH0E28zRUBL08ZJB7mBv3UP04a+96VRDWowCN7QpUCtyxy8ewTz
Q5YqqTfuDecrG3R0tfcbz2z714ZDOB1y2hnyiFF0FhJ1tRlkxPbLTDybqG8GZ+1j+p0A7UILhYYk
hDzUUwssY/AcyMbsSbrI8HvyBtAi8YovFfQ7UnTpXtuIw4LZs+wL0WDv0mP9Dnc5Xd8zbLgtCBj8
7tZBQMV+gt9nVNzhybBOkjBczNAA1MnQeOBsCVxMfBkOC95q/ODW0jzBQyiwoei8/V6jJnnU14j4
tPtut2qoh7DqcB+RVwnFt1rRhRVYo94d1zbWN/egBA02oe/peW816CnCcxpKQa37SBlRVVW2JieE
P+qZ7lhvoSckvWjVzaDl+73Jk/r04fNKI6DEUHPTfePyWRiRSrUR0cVqxvSLeVBxk8LtqM+QQB1t
DHIUnfEd8HtYloRXQTUBfBjwcOHZcVuJQeWoKeyKRT7B7iD0rTxLEVlc3/XyEUZcwM5gZuP6Etut
bsIp4ccj+yU1TSGJAzFm/TMOfa43W8lv0duPgzfzB6v80U8ZdblrXnIEaYs+0XV5V5/yT9TY83ah
bjrtlnyMG6j+0yOsP8Agn44qJg1/SLMHogZGFDBY4aH5qNThPtawjHnc1iMQx1V9d8yLbJWfimfG
/XmCpiN1DvEcjB/fxV0CfSxgXGfkacFEEEDgr5HmGagm/TTlrFGi4d2IRNoAr4kqpbQlilx9Rle6
i3HiUG3zKSMek5RuIMflrIKOpzDQ1dng725hNDlBYiktvCWUVIDDPMP/G/OddQaRas9zA5t07j+W
CyyUXj4RTddnLSxJz0I1zocqlP6tT3WUa0hLt7egnH7gwycVIFFa1lOLOXo7IRX0utiS5VJNT1QB
a8QwTf0Q5daFWR9JZEu6+uQR52o3hLg+fsLM6yApy++R2DFfYMm9FzjOCEZ71Xlo916YY2yafOjS
IYl46Z2ENqIG4Lm31MS2ibRHQNjfJ+mmT1HEdmr+BFkAEmuRbDWHBONIDwSS+UTbuANx8RyikXKo
T0ZB5iCkTXY7SzWyLehTagtcJvqscDAFaD7v6kTUu+Ps2oMoDSchkPKAR/mLtcNC67FYaqOzs7Lu
gr8pT7QWgx6M4eSyNgvONtb/YjpMfF6Ep7hPa7tH1tJXUSqbVUdqbSOwKIH1fGSW/LvvaCxkvDfo
2rq1NXh0Hcys3CctmcTJJnZxvY0BeYs33UyGBnM417QnhgxNyW5y/opgp7/ps3JjleHJTfN1cDNM
W0P8GSNYdBHQ2gzcZQT6X6FPLgXQ4fjhuXa9pmAyFUm+wuf+I2s565c+jQUMtOTF7sj9smf3P6Ko
um0YLHAipiHH54HEkLNmC3XqY+uwbv1IohssvzrkgRdN3/ZLFe3E1xFmXffqaEoq5ULPB4TqcqWx
cu7HDwMM+ljNelmOIYiezYsnUfRmbigZCip4+/Tt7Xgy/+GRrquVwuR7WlOVOz2eXXrkdmxlokOu
EzPf+O85tSNtFY809Wwv0PclTQsThOozK1vCfhB1dpz0ek39ZWu216v/sH3MjoQ6udZyCZCDyzfD
G70yo9szcrzYGGwGeMfVsOa5bZuX7iR4V9ctl6EECyJ5H6LJ/KX6jhPcHXWgu72cf3JkquBJXP4i
ybk2a9wDhjori37f9GBlybh7h1TebZFqhfmd3zvDbfDSoy9/SWfQyUkXIzUll1fzTxCymPkCCOuw
Io9fGJ+rq4K95ILvzCTp91pNpg4OOQdcoi9Vf6sMVPxiHVtymhq7t5o2WNF3Kvp//V4CJ5SWQcoL
+sN/W1gVjRs3KO+s24ZZRqJmcZafX/7XeTvdecckEAu0rgXT/6iYxhrsOWLF4v58UMU2VoyoT7u3
+5I4DKt4qI3Q9mJe0HN40BBa6CWffAz+uGUkJTSnoyrVdaoo5DJD3ldv2Et6Mv/IPLidewCULZO9
8RaRPZvw0MF+KwRNeSOcmsGxWPM1sAm5QgrLnT8qpfx7zk5X986YEdTNzS0FlbmhvX15Q+RZbe50
ozFf1i2aNW45abafr39J+/cD7Hh6SpEvHW5No4YQPHbHySdOKLa2fNDedpCj8kFyO29YaSDQK35P
opcgH8wDAUGtuuUWlLo5uSlewczZBbMm1qRsDdflV9J5K0k6UN7z3T4tHLudkl4fN5MWoYxkALEC
z4lRV983YUodaNdVnVbGDVppCp8Umqr7e1sUaTcVLmd7Qwx1g9geT0VlPJ6lyw6kySzXIvUGftaB
EowqrLyL5iRgAfgWAhkd84CpnoVSc37bWQuQm6m9rgiDvlBzC9PE5TnhWrk8YolsCHNr+gfuu/bU
k4uhNhMJW6kUlj9hBSLTbAHTm52/uHsOcEIN4w8YVhgXrMML+6ZRfvFnqKLqOmi2NLpo6OcFk4EF
YdQZ86SqMpyTwmBAtbo+r0p8Afo6xDXvNHyaTrW62Nyg9Lw+S9by5RCS888k8FwM+Oj5jJsoshVv
oaB9bYdYTC1+rGqOYNGU7i+o22YLcBGnGgj62FJjSqA8L06X1H6/dSrEqGffCs0UdeG2bXA7U5i1
Y+mdd6e8qYX8/42WEKPMKZU4ZYo1559KRBwk4fz0tJ2OmnK/Za94RaBrsObhzGUj635MLt7vUabt
0Bg4ZJyR2hBrmPbHbYNSRMHzQ1cS9ttRM1G2m7nNOu3QmWLR+R2k9ZmFOq9nhUMm1ThgbvDgC7f/
dPKw3JgxZury851Jd4P3KRKL5i22STFq4nA+apxr3GGYbNfPjlBeAyt3KEO6JUZ9eMtO908KDxfU
/9Or4dd9WWa4UipDJ1uDyeXPt12xFiOjQbh4ZqQipERi/jPICM+qq0ud0keAAoutkRq2HaiFaa5N
5GivlSBJUFQ3RAtKaNCRN2IScQIcjVTReTnbCzRRIwbJU7nzFCEb/Jed8tdq95qeflPq6/ETTCv+
lX7lPAWdK0eLu5zFysgovP/Req034d9z8QLDxOQLUYDHf6MxYmbrRZjOE7EK6cxFxWUWteFEw9zE
/rXlbLZpKmzHQYV1Z5cmDvpQ4fWbTTyntv5Y6EmMpNsrQ7sF22WtmwRtbSZgoXNkkB8YQMxEI9KN
9FFUE9H4UQ2t4BgnL9dpQnaDUn/dAV0FHUmxHm7QMkCcRabW4XGTVQ2Tlynd4PRvznyJs6kTp24o
FqHp4jgiQkYmj9nPZMIc9M+ACM8NQUxhHApqoLMcFmXs7bVEu9OMciwr5tjvadJkCX+hL2TpbcEc
PECkQVOLJVeSmdPnpvPwC/JDjNj0WDWMDxKdjftLdLrgTPBgG4O/L4xHG/o+f8+9rtwje1nytzmx
tqSmbf7gkTpXi82wV2RtKshKPMFvib0kVW8r0QmNYphqOlBx8DEOBfTI0bwb//jBF8GFhKgF3dva
9XOHaHO0at/qORd8gMAB9bboSjvyg1gWIbgtLfVVB3JmgOrH2JEfcfnt/vSKPr7m7ecuQo8rlYia
N0tKqHIyDHGYTZqPr75wId3wiG0p5oaivonz7vBvj2EpKSohtZ/dGW56GcErhHrQngnduaP4S/tx
TVMYXY4cgT1gH10B52zUT3WH3Ds5C9o6GCR5nuwFb2ggOA/rPVsykaZLOw1yhFfZqE4J141xmTp5
GYGsgFetGpoxFSc6Kge2Bn8yqHR1zry5ZebjuCydAfK1tGiZYseSrJLqG96yoPegM9Qbi89qIlWI
E92mT6SIBcvbpcgppZ2wAEAELtgf9jqL2W5xklplM8RKQJafvcWIEqNxOBrBwEeKZwES9h96MWNQ
fFsUHk312hI6tEB9WFqApnsNY6de6GFSRnzp3i671WhbUf7HgIy4dxA0AVlCPbMm2C6jFba91zqw
RMPbveEgOUl5PQ3F9ge6XB19j2RiSrNe2CzvVc4syFKWPVoAeaMF0HLcPxyq8wPc/Nd+jrifTQSy
Om4CABERCOld9TM7JWiMHx1CRI9gXP1uHa//4/AcqrXLLt0L5DSPKPpLJYQyIWN9BQsL9bXQtYsP
bx8XzP9XLQcDQOrzOPwocOxmw5WPgQcPiQ1AYe6pEL7LtdF8kuwJAMMrMI/EUeWW1pSKtwcwllJC
6oSIH43jUme2hYdUakvhSj5f4puHz/DXbqdCmrU0oqTYUKai8ME88Oxv59AxNx0g3PL4V23tcqcP
8pPTMuArA9XmYh2fqiadf6dGzAmFHlu/FPBbgZc/s+gZ+kQvK3BwnYPY5xkNs0eeW91uFRhee25X
Pi2LuAv8unyt4rnBhqZv1VjBRiyGxWauGGbVUoM1/acn2+yawtFJCj7sy6WALwEf2g7QskwQkkhI
3ko/Lh61OND82fFXpXS/CzWIzoVXYZYeIwEtNI2TMimRRmBMi3Ht9swIkx1DxmsXxN357tH1In0+
PTOREgXdZpZn8QDnM74KJ9caaWkVkAfwpS0DS3Ea3zBbDkfR9hWL6nejGmMdsRsQaMYbBqq4iA6C
BiIHYrbUhNNQ39SGITpS9Sa9xGk5VIQrSZB/C+z6nTHBgma841ZNL2fkCLMIWVdwbPp3U2UTrlh6
P3Bve6VzgGgml6pJhFY5E2jNPZJkdoTid8PKKhdGfTrqWNAR4OaUzM1OyeBeVV+MML4CRws59N/X
xc0iUVweuzpWClMaitQj72qdXx6AcRBoJAXmNGqeW7fDntvO1hKg7Xi05y04DN7nKVrFSH96mN6Q
aLr39dcogP2c2Rt5oAm2tgHY2bpcbVz7FBmZZBaC6LYxuWjviHMRYqThTXhz5M4pamwoJAhsFjAa
aWLWYTRhyAWHKho2DszNpyy0LjdoKS9TjJrIUXpDq+abDBf2tQ7JDrqspVo4haWCIJ5s/byyCTzn
JKO9/AC7tknuiL54nCIiMNz4fS+BxSXfg9QFDFLlZrQTtPFdWD0l1hj5LMfJe+Q60Lio1/05/b1i
bV+B2rQCT3U4KwvFnzPfZqDHkOtSMdu/sJ5D301VvDZ2fjTjzcBxlPbWEZhWOFKTl+zVAvhiHQWb
WRft7d5aiFnuU+bXIoYCpqs+fGHY2KUOfuUKRvHVwz0pn7NSiG/bO3BiET4H6JYc/4YmJPlNW+wr
rBELKBpL8vUrzMIHltZ+av4J8NvwaKHYBgk7UgI3vUiitEkFDZUmeevEIuegak+9em+4yb5mC+iM
4LursM/DQKeC5xd0ZmpX3iEy4WaI+8FFFPKKHugDjQrOSIlsVu/yQBVzUbEdhrGmpfntTSxYPa2b
8Zsjv0PXbA0n5k1NMv4pJ6ovGVu8wm2uQLZzS4c0LujmEer8FrlNkYS4WRBxs2IyvdakdauXfhai
px+ahMuXocOMJz+kX5xsfflHvFW47m0nQ6s+HFB/k5uMG90gegEsePp7LoUKE/oXq7dBE3ihUS8V
HsDkJ5c1LVh88XMCmnMfFJNeW2lUL818Wh2bpxkyyStS2YbAWMyXx60XcERs0qlLNXJdb4StwX0H
SB1prB+wUeQfeedeG23xWl7Nbl5N4oBCK6MObaPvUQsKzRET9bYU+92NhPNIHETD01ARidbb2WqQ
ZSZu8zG+DuWjtXMG/RuU5cjJsXheX9cZC60tS3d4d+OliLxqh0TLn95dAD3bdXJfkeuVzn+JzaEK
axZ1sahcGXpSPS0N2EOBGahbdeLN4zY+dWFJqbF59rdf/sbpHcNOZDgKSFQ95mJgMWONPtKgKhQ9
5jzY/iV+UI68bWr7NtxGs+nfloSd0z9xNZ+uvOovaGBJ9xouYv6WELrC+jgCDCRZTBpNAQRZ7wk/
MmJ5MvU5ql/z9ItfTBjJzymfpD8Ru/u68skYJgG4LzD/O+ubiPolQ0fXh+1vJmQ27BDKmW1BkV+v
ErRE1yZ1dRbXjkCKJJ+QTN/xj+fhV1WJMdYEztEQZRwRy3rrTBNugZ0iH2tiHwz7cY2qB6i+FZ8l
wuIwvvSn4qm9RI3UbASPVu0Qrqv/Pr6qyw9mJKHuliiIzHpJOomSnafMRunqUhc/IFgX67aKZHZb
rr0mOlabPmG9ohLo23gbt2XMuljSX9/UDEENG90jJ7O8YMNu/6s440IW1yzt9/dRgqu7Ls9PNUKH
hKhvyFTtukNTsYQqmxwRDTG8h7YP02mKQB1AtPGf0nBQZcr37cUswYlWVzwXbeTVg7gq2Vu7Dfzi
wozqREDcq0G2y8AQ0aqnNO4tUnz94eilrOxhfc/ysPwCtif3dAeez+C0g4M9UJzN1lN4kaY1IXh/
r/wMVHKbZMKgcYqwrhlUPWGTc19GWgKjR/S42/qDunqvLetyih681ISS9p/nYLbNoKJv7fDBXcM3
eH9LbHYiS5nQtiH4KQtY6MT2z+bPYmmQ49v236/wp4rKQ9ecfJEu9aK2NjuggctDoYEdIIJf77x4
OtlOcZOv7N6ZMAyXG6T7+94z8nSjkoTawb7oUKhYejNtihgUmFL7kMwl+aEw/Ci92xFsjwTpLpzk
XZM9uqBBtq+FsE/OkgpCp9eqMTjdSbxyKVwlv/39RrNx2pO9yxOvc7mMP/R4J6mcdXwpFRfAOxWe
+jY4hAIsC24F9sU7S8/L7IbgVrbuAFv7UOZBbUPMpIfZlr+2OkSoS78Io0BLGI0ieNLgk8ujqTyT
3yPBlrRq39BCwY9oaVhpOt+cjEZTdNspelZf4Ou7DHi1X1A6CO0utflhOS1nPSOvMncF/Z4C2xEM
OJeAbgpx1ZijusAMRglJsVqw1lO0cnMLttszLr+CokUXOvsY56HffMYlNGpS2hXHvKYjtrv5nb2C
DYTiCHpuhJCqap9nM/VDrKal4BKC7A99jlwAGtACbcAAQnXnW3Ja1a5bAk8jMJRrZhRwlRtBFpfd
JaEJVt2vZyxDMNybMgrKxw7fA1NTDHT+I5MazM6ye6LxG9NL0l622WfZn080Iwn8AlSXiGF4OKTW
L5HlerCUNwKpfpfiRA8r3LLtnuSjZhRL9DbQy1Of37BBH33ELtfXisopjAWX600TO1oB6CNFhkWc
3vqAaNzyR5NheWdLkbc4MX7SD3Rhqb8zs9pOTHhh+FBPQthHcYQsKmHdWJAGNGIjPG6KU/PjOVzh
zJent/7mIqYqyMSqwhDx8lrjKKCeT9MAW4WZ9n4zZpe5JBz6IvzQP595FayQwVg4kcX2tW1vB8D5
gh4aZR7iwJEUYnp1qJwJfxSmWO8WU64e+9Wkmu4q1bOTvo/MJGin32x4SGa/+eoLY9bl10UodehB
QJWdkCYAOSxwkebZQwOJluZc1fzog1SPtAOAuBXQ1CH7Si5B0+Ej7kLcgHMFwDL8AYeObFHV5mrZ
9aga72MKBNR5p0O31QWlZSYxNb/Li9VYlX97cPBJGn83jsDJiRua1Ji3MQJXnRMAfZtaXPsGypoj
zGIA9pE5eDx4KIZs47EscP2Sm1A/PYF/eUDrsS6eqKk8QLzNPdXuJtNUJkZejGhTR8yqRgWk8yCy
X4ATgjQKOKGxlLOkRYqF1sWi+TvbHuDnbePU6RGu4aOpJDVXry8iiwQXuEshOaLl+pd02aSjbb5M
WLIjSju2TuD/P7wy+3yHtUQe5iTfybY4sSW0MYXhs3kgH/jxYVm8+d/c3vWD5Goqd2IECO0jhol8
HeiXaNt1wdZLqnmUgQiE60gJG5nvO1O5Ot+CzLiT1GyhfMxKSdsY2U5cFAsJgPjRzfgeej/Zk2Gn
UQDNXH5ZOvQaPn5q2DhQ0+nlWkKzKMxev0ImOIdUsI5YCEjOLZLGo7BBx+C/stldbXE2NRapl554
W1ut+f5YpMt9VsbDZ5VWE2DTZdP9NKIDcqDHljQHGEqEZjMYWA1xplqYFg56xR1/9EyIhUmSfwTk
oaw2z7McsS7gi9+H5gB/eAUn7dVbnCAXWP+xllJlUJU3vcXagqT2dVGArYN4avBtlNLBp+EK1Ldx
X2SIoRxN+SbpmKOElrD/wx9U+vQsWmJqxmmeGkgEm1zNGBGMHkn+8/uLw9oid0PAsJRyFSqckujj
q5lrL/6ckWg5uIK/1wRd8NrqR2/8T/vSAjBfIrsD3ot9nCqCkDpw3tExK1FC5Xbf33xWwfHDK/UK
iD3tFwQC4Rwt9OJ2RiLlK9l/AdDLlsdVpvuu5esdLHjGxi/SKtjjflVxb4AjlDWfoCyNYpBKmkgg
btxzw0E/o/U14rds4vyE+eLdCGoCjLpMv+e4Djzp1+S61hRhtHsOyiKfJmPNv+kxH5gd09N0g7z3
ttFfsBdMxE2IVKtNZKWN9H02pou3ErGOyUDydWQEUGHuxM0nRVFnPt4tCYKOgm+KfApVVF8wIup2
21QGx/bu7ge0pdtaW77sMBTp0WN/QYPuhZxmAnivPy4HZ7pUyU5IlvuvUAAbTP82Y8OOHBdqEH+i
zUKFWj3nV0YpaAIuDIetnO1vYgL53HhX703KdyLfJQDuLIQbsEiXuFxBgMApH+DEGcdC4/JBjgzc
NDCufepxZ9ijqsBFl+TJibC6xR5GCRKruYdzJ8G6EUMHK+21iIvntya0SuwLEOW+AxnEkrmeXhg9
K1bLmOojfIlqABBGd3mWqDvObrypGfMHWZYm2RiGlJx580BvCpWzr6nVDucINuivBLy+xakYA/QD
TIML5KymwQJAT7erG7uoZ/FHkbXSWwlQKEG1qHfKuYWo+ib+ltBS3HbsZznNEUyMbYlMm1uiC6n0
Dd0HrjpBBYK6qzzyslOgnrtazMFDy6etjWEbvRm803oepHWzDYao7INodEEaBIbN84u5eS6tswWQ
sGMpd5A/cdEjpIl17YNQ559twgjwjZVkqu/N8nT2e9y551QE7CGyd0CHHZx+Jh/lM54EtplzdMm/
oP2zLOsaV+8u0RlNler92IpXp5h8PZtnUSOJWNtbCYKVEb7PjQAlO1dg3wCSxV38ecvuxUM7bjS4
LwYawZDgm9wWIu3BmkoOG3zm/EPOMHJYbGQNuXB2VKs3JcBYGb2sbhuVkZ1+WlCKchPdLcu5r7NF
5SYR8SuozSEcvlxOO4EdfVQ6Ifm7scnHKUy1Wn7+8SXwZ2p2TslQo12fgaR1GTgIekexQ0aaH0OA
2PzXiZOfLI/OVrPccdAgN8jHs7ZQpdIKKqOtL3MZZEiFaGzDA8Z0HHC4F/0TdwsFBhVhNdFSptZz
s03FX8u9lGKtkCVUl8rVrKPCqCwq5eXZYVHAJ+M0y2sYu2zAI785SBL4XtpewjfvQtKgB/esMFtL
Xg1C75hOtt2o6kb/LnDxaTIfLmXMz7gwFNZkaHcfOmITC1aIsncF+meQTu16NuMtWfXril+6SI7k
0pWOUXPCHBiCvJ4UeX+8EiLc3F9OtAuofwTYTWjnK/xr2M7pe2uWE3CD7j6kl102H3NnHo7Ahy1R
OX61UjZ3iYVO2gRDXhznPwQf+JnGll9usU2JMk7g6ia7v1m7wZ3h4Ug33BJD/dsXLv3uFV5z8i8I
uoBoCAXrkU4vEL+kW4J/swakFIgou0IrQheyqk+wAD8ZvBSo1j1cvJRh0BnIlbCNnanSECmWlzKc
u+bw02ZcXRh9CTSoqk0M8lny5lS7tKy76WY2cUNCnpv8gNei2QvJHmWNf2GigWpxLEL9bQ2Inlrz
RgI/zbjU6qy+xPT2MQDPDSjzvAcAmeKHRRataQa0pDNDZj+/RhlKv+ZjWR+XUbuDSUB8g0ZeSMxL
KBp8ucEYgmT6Y8tegyyr6LPqkG4zyw25/UOyTzvJRdhPhL3RvG1S4GR0US/Lbbt/cBvZ6A0Wm+P+
R9XDXM04jvpVmsAPIwTdwuT/qe0kUCcdKeJcLjhV+lrcFx8uDHkgjRFAZQ3bo48Wo9nDq/BQfFFp
grIoZUVKaDyeBkTKPtLjcW/XD6o84mosre7FuUQdFeGjzyxcEeAN/yKmm9UPAwcByX55IhYrEuXs
UrxEMwiWiz7jo6u8RrsTxbf3NvtzN4H+Id/eDpgNXngLN06dsOh35qEgH3ZzBlmpIYfMJlObRxrm
35Q/kEzIjdFDoLWjywEuS76GdvW1oEe6hbaVhfjKtbjWw17hJO6DuYYpBiGlYdsGAyZBQB5HUhra
AqfbaBQd0IkSx4z/BazOoOhTlm2SjxZgHg5G3c3jIpA7t1fiX/DEZFX17WDJy7TVv/Js6FpQHMNp
y/KM4Ve9u/IwUHi7ZoksKgQIwPd3GDir4vFVbbAzpX4P3eIAyUMKrF7qqqMPvWBOofb1KDc0a4lo
PyRolemKtw22jbPr6QUxliB9n85fZYFd0t1yl5srY5tNCy4oPMCUwEupzH0UYkLOVEJ5HyddcOw5
1WhRRJ3ePghimNx6/FpEsNTA6NolfJN7J9JlBtDMbD6fZ5gK0awZlHTL3WD0hVug7BeHlS+qlv5f
wlR2VYFqDBtWk6aGDvf8iZjfXSO65tz0N3BZikP36V5mcJRrkYpSMpUc/YjU0+A1YmYEfVXPy2+o
XNyPJBpn/j5hjB3w2QzgHpqx+ATBm2tJrM0oEJLU4W8NALfabc4SQ4ZsayMhNR+e8qI+CQRIKfAN
BdE+5pHN83X71J4dFkldiu1UDG6GdRv7yBfa6e8hsOapuDsRbbkwky1H5L870bv+qEt4F0CmkCwX
6ertv7Vak5Jz26N/TOxnZlt0yMoBKNYk2SWukWiF09wMe7KeaF2jBWG/bgNmxA9HZWdKXUWJdKgA
XwugRCVxCqm1XdJVMBz3Rw0ZI0psyZMMQmBOHfT9fNPbHUS/gvU4ECtbBCgRbBaVjSQeUrwCK3kr
9BBV8sLxI9uoFWYzVPu1cV8V+JSzdI0uPDK6C0R2eJRqHy1LsEfbu8NKX2oItoR3rVbFmFO7VycZ
AOZQJNcTYHuDtYgFwCBvUaRZNy5+N77zn3oQlpixPeWm75JoXTDvZe9SY78d8GvJQ/VVocdFY90n
GhyH/I7tJHZtNLwqFwGK87N60RnUsV3QMENsiswaJGnHqOxa3mQS+iix1Q5Jm3Rnvk/OJr+WFt5O
OM8IohpB4mo57FtWplzczxDRJsuosL7bk3yMkrSFxBam83FnsrQ1Bmyo8XOVQ54pMotWGMkiC5LE
zlIJzGafHau1mdRXH4OVVWfPI5hJyToOJzhHaRgh/VjylartDKS+y5dJUJ3/+iejQYK7/DpmAtcW
wNaAS7ocW0pvvbdSYr+WImc7Ql1HFKABOqCV9EHh8FwIP0o5Kr1kwLtjjec0vF+wM3GzqV2m4ZXF
36AcAVsc+6qyGBFB7osPzh1TCnddtAnkkeUoaM62jVxOkixq/EexbZ+DUmhc10ZLMgLFiAEkN2xY
ljogEaqPjS+Qlh9EJzkLwyEKT7tUOOk16guM68HrbdjKeaDHMoAMYJNpP6TjMrKwXf0Pfe1+vawT
csqFW5FVgt5ghBzby8E865C+Dy1eBIdmcWrNW0Gk9Nscu84yHs8rwOs3aSBC2h62wJnQY/h9an/B
9jaLugGkfHig2BG6vWsI9tsAL+nKD5k6iuF8UkXvslsye4c2ABAJq43UzsJFnLvVroA7hXNMSTf2
iIpgVkh9fpGx0tY+y97xc4g7X8Yc40c3/LH7x/mCPh9Q38D3k7Ncw2ZMhQuBmqPJdBwoLRDaVGEZ
QMVfu84pCsYXwgp9KqyaV01F8oz5ovfuC1/WH4GHKZCtSZ6lisUsfneRX2Ei1JhQO6F6clKq8DBe
DfwxfiSvfdPopWsbhdtZrS/jf15E5xYU5h9qKgi99GSCJvruxhU7lBXt6/CIMa1yY8Nbi9DC7u9e
1rnV97j6TCnZivLLdY9KPfT0zBbpSDt+zuAjO28L6ij1NMWOpdq5vT8xHMThUxt1QcXqjT2+gGiJ
DiRPnrgf85DF9l+ZFAfx5AOVdVqPsn9ahLt9N7SNclRV66RsxFjUbbdAbcEsFPCFTPwXPwhCSrMv
w+PDN9X63866um+JGJ4ULaq7BYxCe1huPHjWsXSk54M+Xb8LRe8PowI5aWWK0F1qm4+A6A1CQcSV
nta7U+IeVE84Rvjr6yRLRii/IHDacm35ob8Ino2ZAgQPaQHzHYQuW+nHaJzcMRmGTyvQ6MAmovtl
IgSdZopQx3yEGuvrLnu21iqmbMzsRRQ0LpOS9sStdQS+dP426YLm9X6yhHu+bSgMCg4Yx0pV8dzI
ZY7miRPllQ9C7wpONnd6rlo/hhWrzoY/r7mN+hFwp3SO2golNN/957xOBMRZwd8Dl56IqRke4+az
5MLrS+vEXY/VWDG6/ly6OfwsPh//8dCMwYWsWB7/hK0XHvwoziG+S5DVXAIXAFEP5LZEn4SYi5Jc
nKo2aDRPBQU+nzeDeHtdI4ouaC6EAwhKQ9sLJdDDdeIY6GitwKFPljSN8ZZp2L6kzN6hd1oFljnm
nSIH3MnlilobTzFKmSKE0CKMADHMQWiwYZzwhq1hFIPASwMrmzquTcJxco6o39B9ik1NKB0lhHAD
dgynsG72+ClM5uCxiVI0bDTvhIWj2l1QaPwMnZDTOYbB7pJWqij3HrMPUGuQqXL5IG3+nKv26tZ2
ypSpoHyCQ49Rii848um3o6KWETL5lPXA33RZU96ODNLOVE02gKbq7gcqO5G6KiG+9DfB63lgvE2y
NSEBA0jL2XoywW7khThG3/uE+/icUZP3XzejFPSfXlsJKaGzgxjvnLd6g1IHsbPTF7eyd36x5jn3
okqoYMNaV7Hu/b9xhnReBbcnwHq8n7oPm9EwQdb9IdBBNCqCCzcb0e11iCEf8JaY2lFzikhZ1LGm
00xyNMv4r8QJAVRhSmFS+Ww1w6Ma6OlgWZY4NdaKFnZbO6eyBhpJ+MzmRHTuae7LudSMgJkQ3aqD
jhcNni+Gw6C1MePq1NxA3a0/7pg0gmeTzbJyM47VDqf469F5TEeQF/j6uFplsm9hzxNXsD2Ah5qv
Cw9GHCoL+WeKUsy1I3q0vuV9OzLfuJRAM7SogpVutd/FaLi4KeHFvwz7gt4mZst7YP86K2XoxW2D
sQy0IuGVUshbNWNcPBO/YS9AZaxf3+2ygUSYUqfzSb/da93+M63A8cMizPobQPbnlV+0DKUYD6uY
AuH03n0KxUjx5sSXNHLNleb5AfUUfM7YY149401SSgO5mLjf3cPBBjaN6X1dKlcxrl6fAJKuqxq7
WqZWd1mJMP1e62eySHMwmsG00mJ4WaXBkBEHGZz4602sT4LJmjGouFHiG9KyB39tOn1SfHyQY4hx
GjXrws5z13nQi6pc0tCy8qitH762wVUML2oWJHe5P2IYV5Cv5qoZKe+Q2Mo53TOBKrzx0r+wwUb7
d7ty4NvnTwvoheH1Q/6/5JnnYY6FWrzDVtQ6WFVEHFzgSy+JTgDXFFZX6o2CvVYBUhzdBkJ5aIDy
CTHE5HvoUlJHXOpMqEJlgDD4HwcwYAbvqm5Vgu7udm6ZuZxw6usMi5exdLk/lQ45n3an7o9NxTus
06d6pyRsEo912rSVCqd3261tFAEDuOFknzInK+nCZ/tjXkxb+kP6IAdEv0gYVeNnqev9TMFFOx8g
J2Pphkg0jXUapaxVe+cQNu92B7pMnGag5YyKKLUjcbaLcLqqwuwwv133jX+ztOHam2cnpxOS846q
Tlbo31dWs12IJ2Wx0KrdJ8CJUdDzE2486m6QhTVIsf7Gc+scdwhwWh87MWVdGVaM8Ib75Ww5007Z
VLJMwyTSWirRvlJ4BM5bpwPxx0ahAMjwJU8t9r0yPBz387Xfa3UtjIzntHekqR3274kxhxuDH978
O5Mjp1KZyo2VN51lhK2lO0Vy2FsstssBTK5BTYBgPpWZL7ZOlkn7m3nJnHzgnRwfckfj1r4CYEGG
6ivyVfXyE2wdEePGa0nS8xov8sDqPgTcX63wnYTVilI+P0irudQQJwJAeItxfmgnvOcJ8ZhoM7Ir
vBMagtqVhVaLdVjLDpKTdloANcowk+oF+55KrkeX8kCnHwJ41fuR8++okpceHJ+n5lxWqovJ0RQS
4+WZjwqf9Wqbx3HWeI52t0Ry0OIZljJ5pBb6L5E5s7RLgMcTLaBdTWUCKV77/HSRuCSkIhuZfFDt
/Uro6a0koXSjkan8+4Yjdlz61Him4Efe1uD7iYzbg1bxS0PTvg2DymrEBTuM+iXzkGNxrTWBJoVt
U+2ja/FErzw8Npi/+jdhWiRuwQKimqBuJAYaiMNONfJuTeO+yg1iRMl+GzDSSNzaIkRudLblFJvi
DnA20GIzKo/foTBX36CvaTFTdCNbWaPIWsf8mE7O7gl8uBpBuzV6yH5ZdOHYOmSNpBRj8HpugFLc
JNlnvM9atSD3FJ61v2eEOeB0r8QBarxz8y2ENi+wp2uYfSFn+mtzdE9mhQqmaalVgxdDu31Uo//c
pZ4g6mnHmuHmB4yWoDiYe1mTJcG4JwqJOhDPGonImdcOsPbHxKxn+zah2v2qJLU1OKyi7g5oS8pT
s7QiaXopASpi+3roQXOlNCdfFQssSZ7/+ixwJyu+Y16oUDxlyjYvOeHYaCSREUIAVMH/IjAWxt7w
P49PF3j82oa8Jm6LhKAODUzPQF29NhEMTBcvbBNVx8ElkAHQQB7fUiIx1WhgGmKD1x9K9VahRcD5
QSkMRquaK1fEAbm91/DzuIMWnQIJRnczemJWfFxWZd5ZZStEO3gx/tLh8ndX+b80tKGdvlDb/NL3
HbW9tSiSAizPpeoRnJTUGTUzsvNrlTZqjRM78aIFJZXLIw5ss0Pbd1kOZl8Bsmh8tUrGS4Cdix+j
MIEvZVVID+RDr7XibL6iQwy9i9MpBH691nVZMfNVDaa+bXW0SD7q4L0x3V9+L0vwsjpqH0H5HZRd
CeV0C4fPR1ujgxYp8n4vpSzchsubH+hWp99Zm2U4LrVCHqQyq5SyETtm/P2LfjH5sQNKJaiPUoOY
eZhjU6vL1bk9/wJ71OJRxz4kgNl2XOYLKq7jSNkZCut0dXnJc6yYfk+NWHbDSMsUoDNoB0nlkNrf
kG6fYhJr58qz1k93QfA6zQpiMm9LTYrfK1bwXB1ViIcOXxRLeihMKJ5jAm5Xnbk92xPLLkndujgv
H3KelOfXpgzYdtmYC7psgnuZjbsltkdlJYUuAvvDRqncTSQureHmTJgbtms1Zwx9oYiGRF08iZlS
1K7MnTV0aAmez6Vfgt6XzPYD6w5qhk7aSrStL4rsWA5UtPIoUeyEo8TDxBJ7au4feA7Ll9OLT0Fj
WgL8rkyrDukL3AbHaAcN+tBaw9AuqQK1xeSjPxt9KJ/ucuWmauTXh6WWJw169Hl7HqCSSp/1lTzI
4kusN905yuYD4jiBdTJHlMwvFjEiTEV/1PH3PiMlsRPXU/DSBTD1Pup3eWdfDJX21hLlA1Scw39q
FUmc5A0I22IqjuiL1uQS05ucE89kllqmj2m5HAtrX0XlsgpOVpE7B+QxmBxfkUbRQFjkTeHCYWdg
tdUHKaVcdbTmrUbPzIboEkzUK1F7h67HhGlH1oqLTm7cSpDZsD8fj9Yx1/iTZpmmgPPXqaTaYiPR
fBbwkdMReW2sTRF+dpUWR6dbQmzVx/0LpSGMeR/zJmvkx6ftwy5QbdFGeHZjJvF9s7gcZ+avqP0K
o/b80l3Jc5fYMDuvzUCFIbLXluJ44H3MDdhx9IsqLjx+qXJDkZzAxW5hgWBHkkQdZTzsbyA6NOXb
hu3GNNnE9oGukXZ7bz5bMOjpic8gozu2dA07MRzoy5yQZsdtjQ6XS2DDYXFFX+seVmMejeW4BZG/
9dAiDKbodZ9Q96EEW1qKM9Larkdqdap9dvuqsYrF22DMMcq1+bV+y5bsBL/VC2IQ9mHXb4ulvqjv
gGeMI7xWMJz2N/EIDCBZedMPmXaLPO8REl7F1O8bZhszG1zWRDAmXVWGybz+E4uXjtSe3ZDRoHIq
8fA97yyjLlcNIiOdkDtHYXCC4JrdedxI6EP9cVL3Kl9ucQsKLOh8+ZVCuC+6eFP7wqc5iez4YQxH
ntTMEN+te4c5cxi0WPWCbY+rs52KPZLDXsYGSSNHXPrUsvy6kPEpJKMRH6J4o4CBuH8cwwb/ckiQ
fR9/UXbh5G5rsLleSvrX1+QwAU7wDfk+vScYY8FznPYobYogjI/c4F5LQnlsPkWywuYfN+GNsoXl
HpdyVn+NJbc7cH4gT7DX6+oxQeTPImiqU8PNZdoCIqsx9d8+uUDyPFaH4j5j8lA8vJOYJdV+AVwh
F93YYwNdE1gUz6ElHpvHnuHY2+I3BnVpEMDXILB6J2nsH0PAuNXoyKHGpriUsCeBOC+gWrm9CHnu
GJ2KJHWnhDAd/3fv+uwUIG5YIMctwy62hsbWINCoKwnRfQPtYBiNKoLhsbg6kII6xQ6OBCIiRqU0
pw5z9zHSLs/ppmvXKJcU0XmRKJivXscFlJVGcGB5E6iI6qThDpjjnUrSXaE4qk6WQmlkFI3qbK2O
WPNaHyLw27TtTFvFd0DkqZxV1ln0OqxFOzdrR3vBE8IFk0IhjP0IG6i403T59m2XLiA1oZxhGMNd
B61JiAGze37G0jOC9kEbBmQ/v/ekH5l/wbuWpBxz4kcsYXn0jT76pX9W800aQBdrpnuyaAupIpyM
MzuNiNjjvWg78/hx/XC51p/Qp/YIrhojWBT9DeUx2IVI77qE+PviegEtfa2T7jZ2LB7c7eTqz7ZY
CqTtEvRadJhoJjDu9LEfI43MEIoQ/b5BY2loJIl3L+ZUDnuomrRDH8+RCcMaGMaZqSRj2kuVPZb6
wEUIjmpq54Cg3k6wJbiHIr9EN/MpThGvhCqsT4wNS8Ke6hgZTpg9W82p/djmHJ4dnAvZk1GHwHrh
bGMthseF/de3ekc+R5lkIXISmgx6aZfJn0P78JAZNhafmEuzdaCojPQtQTBxgrnAKiIeNY3Eh4FA
LdXpMR9/lcBX/ZMtvu5/P8jdW3D0uxyPlsMv3pNmGZTj9vNESvpuO1Dnf8Fkba/hXl7rzohm2/lw
TL/sIcr5LTW9SimraKkkbT2SpJBDbOLhQw+4zlRhGYifPRwq+6R/PDO9HotRfxLdzKrM5hrisdyJ
EBE+OGF3azzJKo9unnbz85FTCctm4mFcbwQLRnNZNq1tHKQtsV0epT2aogkhrTm1iFNXo7BgEg/f
CPj5eAB9pJydV3z5iKAKGV3IbD69JwKmbq16uAk5NSUnVMSnbSec3YC3g5ylUvSKBzH5pZ9Hw99f
TRmQOVT9kOTgNFgK9dlbHcvoahK28u3ZQLE8/kou0JTndeUqabod2hnu8m2bG6ObI59ShN8RCDL2
c4RwIRemwZvGdCIAfITmOFj5k8kUrpEla5a66iY//Foez4YGn0YKHTpTt0Id1LNl/chju3egUhZ2
GkpgyI/7ODnbhPIHkT0qIiq0b9gojXeJRAdMOHjHBN9SB3e569VOoCOc4K8tb1fkFfFUSUkNDuCW
EZ8fITU0id4k4ovqB0VT0CmoVrF8cX4hs/b1EfigskGZB7YyJUALq1IW+nU8cbKkMpRoKeOdeZvp
FhfhLDm5mtb0Xj2XUaQzsAjtKzX4WjGLGFSTJuWb9kqGB222kUj9AL0/Itm/JNfTy6h0QSWeGIfU
1LRxK8Q0oY7eXyB5XUNWQlqHj8YBml+hd13MBI5ULCNGbbw4lDUXDGCL5IpZiF8CW4iB6g2/iyYy
5pUxF6ETBxdiFsqbXpAFzi7YHHFi7nRgQCM5nJZfKwo1KxdL9wt5CIeviwrSUnToXRtBu4z5y5So
7HarNUN9AKB4G+U1QjbhQwugNaLKC2Trkq+o5wZKJgM6tYzB8YMqnklgYYBbzPl/NBrYSlRnZIjn
5KA9rCNYubbp++qLIoH29MhXZV5izNLAYHUnCDm6XLzBEZ5RXS6JcVJrMLgo561AL4jmw+phJ1Li
ZMHaRd2fRgyXPb9hSFvGz/664Pt5HYfHwnHu5x2viRRDWSUZ5+4R8lRRUFcP0TDyuR1fbToqXNk0
ezbblwzkUaOC0LVQwFLkLu01R5FkBQ1h2T0OENTjWCuB/wdMooYBsNbZ59RmIfsqkMcEkgmh9M3s
DSLsHP8UU4lJhfS0E9C25IvgAWUBGVMqhcCu1sxY5F1NhjThI/+/Dtf1hZHu/Ma0t6BgxgoNnPul
iYPU3LAZt/xsQalDD9S4qUIhk2n6rpE/8xhNbqL6jPbJqgyfF9Kx0QlRZxhRmyydJZdiAEyObMab
elF0tJVDdGh/CJgmXl6u7yXLUMxQpIv/M6psx2+aR1DDxBWI94JX2wqlrjt8hedMH5OkBdHh52CA
CLzsFg0kssimw0KYVKWOyn5OVXdQnc64uE1sTPK3DGYe5MCuO8FvdG/+3vDSvmzf4Mgv44L9gllR
KMkZNW2LZxoVMtNRbaPKHZ211w2o4JZ+HrQ3/tkOM00SezQ1K+cZyYVbl9YbhbtzWM5fbWoz14Ay
xjrf8li3DIoLJE1b6zfHIET2O0jTxeYZE+QpUnmKK5dTtH6uhe1p9pQ6LsKqLZA2SRb2qcFCgEdA
m5RvdmcqB9UxXAa54AmGtvohSuxW03z1F6tUB2kFBWZsN1Aytu8f2Ngk9/WToxQbVtTqaBLZTplv
mGnnDr7oKx5bZGOxj+YGGNlC9TenqnnxTc2Ap/KoyOCimXeLN7lFI5o8wdeMcIvAr5kipkAY/8Yg
wPuNYwvZigNcoXtP464B8RCXEhUdaHq8W5++OXliJVMeAYGLyZOr/lnXWQDQqt9JDwR5M7xEakcV
TLdce9AIrGXijOZ8vEE4d8WSAzXgnkproxZ2VoGWe3UPEfknufxIqIktmzfGf1BFlqcKML/wRYLS
4ofuyEmDD/jMsWHmFjnVO8zP3Z/uh3XMWNH84DMCNxxfF1GXWzx7gBFnDVd28hXstqcFnYbcc7oV
bS5fTXj6SmFfwbmUkAniCbspAWBwNUmeAOcJauCJSAKShQlJn8T4x9bcYC0haAKbcoOu3juWoPyK
eS8TzJZafvInV02j/hRH8jZu+OSz5juQmyTKPFXasV+q+ixLb5kbHB3RXzhHbm7j/BdvVSOHdDq5
LHHsXAJY49/en0wPnbxpolrk1xnfbABmVhsVd9Urff0eHNmqYw7o1x+7Tl7qIV/FwD61eDbqT9If
k94NplXmyHTyodp+aT6YgCEiumSOWSpT5e5bcBMaWVG7X7Ida4JCyLtQknuNfqIyAfWt4QW4e+n+
XjRbgQqNb1uF9uVOAQCuTJjYNo5M2Hi+G3IUw9YTY1T9vBZB5LNcfS/MM2tMagKtq1kPWyM015Kf
SDHe6OT//r3X0a9l4WCoOdBGVlpn7InCDsjfF8W9jk8QBrfYiZAIl9Z7tWYnbTKPHHHb7V64WgCj
/lkEYU4F5ihRW6B2mbJXNyaq0ck05SgyNQmXUUCXEygHWu8glMKqVlsVi1+Z6tYmmkXHA07EFSVd
V9OAte4NDAYTSALwzBjgFVdElui0aQBILgCukuoPwtsrGcxZkEooBjNM067tlqUjP5UPeyCxHqju
JaZt0uf543lA/IYVSYH7CpTeRwM4xiu0hc6By3bpBW5xBD6bPhXSCRmZrqci3DQWYoYpDdflC44t
XrLWQldmgpCIMlryTiTAy89gkRZrV0ZXh2wTn2vqOQlkVELwNKmZdzTkNiRCj+MKH0MSdkMzHon2
rhvSuwfasN3ePXWL9XTOhiy2qoKpyZSkLZW7jrMgbfwkOn/p94996iDBNyduu1MauDMAogde9x0b
F/gx6+z/Ylp/bTeRW35TpIUiFqxjyNMJp5EMIRFbDSJUxuTsvjeA6xBYnnUGR4BGxC2OVUBUxPCb
qI39iepseXEMZyUvMzGzJg8zI9mcgvARKU+1ml0Krfonix759getAFzCSG0Nw8L0nbhnDOCsGvkJ
r8rDiHD14CN98kJm/Jb+1TQO4lPRJd0S5JcnwAmX3eJdFzCQv/MlfUN4OyS8AYr9jun/Yy7hmaPz
YEETS94rSKrPB2QzmhHyae1ImoV+X26eseigU3MgwsNdegJp4UueoJPXqEpTgBWiWkKONprC4oMP
1ythUS4lwkH1VzjNklXIzA3QcmMj+ygS8wzwtMC+P55ehwsQ/I62K7xnhhaXed9LFXH0hD5lD+BW
WvV73+0KKwyj6bdmrTH6STiqkEe/PLk+wbi5f07DuK74iUQM30tAXPmEs+BIRgcu2jp3rTc/AGkU
X2L+1H7C1cjwYyUAT1CnVRedI1Cb1+15C1AUZqwvxBZ+Pt3V+N85rzyTlAiLQqkHVz/7DjvG9Sig
XgeGdJO24HC8KGgQSkAa8oE9Mp3/bh3d/cIUs0ANC39Cf4fFCx7+0JlXo5CAwtn3yWM9T0nSDPYr
MZ50yZsSwgbCOpzk6NUEmJFz2tWoYINhUiMveGKeR3V0HbnZ5e1Xt1khlNnEGZsFCB0aRc7DKxQh
7nBymfLoToYMC9VE1WOhXQxMbI21yXzKqQRCgOadEyRV/oguF6VLiyYaUVYiJ5AN8EIIl7D3Wggf
VHDRLK5HKyWwCxKHGKp+rb3vQkSP7kxyDWeRIix+fjWHnMtbRSNl7QWFfuJadl/MchCxua0Tdhtu
Ii50VuoPvlnDRxoSn1Rs9SbzNcKoVHs9XMCCUH5Cr3WGNhwmsNAdLFL4m6meJKYrXCyajK8VG43/
Yf6U7AyYJkVbNHPWjLAQUcJO4CAlRA3o61HPZhXd9+T9iSqGkPPmj8GwiMVDEq4JO5l/KXUGcHjK
yXIIJ0RhvVYUmrO4QpgqXlvJEeGzCSmEphsBCwpj4B3O9NlmD40dUHYP426K0U1iAijWKe/gh0LG
4c8cQef5eKiFnowuuzL/ZAjW58F0l6sZV9UO7UA82v/EElPtjeWcgkzkuVZ2FXLbYcOFSnUZRMfe
2nG9cMcO0dedolDxqrpaMxqAddor+6L26W0ApG3qRRBmpBX9K5RzWxyl0bXVmZ1mvTQCgnTJF7mJ
Y7NIOpXYdZ85eYTfjoLhZBDQZ1bLh3bjomEDOT4oW5s9H2EIC/NiIsmPhfCrJqPU3RG2j0qoybNw
8mmyzJGWrbxQqL8+QHIS4d2ADjUr8ysyE0X4nhJ5h8MTZMb1rIepTh4S+cqWXjZMyerKBbuoYHcf
zo/LpYSA7cklKd5KqjNBH+Q7E/vtfcUr4qyCppedic/AU6VVq1UHnMyfZcH307B4lAbpZt5c3wrJ
3E+yVmJ5A45CW75gD1Azx4yccbW6z2Bezeu/NW3emg8HdHwFqKdDF/rKweHHWUpZZ0UlKi2sk83b
0RXIKgdMg8d0Z/jcrTCUZTavyR9tCTxKD69HC6ByWFif+qxKPn6CyTn/hscF0IPuTERK9xlid8vi
Nq+hk7pzBcizmM+NuF0Vj9ArmojtMFlPgHZbP/Xjr0L6xyGHfLHCsFVm9HEVnBLzvB7oKaf5lF9R
l6Ilb+ZOfuo8xi0F8Xk/eLlbeqztC77KmLtt7Yu6FhI9v3NeVgObBb++SwRAD6qyImnnnqXpHeEa
2OsMm/2lsRUli3bpnJwJzYAXmzfP7vkW/MrGe5OKb1mO3jnCta82P7jeB5FwLM1zVqnE/CbMhyaV
a6EFz6xB+VLZjpIORlc3+sITvm2t/PxSOg4348+KTD8GEkHi74m9oVQhY1wGqa0bVqi64v6odjmp
i7TWNvI91w/hvYeGSUlmo9kl07JDsRVl+u4IHwavCQPxksGkVHjuSyQGFk/YcvgjWQXNuhsrs5rJ
//UUZU37Nc0bTaTQbusH7F5gOhlvwicLYjwNYZH6i/2SblhemTTiJ1t09/eBBIUnn0gyRQThc2ME
0wLxT8MyVkgXDOtIO8shhwkcMC2DX9nuyhDTENZ9CIyBXUuVuE2gFkahZBSOdgWU3CMU2Vuj4E1Z
6q2Ah7Gxz3cgD1heQ4i4IabdMDbbOQeGvKoGiaZZqSdWvVrJyHfi2QCF28Vnx21JcUU1md3kZGuZ
4C9Fo0xa/0COQLr7TZG2MGOO3SnT6DuUEuz8Z/w3GV1c2fpxCJiGpK5TjOSG2rO85am8q0vvxgFG
/0S/jBzoscarq/Ci/18I6VHSYh3Gx1U9notvdwz+4McgvOKbj3YboIg32yWukfn2svdbQubIKiYM
WvB9BltYvrYUFcbgw/BrMRVW4NfkVXQhT8NV0FnlkjOsy/rvkGHSi3umAalPInJrRTFyAkBiHs/Y
1JMTU2OfP1v1qRM/S7KzTunOm8FV5jNc6rM2I1Tfaz01d2w1V7i8iIZWsvWCKoI0cfcdY6ATjMVc
/RUwt/hyM+qQZ1mLbs8a0FujeYGDwJ8fK0VrGkzKHIQSIyVVKOo7xXlc7HddFgBiN/pHiX4uhe2O
R30f+r+kApEByxrhoAKMSwPFbdBPXFHNCiUaQN+RdnBv9R2pDRcfNGvEgA3VNbhiWIMVYv5wb+fX
AcyYErIJ6OOAN5lvQaonh0QfD5GIOkUYpILD3VkYefliC4ngfVAe0+ZUfibrYjepez9LzC0b4yj9
Li0aKWQoHe9f+8kbb68eteJVaI2b8+2/1fQQGbrmU1sh+VNz+5KaW8O+e+PaLX++jVw/IZztsgX4
E+pwLJVIXnZEOaqaxTDyTjtu+Gepb8Rw2g3KJQ7oRPuaxVY1FdoeJvc2gN+qTizm/aAWZvE4V8lk
Jzwqo1H6Ln/tnNkI7rPgIl4CUJkzTokYgzQtNedGXLx47cXWYrOK3iflQ3HTfM9QMMdX5xrCtXrJ
jQ6wDQECBfvK12yM5fGOR8Q2M4PqTpRDWNr6fFGjXVBHgW1VjPTIvAtt/G4BawZxDI+0eGJUjo/g
GQnGjoRXLyykVDKsIKrQjdHkFmSGdBGyx4SJj3LD2i0JUl34W/vatduhPoZINMygrqrPsycSa7Fi
fmzOOyOmuORaz0/Sz7yj9RwPWC3XelexwMRrZvadnUsrUCRULaRvfdN7PzTi3AFkWfyROBdnMVrB
oSL5QX0iiJ5VennGcr/FUOE3bu0NuVa7ThQTcwU47Gcrs9MBRquLd/hQZtJSTZKwg8Q3r7+B3KA5
T0ud9now6W9kNBXU4wxidyZj9iI2jdmyUl9HzMSwS4FXQ5dDJ+tYtY6OJESwMn3NG2CYiA9v6APM
JQM0qcgmJBWSsCZOX8AiXVE0JV2TOkdbCbKYM0TWAEOByl8cxizpwt4wXHMZMT3GOTqbRuBWFj/8
9kdH+OdOqviYPCznTFHeP1/u6N9Yk4a7imD01yzIO6EFBYXMjWsI3bLcu/qiqFzbvql9QxRnsdOp
JdIv5XnXNeIlUQEitSzglkFGbfHzAgBEVf0ju7KlNXzlV1e7Iqv9O41POlTMJihtNr1c2DEaozfE
wYneUP5T4TZlZ7bc+RD6G6EUro7ayUrQQgBF7Nvic+CzUMEJ8+IhsixP8tGVHkyJ3YD4gTqdtiXS
KxVnrBmWoJxMaQ46pH0W+EV/vTN83nHPWo+edw8ClHhiARFslOn1DfWVwLJy9JhRkyKqytfdUVDQ
AhEusomk4nkO09hCXjQx4bKpbSo3QRhpmQi31+8Cud4XjiABL3nmpE06OI5PfLb60WlOgyWWfooy
SHWSzJFYjJ+XzQa7Cq3fwrCVJ1q4rcUmgQJ8sqQiZpKVIONR8c002pXqwROnSY1Yw4AnANyFWYof
nzubpZ8/co+QqVYKNAE8D+pGP/X78YLDz/xh8s39aOde7OwXuekxtWiT+y25uebf/rXDx4IwizrE
8iqUNoq2OTQK0HuVwl5qD2gQCCAqwV7Q5nwiCYKcTM+dFgepkjTceADV8NCYJAvxr6qIJ+JsA1OL
Qaz5gW40zQzti2kLhA/9F2iQantpDsGUlhoMW2hzmdFNNXs6eQJnXwGg8J9nzG0C+MbjhOKrFxhh
hlDzlmMq1L6KD6m3mnddtYAkWtHENvy4LJ4Avxc7jUOQJHAaddzlcxNUyD2VCGaIntMPbWRJITsS
Q7ts0UeW5CkgAr/+NVvnAzpk9G4LKHmtpeBoB/XU3cnACL/9rJ2WiAML6QA9RWt7pJi+uB8Hi7gz
z5bnABir39/cc306i3WXukzU1kh3KUHAXkWa763BQ3+fnj1VaCvWMUzA2wMFm+0qPv4TCOdVvTqH
5K9IgfRCMKVQTiHFRi+hwUX3QoG01svtl0sjHYceU99TxXBexztzPCiwrhCYW9c8eF5mfe7L4Fpv
RFxGw3PYEcorAalXHwl8ufcCpDs/fydxeCtfteLNN2yE6lKXu2IBjWSlhNiYNa9Yut3eWXkjC6vr
p9vKJ10EukJYT88slodSc+LRixxqIOPoMFlX4umT/X3X62+b6NG5+KckEpeN0SmNOGlph5EHExV6
6dOcBsfC6HrGxdj2dPr04DSxQwSeS9v7sijXX7Tls2MNpDusXeeXggBjBRBsleHNxg/8PbE3oeNd
HSNWDj7BQPoL5CQqT8yIDDuUvNBQpP1oFBbDavMjRL7sk4TPGbhulPTSPmf3tsGMbWpB3kEf67eI
UiUZLuiOpnhsGtjQN5dv3znVvivmNZgDuDJe9vDXbalbq2BKsq6pustGbybe86M0vhdlQ0F4X9/X
G32CXxwr8jGausIMjAQcGxShFZ7YYhwNyRuecO5O9gxibghkUnVwIiskCXu8EDm0J0aEMn9pllvC
1NBsimyshT9eZZF4nT5QILBTCWlqNBK9Sv562MxjciR9ij4c78CF+v4BvzSkuvIjXJAJovlVtQ04
lNLKO09dJPXwAoKt7lirGv1L023F/wyIyy8Eiu1OHSLNIYaRVNezpJ5hfQ0Gsrt26OlbFCP5K6Z2
OW+DP10EzLdGIvdYVdLUz4g5zO+G1LBNlS3M/HbxFtsrrG/5hzTFQ6hRxmHxyMLMIbl2No0gz+XZ
FJNbKCkkXvM/3PifQwfXRhi7qtYI0lEM7p+Anng6ndUeIAQT9WxCKYcfMRuXPOCYGi2/HObkOlc/
7BO1Uz6xRI4UrEREgegofghr67W1+aEhwZamhf0Hd7db5R58tTCMzI9tFSejDDvKTTlN/OsNTZWy
pMUQN9xksK0w6R6jU6kgK+nKEoOwDrruDpEE4kNaHtiMabnafJwD4AmNQAzqJUa1S9vBi9jrRbU7
xAXklPG7lDEJPFi3Y1wY8ydcYRKjd5J5eAAwwYic18CQI4UfizEk7xjLC3OycGdk4prQzsp/XlW3
GUvqMEeOJoKQ8xjKb3Rs45SuKeQawH0prAEiuQ/tGTbE/Jv4N9lrCldqLeBDm4U1z8Cj/chwd/Fx
vP4kMIFfWKcdrw8ZbXq3m9AvZq9ZdXlc1jSC+HeWxVLEmcWviQfrC2KwFzdWrY3DRwzhKqHkh64j
wPzXAW6PnQP0+vEImYOdw3aKfjjY4jJ99AONLK+F02r94PFgRNaOaH/A5sCULOBAiK4S9stULpI6
ggPlaCrdmwTzl0IMitJp5or826kJNdkq0hP4SBUoR/Z6XqmjO6+J2SkWn8u+suquc9X3EZICSNzM
xwBaU/JLtnRWCRqS7bNGMRfPdYRBzDAfEovMG9vpLdJFRO7aeVgJeid5xPiDbz+AAZ+yYt1k3PoP
YPU4gEQgBvH0lW9N9olxSXIrELxz8206LAtoceQXB/4NgxNSh/BmxNl6FUcVePC0NrqXfyRDuXSV
FzpnQ+TputBv1xzyrr/QwqDV2r5YP3oom8tWqEvgaftJbEgRXdiE/KP9/6iZ2M/z0e9mgWKVxr+k
q9hnnhSNLBuhhIazs3FgXAMPca6vATlCc7KItQltocsAo/ge1C9ViPTbHIh5sS1+Y9ne7+CWqVQH
caQbhyj/TBapXVqqclRtMOI9meJREJ0KRr0IJiEhUNPOg7odlZtG6L+g09Ub12tHdMCQitmLDybN
CjMKnIDn22nX0YCYlrD5okFlZsuYuZqahGM3S5cbb+ireJqk/f2rAF88tOgkwOxFldAL+EwHEbeH
9eF104NHJArwVu9PwIz1mAR4bLM1XOu7YyECIzKCH3tlIXTj+40YkP2TPBvE+siotYQa5s9UiU51
bkN+T5GUk2LN90mspukPUOe0TXSUbWizAngNPXC3cEw56+xXUFqlXfQIv1SNBgNEwO++GO6E8alM
bRzWrwId+guBgdrYlPyU4EYR3COAo2TTP4JfTDqdfdkFMRpDdDKK2Nb4sFCxfFXZChgf/dqrevw9
RSaouE3HJw8Flc/mcdRmiVEgYrVwF33RNR1dADp4GiDHnbdxxGNswhEBCqtk+s9ici6J7HocTelK
eos1hYPjprX9qiw7gVbIsAoyXWJXev68PJ+t1rU3mHNhMmODLLVYTOeZflToKv45Q9I9ILnMQwEA
HldmhhUzxgrJRkAn5lbY/PNE2ZoSElDMguwmLRAWRndcuy1/8rBdgZCssDP+mYSD1fX6c6KEiEiK
75g1orOkvdJSUMWhPYW5/DX//Zs3ql2kyMx6jW7Vx9ockYK/KFxBaBLKzT3jwyXl42Z3cq8XD1S/
6Tpy0XSyd6tL44O+oC4TUIdF9Uvdsx6wRCkdlnFGXtjTNnm4/JWdZbUrQnCuwQQnuszbaI5sWmIA
fSNMWtV0PURsUOpaad+DQAxV/Gb79ZV4/4iC8fgh3C52Hf+8xqWpnBt4Pf7bvEPwMefQSDX8OfQN
EnWfR4g6H3VK5hwFqLuaadxBvT0WJN/39rmGdhOjKZgY7ilV2VfsLGC9KcREkYpyX4SKUpbfy3ko
HIwtpxS6SyGZMOC2F1J/c4NLQy3GqlCrMsL0geqnuwL+BfidtW1HmZU4HKEMbuFGQdX0x1m/FuQC
oSnhlZzNLOMwCntjSMIdn/peiyGHOaQrZk54Z+BXH8A1qgtCzBU9aWMhHzTsNKz4cz8dZoyBYRJc
krTpHkFYTXmP/MpciJLuclYDcqXUJM/rqcVHo/AsohZBkZnBnEVtTvnCU8y8xJNZ4wgvWTD630zL
3/6kqHJKlBjk2szC6Jf/QOR2ITI+nPMjAJCgRSTRikGCCK6GpimZR+CV1FRMLLtVY5fAXS6ml0ki
fjm4MUe4NkH+vuwmxk5spSQWZxJ4L6gXlHbCIUeg8S/NfRpC9IquiDa9XqIXxdq4UQ6b5gK91GR7
7eXm9FN3SC+HCThafzV28o7l85M+upTBamrKLGYzlyD5hifW8T2j0GEgXaCjVA+W0j6zwC1v7V8h
JinlTbqJDHdO6+KGmEvJPSGOwfec/NFcFrthtQUnT1gFMHrfB31d15bSJd8rAqfw+JfeQbicXSlG
941XtO2dTauqfeX8l13JmB36ohusD9xbtFE0Cx3H4/rbe4DBpuvIXGJwhyG01cjJiFJdZJpwr8XX
CnqTS6Mj6nvn1I6yitWrf2ifbcQtPUdsnuwnFk5QY7ozk/TKahVCCdbqVFLcOQryTccuHTAsC9oQ
Om4jpMbmkR196p/7m+yOjJknRdWxLbhGD0t9uHCHn+M96CwjX3Q2h/QLAfp/Lfo36OPIMrY+ybkh
tnt0/iu6aBgYnFbEORjwEvJd5/TOxedJt2egXfGdfIa22P0W6vxh/nIPq9fix+5+4JvcujlI0mk5
xMH1lTFEOacmrLgPyMiVyYUB3s2pZKWWki09GT69OTJg3eOtTBWhD5rdR1wX6IrnORX/a2CdYr79
c25YqLfatk5S7sIhwQdnQaOKVLtnPD4PUdY1tHb+4vOFnzvjCZjyVdgD0yvy2Zmq0gtsVCbh1xBk
bIytnh1zpDnxiiabd7fM3Rhhu31Cqav09zkXrwiKSN1zJunHrNdG4CXDi4TXGqPpQio5hniZvdii
d+JLW3MwmQcEeDSq9lqdh+ek1rbT83fX8Amf2nFaxmvuXgG6bzJZwsPt+OMq+dJYfmwZ9VTdS8ei
VWQIueBHl84uBpV+qb7R3YgcbMB0o0RXbnSzARs4mEgWtaZzcKrZqsMjs06njokY9eLpnb/WyVwH
XCRaQYgf1u1f5IH5W74iO+OYgq6Xa9nQS692aPjs6ouJm6DHjMAmEilHamUHJic1lKpwlNSBnrw+
cu9Y2pnJZAJjWaPpdLjmGSh4F9ymSAWJZGzgRAbTxSQYYjskcUTiAPI+gOo124Oxse/RwFSzJnw6
YpFVlAzrXUZi5XGQ5tum4NW/AmFve+tJGHBbvT5DW3OLz+PnMOa+wDZWuCtxqRJEOmFK3Z4bnmM+
M9R0QgAitB0d3Bd8U3CF/JwIJoeSq5ehHI4TUXbWO8a07lgNLwv8rCWJFfuez6xkH7hG0/RKVTxM
zydlsc0jVqWPrmCEipZUIHylDxiMqxAtjtlMTONJ4Kk+WfcY3G/yV5f6sh/GFTJ8uqGUntvWsSzD
S32uC1Yq0TIGGzh88C6InFjw5sfe/tYSk65xDUfzXazzClDDpNJ4xacGJujaDKyXck9DATqAjW+h
ixK7gekc9qe4w/Br07wXbTEH3TuXddGLer+nZ7e0/AryFAFkpY17Q1KOgLMryHPwUALHt7E+vov4
nH88wIyeApEuGm3teuPZdcMrDWt6C5milcbLXGcZjBpWaBVYmMUY8E0Fq8GMox82d0Kfy45KPrY5
ZWWPsNRWM3olNkSQRl8+RWuL7fLbrhHJunaUvJlYcompDEq3vz6Aid54dotopENjbYPWIyo/KAql
5vf71Ko4jdPp1rjFLFQd5KKAtCL1VG4zJ/fjHEMPJ834Yng2GiyFNjqK7QAnzQWDh4UIgk82Or5k
AYFXRrA2pu4TEvvF3j6rLhnZxUcOldxYvgUS9Kesz82tzhJTiktlKS3kpw5TUQ5axRfHRVL0bmvo
0ABKGJyFyUS12YjMy62aGja1CrvIsAmUUoUsSi8CD3JEsFz3HmPRRGOcxmxYqjXEWFA8eeG5SwWU
KxtzRB0EREHSH6Ka8bUKHeRx1GM1CltiiDlqaEA0Z0Rp+MdKYb7t5MEcawr0FeDGL+8WCRtqSqQL
iZwJsJB6LLlm4RgOdIsDp6CtYme2ywmR9P2BmqLQscVgRietrUyDq6SbNfU8GA6VeRmeih/gaHRs
Z8KipqHAEP4MJLAxKtSpqgeUWVGb9F42WuQG+vip0wV2gFZbcwSIu7LLg5y8/P4jZjvMaR55m/Sx
YHttnqq8fDjEOXydaIvswxZdK6ErWdoB3+anNlYYypKMiyBAWivxHX12518qwjqX4FCNpVNy6WVl
Y+dtVHw3tRQ30c+MWiQVBMSIbwuQ62OoZG1Zw70nlIXukBfJ8YXwhv8+xMM/aho+u56JO86iIjc+
z4jQH7xhBSLtokFGT3LgHWCbgOOr0z5zlVeE86MAYI2UndXcbCCsS2H0reW1e5co/5KgaB6QQaWK
0YPF3eivKVrhwU8TDWDTtpAaGqbqaMwS9m4M3jgEjyruotJySnxZ0rwwl2W7zE8S8g0bzd/mS9po
gae9nXhzncoi5lTtRJGtQEyUAaw2N+mxOf1E+2w4E/g1ExzhroNT4KQ6GJjVl0kJWbol0FgHvvlM
j39D9B7zcrxuLavrVWY0UNXm5XCFIO2c1ZVi+ok41k0tqNDR988Dn/VPOpvX2iA2jnJQhV2ew/9c
17w1k72WN02Q+v0+7+l+o1eGt7YZYpEbvv89V3B/7PkLf6+CZblCJt9478EbJLxE2zSfV2Y+1FLW
0Kom2wvyKcknw6LwU4Ka5KbEwCsCQjS6LAAYoRjLR1Es9cTluZBHhFlbPnmNsYC6zX65nd+tXab6
8sDP8x1Lf2gTT5LVVA790EhFOoJEBEx3CPwr6G2mAbn8O+Wtaqyew0VemWRu14CekUn87Mu7BBE4
yaMOs4RGu9IAUJvrsTfjH2b2koulsLZPHhfamOk82PATFWtzuQ7FeaVMlrlQ36uOOTmHRapUduMQ
cKQ132pbHjr0exQuPd67an/YoRf0X2TlX86RX9epIhslyvFuVxAmh5iyCi6JhnQyl6Ie4Kx1Wdwk
1iXtkKiY+UdtP2V9MAtEfehSkBnPemb3eWg72lF6rvi+ZopR0vVRU78jRbUuB97HvJhdN07yr5hg
JQVcJ21mpmud8P/c9QWqdivl1GxKz5P3ka9jbBAN/lTT/zZ5bn7DOBis1oUr3moXQK5KgfKp/Ml0
OEQLS81CGDSecnKnZu2vf8fHRExxqddui+KLFg93cbgzjoQhIBNMIztyENG/7VGa7ygdmjTOdSXd
dMn86WQS7ziytpYzPb3VpAvUwJBoDNHgeJcNx/nDyGW2s8iPy8WosEhA52K3jzDI8B3JbcabjrgP
ocKh93lZ1xMAT66+MNbpXoiqkdCrq6ozSoXYvZ5VO5refAAHJHDsMzPReObPG/XLUcs1EKqYK3iV
emf4zvSrRb1AisR22rg4C50f9QpoIXNksf1GXBjq6mTkcPSkvq8yVAL3Q56dHnpjLAkyvMJpm4g7
jfuDXRlL7NiRIJhtnjcLvkSjft3pHzfIHUqitujNKoRmRWRzT6Vxsehh48KASMgwyx1duWogBX27
VTXm4Rf/T3FcpxghsDQ50LyFR/CUYEK4W1I9u5edvYXilNBTQ6UlULx05pEDy051si6NWbrnUbmc
QBTt8ed2EU9vFw+kUTjFbomsbzKBeOP8Z/jZNfaZ9RRaBpbrXaIdBOqXNnlHoqkjiCQJ42+FnKjE
UGEmV6HJ7QDWfa4eP33/s2ZKhcvxWNiud0RlnP78QNRwEx94P3UNYEFFQfTYC1w2r1VESGuWGzmy
3vobZqwl7R484xVqHVacU4bhuYg4DDtYoNRJ5rFAMGIrJK2CTlFUpucwwYb6AbcEws4JDlvgjXII
c9YB4zHCXReYTBH95sWDzknlrH3Km+DKtx32b+nDewJ68Fxi2iG3Mxq8VzSxUarDmrbEG2k/stKk
wvZ5MKPeGjX/PXCWiVuGUTfCrvJZKrN4/dSWVxNGANtw+qUQhimYx3oojtZwXzd3XNgYnYusO+KH
ZFR8ovCK1/PUdDzbmTmJlyvmKH4hgQYzJWRsM+kyRrdjDP83IxCMwEfEhD/Ory5ieXMe39vr+yyq
K+NxawwNnxBJX89Vd9j3S0DfykFb3lHt2g9ZPvm1svMiBbwGRuAxLUvg8V5kJEAJmqMxeNCDQuso
kMqP8puduOwUghdbs/A9ZAQ0kmGgG3Tn3v0pwrhf5tks9RyTm2AqHC0YUnf0iOunMi5EwqyfVz+R
+dZVvISgbssVFvCeD/1LajUfoOBvQ1qWSjvW9V61TiEf48/NOSETaGAAgCswhuWWdmf3Wvh7ouo5
LkXGWnzfI9W4q+2FLsMAEKjHVEESEPvD9EmZxiTn0fRFC/u2vYXWmCCK4/pKEYVlDfP6DWRnxW1V
R696oQRcTMUif+X8Erv+iYCZxxAfyrgXggFnt/LGt2hfeNHxzgWptoZl44Pi4RgAHEXL3VpQFUmJ
vkKBohGBlcv2+6109wUjqR2L9kFw9mxV3bKhoLd+Kt3TkX0Ywld5KHOIoJxUtBltpl8QTx3VWXze
2/Rj7exVW+AK+8pF/ITT7kEg2nmDTWrcKgiaWuxkoAE4k2RbmpR9j4p93/uayEwtb931mBfkK47h
hXAHK1vsijoZvFOb+UkDOb1fleyrRy2VaqABvJNd+EgrifoJ22zGIqr7Yxs4Qji4b/xWMmErJnoK
ddAYXES17oR1+3p4UpMr638PY5nPmdi1tTN6DUR7ttGbg3l1wGUySsSz6fQnpaPIfL4UWM5uR7I1
Pjx1+2vzswwMH8GN/TBvqOSDdld2TGgc5u/C+wwgled5IZVPPhrptsjOrDfbt52LaAksM2ew8j51
5MWL2By6q4AiRVZjcKMuUjaxz2XGAeuiTsznZ0RHOE0h8XwmR2jRE6PObElBhnFwAIkqWMthAU62
Egro/dsRErCGV0T4k6cic5RjdfVkqmDQ8h90YSQRi5/pZy4az1C9Dx29ZvP2MWiEHuG5WGszH+Bc
l0cverNAiMIMjphDl8bIkJBfoOjlRVyYywqhpAY34uiKSmXcEMDHdAcaEjUgmi8vF1Wq26Dl3bK9
fb8RXhscb+m0zVKcvFicbx8xZAFAqcXv3BMFhU5mG4Yadb+f/M0temA93nYTLC9OJfqu3+gwUrdU
ZrEqayGhzqMVCM9dzBqkIkOZVnRBFz+BAxzoRz2Fv4JWxIIKYrdraKladXNd55O1wqfgJRYAGL9Z
RYUI0NuUyvMQZ/043T+TwGkSwTSv3qazy0Uu+BACBwBaYiusikemJwHzMRxHkJwSwqNqpA356sx7
BfuOYUyyd4whn4Ln6lqONx5HvVUZQa0Vq1SWZ1hjvP2vXG2sLO922NDE8ilIDITjUOdZr5oW2ArU
4PJ+1hfo5mUHxLunSLNs27Vj7PHAAoFoxsgUHv+MqOAsh+YfuhdJs4+SouwuSut0y7KgudUzkkiH
GNQkbnKlpk1ZQWE1Yrvt7s8bjjqw7XZqBgaeBnPOt6+DTu0t+CpePrPDQW5y6i38XRvXHvJ8K8kV
gVwJgHX24K3z63bPifDnIIDcR2jZJCT9OfyCco7eKtTt3Vf8xGU++5+xtpPN7OUvWLLq7LWxdo3q
9pzPfggH3xO25F1AX9illPiAYH/hVruqp+rZTxCgZ1qxwRuLDXig31xfESlvXkg3a/FzcSuJSFHr
P0y9+GOZrU/swZ8xePsy6wemqGJ+W08ijFsgR2ONH3KfWqJLy2XlJ6y7nRBurUtf26gLb7g97nsZ
v5pGdTLgfEcMAXo5hcUoz24kH3dBewyS/VvhuvYlEfWB6AW+3IsI2tlWE92k59bn3JT9bkZA+jVI
V1IWnFzgYPa5uOWsNJlofVYgXQCT7zZQG2DrKObG3BFLuJuMrpF3KqjiaeAQnGDmPewtQ2rNusuj
+9OR8Ou6uMjxpuiFcCLMAy9MVa+Qu5dK/I73tbfNfRXf2gTkfIviLzO8qOR1X7RyGLmh359u1myW
bc/zc5SFt+/MvwNe7PJ9AwBeaQzITFUL9DZzzRk8vYW3n3CwvtzlaGRAOUU+H8b+DNe0bu6NJjXa
SVJBpvVfVdnrAgpKwhzD6jPaMRMHIiN5GG6Y/IP0mRjlGyIIQMDnSOPU2yWdIcY1Tm9kVC+c5VEV
6bqaEuo0TrnNGmIz5IW1z80/UGea0O9VcSJqjMl/7qjJNO3A1AnbrxDXWc343hlYGLSF8sL9qFIY
mB+YHZUj//3DL3p2qJSMkmRWYqpP3du8RYv8pvrZz49NLf8LDuzeZEM448prhatKZjnd7Wi0O6Y9
lvakHJPjc582/xpq3VUdWr66RYM8Lg2r/cB2fWtU7px1ip0J5B77I541brIDBMBliKcb5xZTUkHs
V1C+z2sCqiwDTIkCqTjRmF8QKeO/jnYx7tVYdKxjtwjY6mbdRNpvWdAhuvUqeilADQx7+G9Rklsq
vH4F1JTE2IbayMT2ofqTvgBPjemBl+UYhjkVC2crmQAWg7gwlaPp15fRFvrG8yu1s0hAsHrGdgNs
+SJA1pm0ihJ/L0GOQggq0OHaIcQNz++6DHXlXtAteoKUX0PBE86vQE9f+URZ8yIWeVs2nulrQ8Ma
7YLtovI9fSV11LovX599e8xgm1vd6iRwPCaMo75imZE0LOPxpdfS0HwBQ1o8DM7PxYw8MBknz9Sj
I5Jw+Cn+Qc2KCmaXSZ4JrK2707qPHwfEe8vosqxb9wsLiF7yXERwskQItYdRWqOLbbgZD8gqutb1
4jeqsyKRYlNwT97bWRplovsrR0SLVX6cjDZss/OipE4rbUPgDjQl/m6cVUYYW2tDllXRRNsz7hi8
TJfc/+xUuRakqvMR8+rj3mPAl/t67p5uLvqe/5fJwlw88jbVoGfTVOQYdDBnAMSWJ3CnbUwV62Qn
/UrOKqNvY8YWqd3BrC8HnwkGutLuVmKpG8XH4/2qTyu6vOz/vJsrm6nmEzhz6R8cHWy1QsKu1wpH
zEZH5UorDyCrN+WxqcNmF4R4Oa7u3BU9LLo0088AIe43bsLAsEeqsJCc99QR8NuIskkl+gcCWm4O
A0cTcGikuSMNvlyiExPNHV9Jo+Y4E9+ippE5a+6519OZ7/8XzpkCGe5G8OshW+6IxipWFgbhNquJ
XwVPYegg+h3SKORZYDfQJXYvRGGzYqKMv5Ny94JC80IQAQJvteMTLJfZJwKLmaCO9BkJbdIpXSad
aCgxSEDJf/ofGzdlE7cqX2P6XHK3RKJ0RXbLZIHPJUwthqnMIxUBNeR7bbRb0kOVkDmvSClfCbuQ
Hvd1cU6IlDPNF97rw4POKmESY5V+KA8LeZdhuloa0dyFVV3qujl+1gBQmTgnJ5xp3SyGKkrvdSoQ
AgkfVWAlLsz6M0s8MkwCUGYStkS1QmVXc8e3xFQEo6AEAkz8IYRJGhuvbXfGu4fMuABZBYIB03Lb
N7TqP+x8SjB0Daqt9h4SjtBatEuXD0CMnao6eBdvZjoxjYrLc5XVuGUiUUDvRHCjZ2JqXkbgNBFo
UF7VU63KZ4p88vzJ9RtcdSfe4cp9ieaEmDjKFTPizpF/prZuXszZnhl5lP+Qu8r6o0n1rc/g9ys8
5ulUhacpSvXuaJuz8jHGt9fxh4yKQ0T6bqnEKSGIiIBseS0BYSsLuzGx8osV9+6u2vZrGgILCGne
sbff647D8xlQZ/vLSdDnLJLH/RJVdsgWdUP0nN7I70UlB2SxD01pDfAm3v834gVbtUbNl+Siz7GD
ZOSYC5xJ68kVbSmsgBdtWVBSrQlhlRhH/Mch766vZNW7S7uG8CMWD7xLlMec8+G+hrhrGEyC6/EK
i8yMsN+2Nl/fELFLNNHg1ueBOk8t7yu7zYW/1yYCShVc8mctlBaZowWYhKNPY+6UaFR2laQEWTQi
5MQFxnyLGGCxcojrPmUe786qvJ5U/eDdi/pFyqp0GdaYcfRHedDWCFltZrjfVpssawIUYPX1jQOV
QG4m9znxYuD8/AvOaygE24J7Qj7SUUhZTEIUAAZnFDINfXew2SJc7UpmECLLNw4xQt4HOKzHs8mG
egNzgvAeVZ8IaBTcSk1TfkfpVM29oulWK0Dae2mtk6GtlusfNFesZH9ba0iJYOjKtx3M/kWz/laO
IdFC8zKDe+5PPRNpkHupqXQ8rNX6DEmUQ+wCn8paqx8WCTGX1ZDft286j1SxCFJbV51xkzYsXbTG
4lYaLmfvqWP+d7NLIxd7Vy2SdL+TpGegdHY9HF8xuhvxWcijT/DyW20oCrV2CUIvEowy3sZan0ij
y8Gh2uLMySsBmFLZrznxh/aT2vpBdKYEd89OqToH31HY//SviTh3vumasw/lsLZ/gGnsFMx+Gt4G
FlXZ6zQlzrl7w+ays/67eeV+lHoEXyrufD6GfKU4ly2Tpa9wTkUgB/8pno5s55I6xY5NBnkZqmZM
ZCVv7UoFLzjLVmoOJkzbO0jckde+MgNwkgCZiTw9eSTu8z3ma5B8OEbKauwdKrQaEFqQRUcisXTM
7/1hI9lFte2Dp+FoqdP+6eq8Zo9NE9JqrwRYdl0x9xec6ghjzHTt86wybak3GWlPbmyo+6V2MzKn
MI9g0hAW0kWS7xwMTB8kX/H7wII97JEYsDpchSzTfkYxa8BiJPTtMmJQuLE52e3yCpFHL/Zke1S5
saXq4SxOBeMtYAgtkH9tirtLMn5nP632Kh7msIn58lDxbpksX+BC9tJNrSkTabAmrzpCzF0cqXH7
TGgIyNBCDZNLieVlLStFiLaN89v3YHd2qgvGg4G817VDa/TMCHk4y+7lqTwJQubqwjG9sgFbss3D
CvIsBFp/6d1nI1rdzMNbMjYp1JXZGP9o/St8mODZwprAHIkh5vdXZtHGicBxGUYHXaQdRTiJmDaw
7lKqcfcZfeH+b9+0dLeUZjBmOFrSf/wKTWC1jX/XwcAXAEknolY3EBs9lixnz3JthICEhlVQcy3i
KPNsnUhdQfBD3Y0i93D3T9iqYaoiueJe0Zx5v08xM9ZTQhLFMnRcdNg5VNkdWQVyozAH7/KIt34+
GK8/X2g78SDY/8X9VukTQt+KSSxlRrzfaK91oKxwH+IfCHCx2w5znlqoSiUh8M45ETbOc5063VB4
bxO81bqQxWPiOVbQmNzn+d2CilmwdV7zwwFg7EuTZLG5Rsk2E7bdVFBw8fQmbJThv5eJfSHk3DvA
pcL2Pafo404uGkt7mUsLVkfcZxxcWaNeEodjM2veJUD6IHQy6TNVYoILQQAkGehkZiI8KjpBBLCx
0ZWAck+Nw7bv4xdwQJ7J/05/nLiWOzt6btdwkFAKOVS+K6Bj0eB9XBUQCl0TV85nPthYq1HyIkVN
GTa+hIU77X58ukgNz2hb2IwWcAJuXq0uSZf+frR/m6xwszEAyO/Bq7S5h9n6HkDyF+o9lG+8t9hd
My25Z7pbSgKaUWGfItIX6Wvpf7XCe+fI+72Y+9QvrTGzLgx7Aa5VdTwvKIi6z1wgqSxFPja1bJIz
wAMYnSlye0clqgenkdzs63nEtAE8kKowuODzc1IaAKxJj3t1dDj/2RAtnCKzI861NuGVLndPuSBs
3py+lA08faAnJTgvaiishLC9iaPSIUZI2l7siWKsCAWlDqTmG7Oxz5esiChovxtfV8ic365aLQir
TpFZQbZrVTUBhgztTx1PkAQDkpkbU7NFywp5vaOyOzZ5N3MGfE6oVsZ7ZZd3y97RjDuwq/zO7VVn
TMCheg99NZNZu7bn0O7fr/YLPHMP8FwFjFuzk1CQS+0cMKA6gwQ+LcD3Jco06OLJdGjOL3I3EHoc
Q6zsIy1dbz0N4s9gYyseUEaIzgUQ1IL7EDgvjD7X7vyIEs6oROdydTsTwnopfLJnUgwrvVCbPn9f
gcLHcEzfpCOeMBLVDVcxsMlARnPExCzwKfe9ogfAb3ZvGbSYaKn4AZFUjDtv0G49dr94vV86vasS
5LPG4whB5Azwqbtb52a3DQ3xGz7rtE/8rLNE7phMi8uliphubIqIb3iLdJDGAa/+IyPlnOEN3atr
nzmz0TBHRf0SgkJAy94x2Wuh7t6es5x2KnUhRQm1g4psSY0vqObsYV04TjK19TuawCFQfeszcXHU
TefNQZPm+KGqkOI2Fp5kqBbx2nDMWFYyWE5Nh5mHdUMeZHAHz2Vw6xVKaUcDpdlqig7Vf38Pswn1
5kSvjw/k/wtf4mafiMW+ipkuCaMXkMukpc+xumTkDCPBPkZ0+9JC31sqwfOpoO6ORaRiVyKyFOM8
5Z9OzDHmL569uBNU5ppWzgO51OMrfsktlU9u2KVYGb3J6AWUT7SPIRFni++07dYChysJToAHsRhH
vX9r61CNqjZmXxs6UeuEJOwSYBoSZ52xNylimDm4C6b9tdr2/M9YiYch2UvT+6Ucj7vraeMih9h9
MDD4HGZAkHpOzINVfWO9u0N7BrL0vso4THQvRRuFO5ewIIU5FQPjlETne2lLmOdGrJikcHAmZLGK
bbF6ZgvEmHAA7HcbsIhHi++Vh1867OnZLTP8BgcCF/dik/ujx4cg6mzeTJDgRZVdKT0kmGWcC/Zf
7LCPLmgdMMcFvGJhm3xYlYxjq9kSpDwmC/gp7/s+/lmoxDrgqB7IUUtEu9uDQBLBi2iWuKX6vybS
nYeOw7LLaYu2uptHRwZZH8/4O+Yz3xWI8HGAQ3Yr4V81cPVMNiXLssSrDj19g5j88SemxL71LwDv
aCHDGe/bTmOR89IfKM8Fxi2H14+eRChQ+RH6XdnJStLRCth6xQa3gfZj7N4PPNNrpDC/PqBYx4Eb
gqXi+YfydnSWo+qt0hIjuGYLGF6TVOWnbB5nvwNh/1yHtcewRu8T5/sZKY/rOW+jOjapiJmEymKt
umUt9m7iHTAvEl4ps/ffPMCyitL6nL4WATNjmmRb+lEq+WDJc35mSHDqItfmCEiu/9PevxwTwomB
fiWzFImoEZ4gDSILjc9kDOdaB+2Sum1jYUyIA779qtQ+XCFnEN+SuWmYjIPX0e5xb2iRZY05Dzy1
/N3ZaQddVltfGAJ95bULuFG6ICEp1z69PVv07Sy1BnDfXUi6Uc1JPCzuILQB60Ux/FGzkwvKDUM7
G6whcLOHlh2CZEGm/NSuVs84dAQ/fDvK6IecVPh1Ay9dKUxMGOD8B3ysWmR0xvVf7OhFmfU/GPfH
LdQRCc6/yzsVLtj0LO+kF22MJKdmgvql+usCaRtKLR7pjxI7JloXOi9CwHhSCFK58/10C2QL6ISn
gHfyJ5nx4DGd4NaQ+TxW2eUJjt4U/YS2yDPv62DXszhPbWxKMSAY7Kw2ZXSGkOR/qFMpB15Xb+dF
w0Ndm1pIoiQUff4aTLn+PK7Hu5aE6Vg30UIhC1znAvu5Fh8q23XmINkz5eF2/A96rWg+fwylAnQI
XjVlakvbNMxMilqyRcJgEF87MR6Rk8D+ma5GVbuAHepbF3gFcHoK7vc4sJ/R8NYDfOL4dx+Ylqc5
LJ3MxjvHv/rrYe5leRxAoOTH17fc3tDThOMNgTZRDKQM02+dOZMS+gkOWzg0PbhbXuG62LtFOld9
FS/MGwW6zFjCVVbeAyyi7gp4yAE1hKL3vurCrLvvtsbCNFFz2bOgHdsBVhf2YBKrXiu3+R13/JCy
ZjDPEZffkeHhxIDoMoccrwimr8jo6+qFEqzurtVMemdOgvYyroZssYOg/q7zTh32Dgi6RmqyFBnL
SHPugdXr9ZI9W5DgoSGmc1+XHMlGkZrxviXAlvGBNAuMoSuWK2ZiGuP+vZFTREnfMOlC/Fhi52jB
lEcpMX/f3OhKjPFAbCJrTCTnuk3P8Jho+FZO6g2oBxj0MCMIIhe4Rs55bcmneD/NV3Ywwzdh5ZA8
AopUFnK3Fwc3L3N9K6Xdl/oTuIEwJaKRb5Zsk+1aDUkWqJB9ntP1vobw7XCb9QiGfZJyf4FsGhDH
L4OZZ3mlpQkrfpVBDfaSRf5IokeINaL4Gcs0fGkMU9QGo2k/+P9yxQZu3jPy+MCC1VxjIqigWoAy
W3iTbUhE5EU1sxkSCcTorvtK5GRUqKzb6+U0iSkGWQReEZriMCLRGBczExT17hCiMWTbMhquqet4
VRui97idXumHxS7ni6QwOs1e2NC1qomZLlNJ4Yt0yZZjqux3V69BHy1ZwXPKVH40atYZdmwnFICk
s/mzBPIUZdtuTZwm9cMQFcgk2iUcB461bs1fkWPtFnQlZn68Cj5c8MiIsl4Yym7jpo7nRR+5cA5L
pSvSzPQSpjp41VwYKdyo+PJxAACKc1GwqIBPL4r4ic+UeAScW6NVP6wOfvObuEf4E2xOwPbJpbF3
ywf5IDLmUAkRx9865j71P0hTgadvVYRhqkVgF26by55Nmc0tjoc2GXQstmkZKtIFpT3FXiBCmNCX
tKpWqt5ORPD6pM5H6jC4U55702uxQ1UFed+54HEtopg8iKflZZF5JHuY83iyUt6F5EbQVaAPUqRO
TzMEB6OvUcqO4+iomvZ7tHgo7tpcSQiqR+JOB8MJGn34jk+n39av2OlWCyhSKKYl0tvZFoExGlB3
QJaV+PajVlIAf/hwMeC9/hM7aKO8TOMVwxyZCYGoon+CGA7QrJdHwWb6aRUZ9nPPsHSOtHAhVLuy
yyxkPyRwU5gWIi3AZrWKEBu4GQJnRxiK7IpVselFJnWM20z1iq5ViHPAkLlVZ3gQai6bog/RE1HK
KSgVU2oeYP6HUyfMnEpYN9Kz1jJsi+8n9Jvo4pfQmcQU6S/UhIMLa0u13iEAKEeRU0Hq2BDIATiq
drHjKDN9CSdcH6gQTIJrR04eWWOjiOx6Kr9CrAxtnq1KEU9bfm/KR9qgVCJK1tgLJ8uIfeWVPeVE
TphWkeW0/fmLGJ20m65D25MPZ+7tSq9PGeorFczkLwtL9YE5v8eT+klkXpZgjxb3YpQyFH1+93hA
sdnwJQn6op6pNGrkLSUPvyZHv3ob/BOdn2t1VUc7C7q3E4vBDCz2dBwMQ6Xsxf93IynG7VFqqVPD
E9V+2LJEbf0E0TI7f6rlzu79hB2/fW2l54bQGXko5u1khns/Cc73TeDLtjjzfbLoA/TZU23YtkyC
fEQPmBBS7wO6O8n86Stf40CQtFlSHWiI6JWSclIfStjGxWdTo66HqqUToI7YBXTQ8eYfJW9CHVgi
cxVlS+Xk1w6hr0iaVxZeVuESK7qQgpswrDGUXzfB0Oe7VL15ker2qpZxMRy5qKJYVy1fgtH/H4vX
DQqff5dM6zOiCI2qALQNd45SAQ8su/YeMQ0eexoGwKR3p6lmIjURxXGAlnPpqUPtnjIPmaIb6LKz
/WbJTuNxyy1Ss1Ta3XcFdtEp0qMEjwn+z6l0fFSLmwlcX+zcVv4xK8jQAm2cwZU5bSVjeu3CNMWW
Txj6zKMkM7u+hPn6bVdn+/1VUDht0jhfwXLwUNALL79lj10QkXQJOeXnxtAV2M6sGSU9Y80mm6KV
Aj8SYTHgJ0YSW5lKvdgSN1G58lL/rYyAmNKz2v1ZPFGMlQrmoU561JI7p7GTgfx3BldYrF4VBki+
swnz6NySanotykL6jikI8FP1rKGu2ZemExn1e6rxgdFu0FMHXAgZ+6hzKsq+Gti+PjXJ/fgiKqoF
KuHIW7G73Hd7/KzM5Lo2RuCL0btHBTPf4b7AdTEe5garK+fBDiX+zgxMnhJqf0uRj/waw0l2/lV4
PTYiG+S/8UO217KqHkrX3FpvE7l/xlaizdEQ6VnwAnYtdq7tVon04c1QrASi/wD+FVT1sazyWSJA
/o+7fyOLvcZ1qK6J2afztXNJrcMXu+JDRRO/igosSM2v2NS6jS99eMUKDQ87eK13pFTOMQOtuANI
7XmRNKyO2AFzUQ7UVWPDAJgdwTlBRXAeAMX9Yk6UkKhw1hfjSdksIylAeAmynRr8eGsbeMvuJcdh
NPAkAJF3MiLt8HI9fLQaq+VVDN05y6+xwyrqgsSELpYRnkHqGQzP45x0x0/CwNH8YAdkTEIlJa+8
IlNLJBOR583HBJM1R+rrYtxPg3xQ85fkj47JnA88Kyr+PtfyEEyqgC34Mga/tDQLlyv4GRE2VIyA
+UyDyVgJ2akeSPonuU7s6ChFZ8Bfl/LPZdT0hAzPCbgsROXLPXxavyd3n+cEc2VcKjdRI9wrD3Gs
otJ1bgZsatkhVTIa+Zg0MlBXSUuqBSIv7c3rNL0Of2OHG5GUFPacVHmKd9yV/O77pBA3IU2rhysM
ePzKYUvnhL9NAj03ice9Gnhr/t5sGEzTD001dAIwkLVoCDvSxjsS3/rYx8YtMfVMcg0gYoKNTv6a
Fhfvg2af6/RPgnqeIvxDur3uou5IyNaTUfx5KT5B+2UMfeCQ7MyFiJf/RU8sjqb8+SXiYIqXV+Q8
uWlTpTNTocPTTRVtjeS1KNDiq2+/tIp2YdbaUnbOPtvsVmYipj3959tvub/hpau+8dpEwcgdKo4x
MCRM2UtpgeSZXa0fVkfMSYbpZv4tT1nmPwjGBsWyyKsFYVycu+dhaju1sjh1CJon5gSZPmtSAySX
/e28h5UiS9Jk5x8wZPv9zJGXOnu2eeiA51hZegjZxH5MC39ct+OT2MFjA+cK6AmtCLiFxowRWrHw
4X53XETwOjFASxr83dKWmwXfBOlBckGEAhTAaEkjgJ7I6t7QTxXLMBsNDXHszbgyhA6OP+htH6Jb
V4epFlH/H6xQ1FIJLzInfFFuQk160UVQia0ersyZALPsTmPFu6Y/44DYlsim72cgOmZjX7MU1mT5
r5jdrcfy5WMalcgCEhwI2u//JFhMSsHgbxP5RaUvQmb1QfE2lvW+sU2I01bEmjVKW39LMDaRxkGb
j/vPi2AT5BcnaDUMEgm3FwUctFo64nlxHJk1dclBmfVXLdKca4PqeagqdnrZXerWajeXPj3JXugH
RG/HXLQvWu54uKrA4ZeJKJ2CcntPA1inHDF4R+iSKVbLfVELGXahej9A2/sKCLE2QlXqNFcB/h2F
qj/TIKcoATnIremoMMRrUh9+iaCyaqIo3oScFTMgEbL9Xv3d7uG1goMyI3J+sdcpX1FK0Qni5Xgg
uQJa88pdENGWTRsnC47GwbrlzB7TsiMYZFdVea366/9q7faYxqdTfELTx9MWnD1wdOy6nNUrN2N0
cLoX18fXm1pkqiR3heqF/97DG5pIdvPl0pNGeYrrz715HJXwbqYUp98RjvfDAPzZrZiEm3q+KV5V
R2HFzsJ/IzQ1EPCJlFdc6GtEBshXUPnjh/ku+3pJVnjAWvvwE7M7Hjh0lWKbJYuenRkD19coqwbG
lCiM83EPXbBve5Sa705fjBguaG8a8go53gWDXTJnN5LaP4QFT6DOcpBZV9j/aYmZN/Ke+QHrGB6q
u5JTMztj/FiKodIhSgp9PgGUHi8rqphhzqCnjtO9jbwYjxG9W/HvH2XBLqkC7RovUQ6xLVAunvkN
rHFoGL4MEF7ZGTh4G3eaQmvjKCjVh8EXYAfSM1n4kPzF/fiovxS/L4011sPQCooRvvTpcOUhBGjM
eU+vK7YGqlt9tuPgpUzQILlK8+NCSgpq08BWVIl+O1kAOgJA1H3I5hiOy5OuV1AhCfKYTbhKNaDw
4K8Sco9/AiFCKywJcFpGjfXTT17qAQt6AmAm1uo+CRQXrVYQyheMokHB5gpzUC0OSt4nXH+wno7r
Fm30SreKzLhtAnifcp1DYLqRGQM7CRT8WoO1ZetOYnoYvwUw6OHBw1cvzBYBiAI+bZERmoZLFJjK
CFXL2TZy310fuOILP7+m91vpHTQ9CMeHPKn73BwoZxKOvxBuFL8RkrMcGGU7cpqaoEIP7bGQkUcN
b7CAhud1zFvIws3vGmxZtjtEd3M/hTBWfD24dEqvRm86K1hQ9e6NAmH+MEMf9WscC+bj5EvHEFky
21vyi/PkPVs9XNkYRECbvggq7/0Jd2mglCnkpg4z++i0S+Zg8o0VoJjH/d88d6r2o5wjb2a6wDOZ
J8O5cK+/OmwPeis8+yngDg+HIKwjqP/4C0zA6NJi4JjjJX+R0cDPVKrGERQqDAR/bN68SVjXb5wa
SwMH2OgA7nvM3AoHCTRhWhm0mYm628JpVJjMsng/jYGoUM4M6eaTys8Yno0tzUSKT7In59j2uNuu
UAOeNwpcLos5ZamLIdu+TY+pIMk1iSOh+kWcfZB68o3HrWj8CHQgwc/1F6a5ttkR/s5GrsU42lAL
kVFbAuTL+yNwxZdl69JPCb9nGjk2vJznuzBljCqmm/dejREOp4e7TlW2JPCNBnxs81IfW8m20Kbf
apfmR9Co2ysaT/6ay3tMd1XTiiwsRJIeqt7xqxCDb32sMaeKr3oFNSwgWJHNVWWL/G6OMdPhHN3l
Z8ayll3oll0KLpjKrSqLX81lhn0uYKRSp2BYF4g/kt7Nj3NGhFFyLneTDqFWwXTzNYRoPO5fWXIW
eQK+B9mGiRNBjsOIVmoK5q3Lyafu6y3gpSN0gmIfTeYz/DgEEW/XdPQQ1rlrGUICtRd5fv/Y/Apz
l6YSDbNhc8VnOCQxqYp61VwgkM3qUY2kdGjR6hnPBNjE1rkkxJiCMM3UJXA7J5EmPi6sGHQFX4ug
32jM4018/w52Cu7VmCgNpMpKU7bcUW7MNAxv9XEzWoXPyCLBHEzF0pJlRlFlCKjp5W5vq6ThVfbH
ako2cRuMiHsKcdtfzuDDiL2RxMhaD3ep0hlnhkxNytqDRGcfaYMNmC16xk1ZnyimtALFWGteesoT
jLapNq7Qx1/HqFlQl5FPKHhtg/rYQ9UzWWrkC1u/cKUliih9Oo87YaY6PgThP/XN4rU5NLJ/AqNh
wFnyoYIDVs52D2CxMkf8QrTOEdAXuga/MfmU0QOJBvrralntrVLRKD2541ftscMhPrsJFMMY7f1V
tgaKbzUAl+b7QOqMcgMNbW8LMSq5cUb3gDoWyQqDXQTJ/GiiX3E0pT/TGeymVJvoJ2l5jJihb40Z
YQ4DetiBQ0Mrq6le2CcfVHIAJ8j1qgO1EU0O/FiC2Y1QccU/C17kI8SzxTlSPKcPjD9sY7nWBwYG
TxiXPGj8w2NgOmNzKjZ2r4dcgyokdITmGjVs6moW+ZwFLfh6RqlMARvONRE+WMg+I0OROTOgUCAA
1id7MrdsKfQ9/OS2vShaAE2U/5VsZRnn8FTi4IMuv/y48ye+9GdeFPmaFORQvqch7l5O+cmelZyX
pACPgybAhxOl8PJacPvRapvIE0zj73F1uNOSc9COivFDirx6GSgSdruD00tx9ddndAbFdEvRWLe9
eVEib74lWXXFplUxHpb2AxSzo2loG48Kb72cP7fDst60ukwaep0n/As2sk+h6C5esi/JS0NZgrbu
oLim0DkOy0zGWX0KrSKWPdeK32SzXKa8KopB11srBSofFjlr+kfb9IGBt0hHg74Zebrgly2yzSj7
MoeGOazd5hiwdQ2uQ307Sonc/rjlmNMmdJ6TtRuPcgJtqXFqftihF4vUSjY+amd4af7EL4SI/4ww
XUBeEJYvlcrzaAHd0WRg4RSeKQni/Pa46/P9N0M8FNhXuR0BiguVN/KGGf0WnMRmuCauoFIJnw7w
EybfRMujcPepQxDdK0sY94IMqRhxErxWKBtE00HAhYOdrgWEdG3pDrZqKEMmGz3YUhOaYGOxcwFv
OCeohN1km1VGpl8jINi1lYPiiXkEoQhTBz0ZPpXbDmq0hbvoyHAFxigQr8B3p28ltyr1a8T286Vs
GszzD0gZOv4mcADlzVky95Asa7bX15IFKVIUeYnosxnsPvlJfUY2aML/Z0IEm6C3DwsWLMjW3G+5
aM15TDKGSyhbd6ZXqK2qE6MjC6943buEyJtlv7NOfuYQ14bLraQRBBAtag2kABJoZQkWgvNdYBAX
GS6kd/WrDN/gTX+0LaNMq527/+TQRWRNPiNU+r6GDKJblOFexapRqHH6EKcmrDzp9YtVjY6HHfVh
DDHRTwByrF4v/ahQKJiMYq3bz3ISIKSSqJXBkKIAMlR62UzpmxQinqhZDOj1ggbB07ACIK659I84
5qOM1UgcKdx0sol/t+Pl3yqsb5KXvV/hNDql13Objjd5ErxpQqT54R16HmEUzaglD5znUsNsGoqq
z5kZbE7EueKRZfexrtMX2pgQsDAoeIcUlHPiWRNO9R+e6pHM1L8UuXz+ycMDoQl7b/ZvVt9YtbYg
vmhkb/CseMIGqbZCpLAxXGQRivwPnqj0J+Oon3zgUHa/F3I0RbJxBho0usKsaqJSJpzK/fl7Wq+H
rwzbEhcuJtZ9qROBg6elqhciA9bzrJHGU3iMYXwnGvuxCjFH9n9PlsZNHdoD1r0W509HJbmNmULe
v5laiLyn1Yg3WYR6weX4nLYZKvOZTZKdOSOUotq32oYqVGhyrO89kLYaYYvfX1AZwLLclbzh753O
//GAweCUmHKkeJ1jR3PUXbLFTCrW7z99bFyDfyGQpXFlLHBlCNtK0+actgvGkt4RPGjA50qY/uiJ
RIOIpPUv6XoK6WPOeGh/6c9HRxULHgcoEhlI62XkEGhQvA8ZO8Sk3u7J6DUathvvMGy47I4WKkL/
6yfBS0eR8C4lJ5jdPEYmniJGBq7BwMk4o3c+N1i7SJQ3u66w9bLfZq7f6VwzM93udprUZlILfw8J
mw0qeXgJHB/6Y0R0OtQCskk+ghnCTlbFKEbEUuMsn0G0SVUhE7YF+DJacZSgyoEr/Qf7fH32ME1/
OuYwYKQMfdGhvQ2iCHZGGfX1+cnNX8CaiQRx8D46aRR1U7HL4uZ/dprIesaRf5bLu+y90TapH5iv
i6uJ1AUOn6qeLtscaveLv/3VoMrfRWhVJkzF0Bxdeh96+xv4g1LT25XY7ygw6pxonFCOmULqzAwG
5dGqHK9IFojTIZ6qZh6wZ8hL5v+neLBWbwV62WSQRAfBZUGBMUbD25vPzTPlWNcP9DSO2XM1zVAz
Ls023Z99AMfbMGjqgWnZs6Q5PjbmVBNZFz3DlIwwhAK5Jl4SY0FtvtXx50NCrkOcvZgmt9AdiQoc
WB6Xbx3Wg0iXbE6VHfW3d4dPpOpWeGzY4lMpWtjj9OzKPgYJkD3V85ikRFnPJvMJV7hTlv3BJwCx
I6d5MAcz56CEhreVsxJiTbo6GgbS/3YNDstT3s8d5HZTfOllQNp6LKjo/YjTKYtqPHgbuZcpiIoY
QJCzslgTOffNMlHdnXHAon7LKX0NIqnZEbXlkEc0SdwqH5qg5Dc//foTZpjFKiPrIXUZeCZGaBYu
rH8u2DSknOzivJJhXS4FJwp9m47LH8lygb5Vh4RqRVkE8hujb6bYPFejuVi1WN1c+L4sBaPTyhz9
UuJPs5qa5bphcjYberEqOuZf7QhvMybEzrw4juSZDvvDsHI3IFFp47rrotjrCp6lee+YmxSBGntj
LRh1I2GsSrIeY/6LNFhkzJx9wNhNyF2zcSoZMYvuGueIyEwMULJXTvjv2jV6BCBB9/M9moksjZ0v
0rwmeRMTcxb0gd2BBJqnSmjmlszqm3Ys+Fvjjr5IadsNKL2Sg2r8NgokmpKWu4ax5HouOOX7Tjy2
25CTBl0MnEIT9Lb12y+lvEPE1ygbc+63+udqxCy7KyDOvyla/pC5EcNSh7FUKJQxxE6pUzE7uCYd
wgwhTd5NO5DkqadbeTMGG3ZGpfoF6IULfnXR8sSd50cDBbeSj77JNc1IeaRgrmMjzblwarRVq/uZ
IqM237cZQ17I4oBCFhBy1lsBsalwKOUCY2FupWu+ypfgXRo8S9JfI92Yk6BtQ5GX8R//R8I+yVY4
enzZhc4VvDjrjDzVnkCJLf4g3KwBL0te6bhqFAcnHXmm7k6XxPZPZH9YtwyQYdf5LXBk9nYfDc0c
cncQZ1HWwCcQqBZtm5BRaAZHCdqpPby8Jb8mgr6qIp2ggNQy9RFD+MnPr/UvmGhSBTvkDV2Mj+oe
MR4jMec0VCtV3Vi5e3s8ISmhjxtL1cLoh2orVB5QlI1vt5Idr5FwZ56k8FL6CCC76syJ4cX3GrNG
TfGKlY1J4Eqr6R0cc8oxQMudr8+UUKg9ZS9+0nS9uDkGJSVgefIqB9c/vsC4cfvOZOZ7hxFjG8cM
JBzLL1fxbQyPh+xZvoDn5BFymYtv2gBkF3x9EmV90PnSSEsTJ9iY8slcnNkluUMN8Q82x5NA57yk
OTuAKO/InVOKJd/VYpKN0fD9+u53TMigFC01eRcmsPPU/m7fEHiHvHtzL45a80+h9DPG15g/n8tX
IVoeqPGSB3mc6bxoMX1xv40dsGNXQSSrTu4nsPlacN3UfYVGOJkfDV0KcybrvLD27+prmaGFcYoG
Q2TdT4ERk/gmYhsuQPdLB/AH/DGSD/DipwmVlvFLWP32aFfNeYKSG8esaTXfaj21Fd/E78+A5Dda
1/DpqFg9FWkOTi9tUn1WBNfJP6LngPrwB7HwPIWb9EIK0ZpkLoX6DkTuKydPiRhdKONV3Nl55q4p
O6Va4lHthgK9eMUQykb3VBBBHxd2O/sqI3z3NQbZ9YZd4Sed9oVUrOs6xdx8gnnHsmW0R3Ab7rOP
88QRWukLPxYy3bTusQguPUp6vgCtyrJP2/LQ3bWKu5hZ+7J5uFl0XcTyG00B+u5e5ZF0hCqeCZOY
vImJsNTWi542WBBX8xV8pgT4Xq63V3k1xdTah4XuCC4He6wwjUqFbtMVOqx0449ylQ62kPgq+H2P
c9BFChh7BGvopadpkoY/Lhq9aYXfKO9tWHQpLHESb4jsEFpOdZFU6hr1JazqJBcYKBvTBGaVQclI
J6FosvpIN7tKc8zyH8sPtcdqG30LFgEff65d3J5AAXlxYTcW5C0LZ90f64kArb0HWcC28mS0PmNt
fMlbu5hTwHd5tn08FeFvmEsJh75AX8qV1XZ/4mcFbT4Kd2veM0C9bwM/0twsmEjcYiAcfzTv5a7T
C4Le/xiayj1uGEpalVyVf44fTxIAZh7tfnLeYr6yGAi7AMKQx1n8X3h1phbaSeyZaL/DdoyD8Y8T
qM5Ym4nQShM4MacokD2J9mCMklVAwQLReJvG4+Aw4eB9GzV7GL83oY1vKhMUezgSCLWEPTJ0q0vu
XDSm2wySur2RfJWR+K87FXKsGIZCpdzf63HWSY2XFO9qfmmdugm30b1TiMr4LlO8bwEN202Mhbzn
/IvI6lWYpcL77Cqpyv9tNsGCDTm4S58D4Ojd6P9fRZJRAl8e+zfV314ZVK+tImEJiSi4o7dwZTIo
qucI4SRTf8ON0y5xFaRwGahsI/0Xoj41TZ1nPRYn/nCpsoelcfiZG2JyW/ufhXSUxo58RpQx1xOz
1r2OSdlbxKiehj9taSO7xYPKqU+BqnDM1Q2maj/jmnn3lK8VXy8mPTNKE05WunSLILmfhnhI3XBd
uOQzl2xaNx3GyVaJPrG0U4ynR0RxR6ftw7zceYZZ/YGouYcf8KA7op42gKZLSaoICncP79FAv/Fe
gvB3+HopL8cxApR3099vvaQu2xiwPf/ORI7vUHuOHlLyktKF3f8tno6enuIXCdsjF57FyNxe9Ssr
5st8jVN9jyJRjsgv72PGBm6zaml+o4znnvAnvREDQ6DB7US8L6utcBQo0xYVqwSxk3mon0GJa1Li
Su2/RveWaeKh35gvpz3NZU6qG81BnpW4XX4fb4tY9pQ0QlM1RJnfiN70ykutYoTzd0El0LmTM2Ci
dH5OpnYOiHrUt19vJ8kmtQDq/HACrLO7Vqzo/4q0ge/EJX2bGxeSKrk/xe/hK+KA16oyAz/ccvwb
4IHF6146I1n5bCHsxfuXT9s8FNs0d/pzSjyExYQ8RKEubcUschjnvc0T6N8GTaVX9Q0dMwwgTyuT
/OMJxY4MmrUqZd5/sBXt9b9WPp2yuhkeJulR2k5xGZ9MMqzDEyqz0atd0q7CmJKqN5XrXNUI8sUl
34m9aVV8Yxs3V9nYj86w+HawsG6SDzVM/vUu+3XDn54Z5KO9E7kDougUqxiC5wZBPHe5VBtzpKKO
FL41CFu9J0Ohg6dl5njWass0QITCotXqwdNvA93Itj/vJknV53z23SEh1StJjWblH1RJrsWUfsc+
EzbxO/X0GXcbX50S3RUlsnG5xzqJD52SZ5Ti/wggSxyZ/zz0ZaZwpRhfUyhJkrCBDinxVLdMh39U
X710ftMIcLZyMSmm3W/dD1SR5pcGAq6jmU4h1MtgNMCs23kbJ/XWv832A37gLMw7XBBQBPRWIxrb
feNu0JmDhl2Rp2c3oiurMf7zsRe3g1s2sClITuf5q543VQZTNCixNamB5Jny71G/M1CToGZ+/whm
pfx8XKUuvUd7kg51NnCZVIdkPrdVcEeSZ3h1FPAFpmnX/v1gC8aHboHEKmdoPeYagFSUPkB21dG6
YlOsjkyRvY+d+UHWluQdkaFrsLlKmp56Ar0qXA5IeHjs2hRsD/VoTxp75CiwijpVRlWW/6JOdpKO
wYZKp3V0KeSDcgWCxsva5rkwnYlNdgKA+CQRSoxV7+l/eUSxbU+zpTzUPVWr/ysAC4k5DwjleaHM
/B7Ckykh36WAS/mXUvW46eYmlNoQRMmjFSTVFQJY9Hyrpc70/dqZqMEWAelnA1Fq9sRydF1r2cWt
4Ep0Z7MaqRlBbu5PjAGKU3khDlujU3bmDD/PzzbE+7i1snS4t7cn97LTg8nJdTDlNl/zquajH9j/
IaM0bM4g8CGgPXXrIgXXk0S0OglRr0zNHVxdga/admvYPGehwqbZXE1q/a8fAhcnFpnpvdzPYw2o
yVz0AOCahNc0HhkhQitaVGG7a/X67GBZVrATZoju6sG9hXBdCQny+UVBsQdEeFhDJNKYE79TTeAm
3pU0ttPUvldCyNHt/Tv72qBsXmV3hkEum1/n6Xu6xUDIc+VDJ/6h8+w+e8tm0qIegasMMCxbH3YI
7kSz3fQ6YPog4g6fC1XBfHcuT8fkbp/Vl/QzfOHX7v4VeXoKC4keg4quJy5DSNO/2NQ8AE8DVVJz
OJP/RrtFVtzP6NgQuuWYoV8CtMtf5FmkSsjOJTL9rt/UPDyORuJ+BgLxgs0d5qAEDwTNJ0kk9S7h
7WIdQDUFrFYO7duQy4APhBNrHU4vTsovkVRzIz3tGtKHg/gmRcAzMTRScRCs1yCSeQgOe/dRFW3o
LNLTDUieu8Xi6pn8r8NrirlkeEbInRuo8jDeTBI/q1R/jSszuMo2OMo/I8cdqvXhNqvWW68XKlwz
jXzsgByNyuHl33WmxKw3wUB729Xg+3nqTJjWd6UC6vBXWMiab/cGrd63rnNdObT5JlcT0g4vhhmu
KvuY2NhNTgElYvstgcS0+GRsVlbHGenoNjh976FIDYW0FsgjX5hb+Xxc++sXkbmKyGQ0C9/OI6tD
bpBJzzZvywNt/EYzYbihdTka3YoXy75zEoVC8eNdQCgie7rJpLhMuuq0bHw7oDIQ9cuxtIPJEi3H
YMfQhvaj9QZAS8aX/P4WnrBYeulJP4e+kM0r0PUnAR02DcURmPfHEPL4m7FDgYg+EOjwM47Tt/Yv
mHp1oxSshqM+gIAhluCujkNIcHPzbnA6h0G0GXVjwuSKRO3Z0bRPD/ZgBhoWKJLZEe/4bJAPkoy3
H8WJJexcBUyd5Llm8mVnfGiSekh6xjtwcdfygfWaO4B6Kmu4i8sZ+/yTL710SMMyg5a/l49DwZcp
D3ahBDfz/IzSVEjeCUUbPtIHgryZfYySxAij+qZQSAssHmP7w5wSJMTAMjEOs1k1coi2AjxDQPfB
WUb4erlmzMa1MYF25gUt5jythHjVRk5fBZjnf9SQict8B0SmtfeKg87DoyOdzs6bgpB2J8l1x8iZ
h+hEF9QeGciQmFqbTFvjhOirTBvidN8Qa5UDfFe6D+Y/yxA6KR+a1RYmFk/dbQfldOhbL3cJs3au
o/hkbHAf9bNq3YIu8UiE+Kc98f0dyKmMgfTStNMr/k9UnKhElwAUZvJLYA7r0JaKJWAW1YS2kioH
M+PBCzRuTl5XG3nM9Pxf1GKFJ35li4HWlrA671JjFoq6rYCT0+ULsFZ1HP7uukDLTX37CJycSGYZ
Sh2PC0d8xfsuSfyAC5LAtVTuzoqXVTvguLxd3t3vYc3WOby1CEIhdoOFHRNukUe0Wq1sEF0zHF0T
sXrztat2GMmdMu51ilER5pvER9yJuMIz8bDB0W9i0OtYU5CsOgcu0VhXutjNEtBgiOmOGfmu4u/b
U2G5Ybt4w2yZaY3TRm1k1i5kudcohZJeQa2YFCM8r5krX4NTAGcn7G5fJGAuIc96N9KNI/Asr7nI
uMadUkiLkXsr0w2tknQ3+X5oZAzI7gi87Mdk0GTHfLvmGOtblObNmpTMBcDjCueDY5S/+FXa+FJt
B9YI+6/eeh7hakzN4ZFQ+Lv22lxfcZt+AeJtJVZtrOs7S27IAleT6TIxUu4Rb+pwQpqkHiOCV9hv
JRt2NT0qafEFEOAiZUUiUBB/KsctkqPXFLHEP19LqTV2QNMfGXliKoy1upAFeANwc65/ZCSwypYZ
VNSj1a2KZrot5w4wVYcwMK5W+0Qm0FbLip4wJnEA3fskNP1KBRVGerhNl0ZiciGUkrEyAgTY6Nlx
fxcCoOBmKgLria/GUOXBmSGcWq+XZN0lo2rYHN20gxmVVbzmn58t+4US77HgFD14MGsnrvRcB6xS
v09+eeGFesEwB7XwTmiKbWRW527FpE5iV+bObAfMyJxVi20HsE0XP1WBftsW31sxHKOcgLBaVzbX
9Dcpg1RLReo/N9hn0eOAohu8CvjL4JczYSkUeXsukjaRyNRU/LMRLITBZ1r/C18znGVnEmYoBaOZ
Ob57Lvqe5/Pn5QoXxqRp/hdleL0uFNDy9Wi7PMfPWSD1rXDSQQEMAc6arUgWXhCjNVo2MAi5P4ah
/ui+fdgMXmFYlTDXfXXxDqsTdzDs9AQhs2CEO7XuiYoTiMnR6kNu52qTW19lY98E3bYaZ7REi80d
Txb8dRBhaZKKc/Seke3WZbptCJTRBR1nDO4zO339yIztyIpoF1wVQZwzqKkP31YLif4pNqWJoEiK
hnxDhYC5iUtgZPdMLz/HNaG0J69We71UJ1q/dHRIgZy6uVfCIY663//hujYktFz/oGbmAnWlWg5Z
X2oq/zU56YUt8KQeS8+I/e0fJhVGwTqd19q3mSG9Co72afQmtCyUSBU7K8y+u7owYydkUK4cl4MF
U+8RuQnrz29gtgrzSBQ8xhqi8MKaOpuG0l6JqFIoVAA1pYuWBnudX0sVoO1jTfUc+uQJRVQInZuV
L8yeqde/Z//iRlN1DhWGidV7fSdLe5/+IJQ+SaT2oT6DYlvwK3n+BS/WY1tYJ0g0fdooBycpyK2v
qT9vj+XFdCu/TwJ+spjzgI2tyiejcYtycD9ymO3WYYaI51ocu3d7eQNfgNb/RBZlG2/uunjkRr6x
eRsvntPIjrwZPZEkKTo4atwRVpbuGSZadec48VM5O/FJx0EUvfgWfr3WRD07RbYK6stRMH99jejm
KwjZAFo32e6Vi8QLvq6ATlJzxtkGJ+1o3QB6lVTxb9pynTt0g+G1tTJjYMOl83soVmrvTtNhHYYv
ssnCQByubWLeizbanIWyjYp0n70EA8uiEI1FNfoAD8Yrprsm8edy6VONzQArWDgzgMRGD55dKhMH
N1K8jJPoWLEs/HE0DTCXGIw/hVLXW4ac9Rcm4K+WIa9d0IifmhjbPPcddGYf9MvG65zfmriy5gc5
hu9NWGDN8VmdY6nB5sbZkQMSRqNUstNrOzb4QVnLdZLLp88F0UeXtPGm3wVWO1fYAGasNUQNt7Kq
Q8QzbOBI/vUIDFUtCqZsdIiJWosiaINNc7jjab8rSpp1wa8DzEHYrLEljE1Y2PkkJg4AthcPlz4u
6bUFRsY1viYdZP59DRDxx+lRuxvT1oBQVYg3kvz9z4q43RTl1VkmWAJOzxIs+QAvO4GLzXLOYOCN
6IfiFHQyA3o11pjv8ZQpodRPjRy57YP15Q4odSPTcVKEzx3nh1kiX3l6f3ZmVTcOhf2dLI+bbWLh
ovpuljjmiHbVUJBNM8VVcPwJieTQbuu0Wc3T/mulOPlF207MziWM4kGgEZYOqQzjO1TaZt06wnSj
kNa+TkIdw+Ci3GPtN1guSmT9/c7pNzeagiEjdUuYQ7YaHBV5D0xf4WmhWiirONpCnJRBrnjox6Iq
TSFjfrybt3GXBqgQZfuqcMG/rmAmL6CFT6OcU+CwNIIRmWyCqReIGyPaiITgmLjufRMRVu34/rYF
SPeTU+9H8iOacIb0lOC9mkSB/TTQe3Md/pQJAZ/p0LgcmssvSbbrbuuJoLvE5luIj0BEGuWcFZP9
MXjMUBhq6bTIv+LJfDxIkGeIJaIfLuz37k5vUrxgR4Oq+AChvy1HWTsi9CLaVU0sdrcElDTXZub6
jsQaCsmKlXFL/3dnq2W54ay1XVb76o8R6N0CqtuqUAIFoAlciqFbiC2vtHtZQDWDau0Fg13PjQ6y
kC7mxHtL1lmzkC0OKTEAcCadSVNouArDlVf9jm4Glb3STVvpp0LM2o14gpKBMcXCjwZZywrFz73d
n4AaMkRVzB6NAZq83ZiiP6YBaq0RcL1hoX9tS/IjD55OAayfZuI8IxYQGNHdGZ/VIuVZ1CAX6Dvs
Y8II+WKJYHWdwOXMCeE2JyQtiQjUUAY3csrG13Ni8ozco3P0vgJQz1/KymHtEfB9PpTX0qgnc44m
CRMpKp9ElsCJokppZgkHriUDAUBZ6UzsaFEDU93MsrpBo/pmdBLf8wlguQ8tobh2YqiWq4qNBYXr
a4DTUhMwsCpskT+dg4JfNFNX8PX30UMK1McyZ4WurU+8dl1u1SjTASlIw+bvd9AhsjYeIlXeayHo
dyJhFruEHNkY26qkHtzyRlae7B3PeFIUdqMu/PDHPY6ZSM/RTRKp3qtki2ehX5seRslaieZbgiDu
dV6iUthOIECPm0pdNPVlxQ2GPCCiksunJ7HdRLJX6AYpFA6+iALS1v5Zuq9zduxVCzORgDZccQ2j
0+P7d9Wh9nZNrVeehV5ukQqp6r2MjWnzwQqSsG7N3Vk652jriJ7WHZltds/8QVLq9M6ZkXV8rSrm
VKxN7y/lgpFxQroGyC00ErYNvzPs0hHoZ5O9edNjlW0rW5n7nKmd8T24+gbj6AoqwVAladkFGua4
/dbXVQ6d186HnibpkxIvxRwT6vuWAA2JH61D7SAmANKwgAja2Rs0aFYdxbQn36J06Q7An8fYkePi
M+9RfCqE/VIquuthloczBZCgoS0rCbbBxgt4cSLRiKCYHxNgWHsJNA99QOhl0r+inyEFwDHMnabp
UUY7OD8OliNhSV2AZKN8m5wjKTyOuKLEM46a03Zyq15CGtdCsRt5d0uAgegRNBHtwarCVvGqOijn
scMEfk099v/n8bWjhU17QBrl91Q/CHod54qV9fREIB5V/GTfVDqtgFU7LXvEjZSwGJKjnZfQNIvP
4wo8Ateu3IlhpLZB6tOCKHnrBSHGF+kRm+ySt53KzrxVSMuRcgaNhna2iwPu+qd0gmSVGFinZb5u
f+Jay3QtL37f8V8yY2pFDCiFdjnlnOZK4LmvnP4gnQevKBrsb/lI6MqMihMzLeY4g8MEeqHtow2u
stXDagq8ieG24WolDDjRhxihC4VJbr7q1V9MZf1VpOBwim3wj38wVYujZX6pvKEclXie+aOYMVEX
AJBcwN3EofHbOlvDCEicIEaCNM049YJg9IUXWr6w+CBqWfyuNOXuhCn7Aak23CgfdBQfHjGPw9iZ
rPBHqW0+4+G6UL75jcLXAkZ+e536KBC1T5aFdUKNm/qJAO4++Wkl1wzP/wflGyeGbb8Tftzdel0a
qESFQF6YtoujQ6ueyCdvhEsPTecn08ul6OrUT1UxZhMMB8VXb7VgwXCT/VkEsm3BS37+7jxV2TQn
/xsMbNl6YuD4rJSxqr8DzYtht0GqrYKAd5c0l8KPU3XE/gxYWoD/rTb7Qu2BVtyX+5vBCIJGdjwV
1JJH7uq70ezoBe1WufyjPwF66gTmwawF0qe0u45wODajfl4S9ITbf4f4DuOfqbAuJ4x4nReDgCFh
8H868N5M1SOjtdpzO1XKmiBoSTSb1njGJagBFwxHwik4jbbYUf5rNm3cC1gItTfe+/3IICqtenOK
ECo/GOBb2YumzQg2EsTsUwvOMNaIR35YAEZyf38s+HA2LDxRjHAs0MTJ2MjpgP3s7GZxLkSPx1/A
mZkVk0DtOlcrOww1OTam236Kqmse1gWqJQLmBrPHOxE/2n07bm4tu/Pal4oAUUx2OxdwEJ2N1OA+
dfpBd1UtdN8IsamXud0Q9VWbd7J7vRU1M0ewiaacoG2h/FiiuaKKQrcH9aE6yyyNkB0UxKfyMClE
AUIzp5wIB6wIU9NOBUDSHispp8I0Rrs9F1PczFjldUmpaHzFDcHAjwRKHzy/xESPAhxHLmMuTluL
yERff3zWfRKtEEVg26cE2WqRNor/snCx859Jw+u2f1kRdDgjpigOnqjdwaTghBUMrokaMVJ6aDcu
BZ19Jt72qmof79kkPPF1Hv8wmndUmDCdHVbXQMaLYTlhYBMXPI0onjHHAm5D3C7XY5VchewOUpVd
pT6cCP3W5xVwFmRODOqQ6lusWCEV1TgTPDFTR+7gGKfvGom4XwwTDlAWITVp2+2euDba0DIKctJt
01ALec60YCxt1dIqOpVefgTgiu27k7nGMZFADZbp0vnJXFjD5gtt35S6mA2V5ynyfcUNCyHqL+PL
Jifr8SzkLaduzZFsa91WFMq2gO5+YA6IH07+6bWIFXKuam0XNWabgCTdcPGj9IfoSXpRlT+6UZI/
a7EQ1jQH0Gor3LC/rdIAwLY5NHxLq7MdXbBDx18k7N4bcn/dcHQ2m0WUeX5wcdNVAtjYj+EMGWG8
pYJ3SyDnNREWxyZy0ThkvtIjzJMKGipl/hjUdaEYRtGp6rTVTROmTyNi11mrM4X2NrBRVVdhYUlt
uuBbHXr68CqMGTakaQxsg0rmNF/9/CSFHtes3jlJzP1zoI2K8uV4nk8exp68+0MPqrzEaWe1FW7r
zxPRL6N+/gTweQ0ACKz7Z1OhdGHPyEmIz0C4Lg3AgA/pBvMkGaRaVbGvibkbnsVUlRVUqdkzb4nG
qwgzgMSqFIKyygvXcOGf4JDWea0OyNL29fj1wWx5WLfdIe7+YtcQn1dqUwTdwt8BGn83vbD41hnF
K/1nZbjdkL4xhQGF2ZIoSgyiD/HdojXb4jZg/7yfthX3UYfyqQoJVTCRbpz/gG6vwpaNJX0Bpn1M
Cl7KjiQFs8/wbZAHNYPGkc0hrs6tchnTZEh+4HO5bn2k4/NBXh2PaRJ7nT63Ipn+0JldUJBNsCsX
h2cov97e2emUjL/SNgy/e9Rr8FY5oPOdDwhWaeMEHlxkqXmzEUbzSkUAVGbF1FENcUVflnZpiQRv
GGZiCGydIcwhypP3wjHyQ/bP4ZepDNrFC5wQ88HwG4IfKD6Fo81c/+sxF2JC+3uIYWCQh7yvVGo1
6urz6BMEC1kRoQoDWiS3jsw9g9yaA2FXqMaAVBTKVVmuDXK/JltH30t3xx4Xtc49NykZm3hAdpqN
ZoAQhXKfP2qLiHb/2EQDfQsU4R1qZgFajvOlWiAZ+M7tvSM5VXG9Dan7mGtkqiyreJyUTaDboY66
gG6YRuhDev9V0gSZYUwr2yKBl2TtnVmqWQZdGkSlTGl1pD6A3DN8tfNx1IvUh94QapAo4WQIyIfA
H1DxxlukG1tZoTRlxZG9pDOYXZ4DoVbeXawew8KHCns6j5inZMiLFU7VNmrRkkEQ19p6MCZXJtqq
evSUhRNGVOg7PNFhQa7DutEBLh1rDQF0gzFGICRlQiwjuUjWUMj2EQQh3ZUhQMJBIUJYtJB33YaN
c7OhOqrt9sMWCdZnOL3Yd5bOELJ2dDw3KBiEJARnwLo+5NAD03mgnypyZpynMLd3RUmdSFBUgj+6
AzB9xOrLpQVA8H2BoqEYWKOuGdi5549MHFh8+MkB6rHFgHr6or2yL3ghowkmVyQpLyyJgXhC8ZnU
zM33Vh5QQYSae+jwwxeOHiby5kvR5OPNBSDtqISNCki1NVDt93v3/rkT3EFUMfA7orf7y+++axa7
gUn8Xh4zUq8lw7PBOmFCgR42dMjywcX/KexAa/3IK9zumhRTNchItqvFvfDqgNBf4lXfSXSG08qz
oVWavffQZTZWfhrMovW+mGh9aLQn6XUdjt7gxaOpgrLqFdeYUhviIjiOp8vSvcisWzagVklj9jJv
tUh5opdnkN5ntE/Q/lcXOHGwprd31kbYADmylmiRqfvzehq7UT+qVts1WYSpfZ18JZWn6dBrF19C
kFL5q7l//Jgvqso4/+Png6NgGT976DGANy0oi4UW87Hm0zFTlaxNozSzY8HPCDmE6gfzXTKuzkSx
Ss2pxZcH4q940uIYQMuh5FP6su/49KtVIMQJzsIlxPTiOzVG/LRVaLgbIanIvn8ElQdrVOVE4Mk0
RhAM5Z2vIt2x0IrAej+6QGNs31WL1RLE4FoTHQPFbweEVRLkHrKe/CC0amOD7v3/xqFD2ZX36M73
ZyqTPRLlbdoDyHkoKtFIBBNOYfYH36Zug2wTxSMH7UcGwc28rh8xoTo1UXYCUAGt6CQwSLpQfkEf
RqycaeLq2fe0tdhuKddX31iJZx8wg9XJFav4S3519fb5ndt2ltGHgG0jQn+hfcE6Iwfj4wuDuhHG
YYB9sA1/sZquBFaNQAWf6qkMcZVM05G7yZGBZZp+yV2k1EXxJTjaGKx2YGRQjK0q1vseJaQJTNFi
lOWUp2bEmjha2s0VcXeoz8nQJaHSpzf4XBO9Gen4X9z0rSxGt8Rz8LRhrUBntfzAnPTMbPl7LHpK
vTnbglgyYPVn81Ya8zXMr8ig0gFyNwopBRm7jJfG9g/Fk3CrvrmX0rWTnU3sDEwa2PFIXQseRv/5
PvVVgdnmb4DqV0kGS3YABrHNMnQ7ZUP874nsncyBiPK2Tn7a4KEouydSHxRKr2CzTdYSg4qMZxAs
ty+bGS3Uzv133ZjzqKjEzYqC9m46liMN4EKpi3cnIHjL7Fnu7+EQ89BKFNn+JOZTNvvFW9f0OXd7
xDg+p6iCEJbv6EHNRxAFPRG0XjYcjcJWO81/jgbfskbZVQhyFvPSnXMSm39osYubNXI2zGWXoMdG
MsokKibeVkRBjufIgVai1jrx0lUlPQzRJseCvp+ODL2Qj4lbucqvnpAbFM0tDoXNt5QvnseRl7O4
WZkKJ/t9qN7qVX/ciBkkMLsg85T2VJescujF3Wiczh3bpAD9HArrjD5Hjuz1ChNFWGsmmQii1CuE
UXtLroKkxGGmt4CWq01Snj7x+fFEoJiULcheaQSEcuLG5oTU1EHwnzFvC4sfngY2ohQsHzci8srK
FS31M5W1z08L4MoHWXQPgOml2yp8Gct9YRC6F77tcetK8LvV/cwTIJ8+JAMc3oONfAo7PRq7q1AA
8fueM+tDtHgJeyOGO+Hhvqk8elDLYEaISeD5reDbU3+6g8bX7QjHZ/GFLWWGMA1LVB38zPZLT01O
2XgSJ9i1trn0y3GZ+pZVJQHtuc0wMXLcm4ykEtXZ0A1bv4xN9xwTbBa++UELmxO+C/ZBWW/IxAvC
5qSRLyc7CwI+3Ha2hgn0fmiisG7MlCu6dLnR5DEbqiBeHGbbx1Kk5MR0l7WHtjedtbYjPo3Nzt9d
6LPj/twHhOHMy92HDR2p9UtWiOdEytRFjpA0ukG+1EsrI4FO4NS46aehfHZObUtCez6FzUYcDN5N
bOD7FNnAQII5jSF2MwBKVK+TwaAN4/LsGry6qIRUtYtazDFvpo04G2ea9EEtzWq14bN5o7wZcxC9
DrA9C9/k407/Lei48udVR1DoKBM3fQLlQRxgTUSFYsVD+RccIBTjalb4uv0/DohamKSeIB35LGLj
vITashNcn+LAIq8kpFZLKbLfjt0aauv+hzIZGQx9Wl0uhsH/9dgRQtC61RnZ2t481Mclu5l42nJw
TvLHC66zLN3AY5no5suMAtR4Aqt74teZLSidRd2fE8JvV1hWe5xj4zroUqNHd6YQ3zONjL9vHgqj
pm4K4GP260xvvQAZW9CyyJpJnk4s1U8akENasHfxTY0PGo0tVd7XHBgFA1uGC8OTrBCILn6gVlAe
AomYwSlyAnl0PcXUNe2Luqqi3NwgGKZqKyN9zfzPIBf5qoBHgx7Oz7p7rnmZVMA0DgyWAxqczCpo
UY9DxOVxMsQX8NJUaQ0Q/Ai7nxqlUD0THGaEZYSz+zuU2YNaWarkvc+RDu1bvCGvml2+b15D3Fm1
vp00AxkwUBSDFSVkDAkrPYEVYXCLC/8chuqlv5gxzvpA4Ztdmha9VZXjW92bJEpFySolCI/HtM+Q
gkqRHYL5CINZwqX92iMrRwyy6BbxnHBBsX5GRIlt6WAbXqyFhYHAubasj078bcnrPXHIbgFLu5RK
dCBr2z95/P8dw8UIaUYQuX6ex2slIoKM24T+/tyKBWBnAi3JzpoNdaHVpwDZ5791Wo6lGFQedhaE
1gNFeJ3Psk6NYElaGzPEuQzbET94nl7djysIrbcTA5Lsv1sZ/RWLJRxKev+ioVWXRKguTXOMU1dC
6CYlzWB9rloOaG8ajLrF3QCXqNY6wbienviZOGVIw3RYd4/Lfxb4pXU8ML22YcBoX/oUuyO39NIk
B5s4rrA57Yt0q+Mj/9xPf9e2/rFFimbtO54pOFMG2T6C/9JcS627LXZn845ZOXhKDtartNmeERKl
Bo56QZyG3ybfRlOtAxL+1QV9x06FWcO4E31skOWGlXcAwySX1qVOQTAmoPHqxnekX1cBsnu6tiHD
VUuIzKTx/fiUCpUXpnhF3XP7T30tiYWsHIfeGVgZOpFQW5edp48qmBGOnBtHMLYBWTBiFCe6cdg5
k/XeunIU7w+1g+n+aq39QTr0i8Am/753vX/1+n3O/r1yAQplj+yt05c+OTF1XnfgDNTGPZPBCzts
WrTiunyH3jENVi6rHvgh/PolgcdYOYj6VL78gYn/EKHTLCDx0KMyiimZ80vYvofm8F0bQKWNYVy6
TAsQ3KOKIrBT5WcDNIYN2cX16NBjYq5soYgwXgCI5iBO8FXS6YLhkrkkn1nB98v0A+U34rsTQ3pb
GNfR4x+FhgvBYPBGQGCkStxN1ilRoJznnxSks7OmZPVXK0xQipMpkzvIQasUtQXupeHSE9FlnXne
4coBUrR8tLesHt+YMYW4z90zPaBUwgKpyL+7P35HD6roRByePZPGSaysYJiE9DXYWyOaBihpAcFL
lQTcq4Hxi6NGxjyYgwG1m/yr73SBmqIz2XPbXplkzayirx9Qq74520hPFZbas5481cihB5Q2i1FR
K75kBOIIFzoOiMcIEeTgZ0fEFLE3qkQ2UbNHECk2mzSMH/7YUlm3aWYAAPZ8SCXXJA4buDh8l+xG
jZ6GSdOUjjwIegDdqQLMzIrhtq+9BQIT9UrOkaxgm1yCAfUOiXCPhwPRwVG4LAWfmCs2ip35pJ/q
nnAomIs0ZpR76FLeIQebsjlNYyxZyek0nMWJEloi6qD5pzRtPdUnjH3JrfJ6ovSojm1ESV6UiIbv
XfqD72t0n88Psty6EN2Z2mSaHbUWErORxvIe23vQYPuVO+G+FJ9sKL6BIK4u4//AL7N+mNWB07wk
c+X+KDGYsIs4W6fecV3Dv8+OR6Mv3lWaQETf8oyDyraHxbzXCeDtKQmNueS3UasZmNf/DsWU1Bs5
Q3iSyihpbEGo5fzzoFTDmwXXqDUKuP/eshSWk7QCEDrrmlqaVmtG4z7azqYQXk6vhP9MRZtqysca
m36JTqJ6+PjTXz6sDybCA4bhkq4co0mRE3ZdH3WSYaNgurh/EnanGOzYPM5Hw3xstgNWirfH4s6G
c8OMJVd4qH1nagsB3k/aRJ7BDfgSrml3N0re6GYRdfHFRzT+rASTyb7qd8uBMzL0olEDF0WVj7fe
HKW1U90N+Q8bZKOjo1hMY6JOAkFd5XbF7Bu0pDKZzWdvS9tY1qfkw+uGUDEobST44CPzeM//Sm0R
b3+6MSZiI8d5wr+UwFc1EziN5m421yXze0LHp53PLIu1cNaWvfDjy/cM1gMGTqeOmiyi87tjSgp/
TZmd4e9pQMXQhHVkfuxVFhB7cuIn6v13dV7pY6ubGBJ/NX/cWuO42WZCW27/dcbZTgg3P8qbhPiu
E5FvUH8+61o0QB4GxnOg4BNYYeChPr741p1tnsH7vCjsUd4dpDu2qYvCqFkb81qbpHevo560ZXi/
CdNv9BWFblgIjPUs4iDQpQEKgkU1nSUnT8TrYz5Juc8IRa7bkXbZql4+ymg1y8WSWHBUyuAdsc6S
N3XBs9Ilt2XfyHmd0D4gDbfsd2OBXAzCQw96+AWTSTI1C4EuFzt0vASY1Dmt35s+A9xWGxKM6tT3
frnGvcN9vHBqP+Qptv0j/9/fmsDN23Aosi4FOJvr/XrrBEPVDQxCnGhXdua6kwshA9K6iO85PiDi
GWkmV5xJSOwXiIT7BLelqFsnO1EObV299fIIcAqZ/5lM0nsbNcjXY3DRUzByBPbtlkw5ajLBA4DD
9txWA5O1pvWUayMDvlK4BSvuqzfa5VbpU8hxR230sz3Y8K4zJ7FF8jCBDrRrhy2YgW7yHle+1NnL
6vW7rZj4dAnwTY6nHRLIHJktQvBFho7It4ny7C3avPGKRvdkuS7akt8kVhFVzpu+Qfc6w9lAt+N6
Uc64xlalHHerF/FB920GsoxSgzi2DoSJGqaym1zKFoyS4Ku7WvjPJ2ExwNQG1/bhBu7TXubCmJC0
PMJjcPSB97QQzS6UgbphjB+ULu/ERzwTS4ry9pj6y0VTAorYTNFg8Cr3EMYWQgi25UaCxHUsGOtI
R+hSZezb+aJBSAYPEGNVS/YkcRyLOXahbCB2wfqyOzfCAcx4oCSV5teaLH6849fcOQw3rTJztntT
Eqa7ENabO+12H1zQWlGeC3gdSIe1KSX4eazQkS6/9C0fsLTtIRyj2MRlxo0SYUpdyo0AQcvG9erh
dSN2zDnuh7x4gsKS07jlc7OaTeS33yNIb2aGAtZgZU+CeU9cTI8aEGPhjsGCevJ0HtGtTDRS80wQ
Zf7rtNt42OEdxf6dHNUCBBT/cfDGpOdmL5xMU+53IjG4TFE3RLSyG4j9T+oxsbFK5pHhcKZHES6m
kPmJG+tg2jzetA+hSey0EZ6GzPXJFR0BYFedMPUjyT8FZVguGrMAG3IcyNOyPSHj/Hm2STQ5sMAP
TlhHbEiWsRqAAN+TNP9qYsfabqFMgvEHbM5uvDWmS2abpKpvriy4x0H4aacGQt3boeEXhOmk/Hx8
5/Lye0NqxTHW/Cw1c6OTgME6B1AcsMHK7CHl/C6jChIky/VFz1TzfMItWErdBJ5acU4lz9Qb/+0F
Kbirw5c5y8I8WHx1Pq6gsueUuBlAAzMlmA2P9wJRUxMwe4+GBjZ7lAlsrS2cR9oR1sglXvVR8NSb
tyC5ghWRkjGshi8AXQz2l61DPPbTbJAmgZeoqvIBsSqXA1SZIy/CWYumLDtY1u9spyGwT8mFI9Pl
UvB/T6oVw2nQwULpCgczfNDG3yu4U97CHTbHA5AfjVOhLg3/2XrQWjXfphatPEXONNwZsulPGfEC
q9TBC4cRpmxtSjNTp5U/Nlzzk1dox3CmPEQx89czQGtP1fo8v1825W38ql0gcaoKXDLS4mX8Y9Rl
TQlHSs/2lM5nNnxQJkuEWnKMXq9eKFRBl/HDoYtTfzwvv0HmjiJwHRMFEysS3AVrapzFT8mud5od
bJUjwUfL8Q7cP0Vo9BM3nC60vAI9pQMtQQmkptWDP5YpgmYUzDLVb9LcBTEZ0rulDXYCK4O1+n95
6LiPXpe5AISjScj2iU2uCRKDgdxZqeyz1f7obEkgtpKjB9ECuywgT82TYla6SgTrMzjVQKdQa2Id
C+8lQBjQfd3BLOKLgJ/4bdn1SWgTgRcDhlT+hxPh9UFCgyXviVXO/X0NFarC3MOp0m1hDr8n4hjq
j6Mw2HkACjzUjI/y6iaiL1/klC203cDnQNJV18pMqSqlX3h298vsr+w6LRyWn+pIpGYb9o2CMzCs
F7IhAnGJz0TWGC0Un2KCsau9EVYCi5b/9VI9PFOIDeYDZA1M5XdUq1dFZxGNuZ5/nzevR+RgwpvL
vpFY9kyPWrEQbUYbQj3G7D7DY04/7sbRVm84UEM8tGfb+9f0O/UmM1A4/wA6JstJ0mAebqTA/pyc
Dl+ZRuPGrnB/MHhMCu9tdn7yqD/yWNKvTgMa0ZJeqDsAvVJQyEXFs87JHnoks9fngFi7jjT7pnM0
XTInmEHlsK9a9S3udBjMeT3IfLV78iSwLv+FsrsWbgS8jGznJd8qu40kBSCV4YHNRTC8JOpxPh8w
wdDn+ASBedmTCvFkNzYgciLqzJQRubvGX8ZoIT/WV46rg4lezPG9ujawGPcoyWxwvSjD0rzlkUz2
yfK7gjD2nWWkmvtGwhWgmO+vvTG2W1rSlo++G5fh2h+vUAPonMV8SRRD8/RBQeg8P6p7WoD/HEyN
G62g2f7oUmqv7hv360jzrhfEULqMwYjlLJTOoXaHyvWBT8rBS3mZWfbwi4hPPjCVQVGL7ixhkVRn
lr8xVlL+3MtkvLdJ0X7eY5oyYz6bAlBstEknm8kb8mz81U1D9nbtHg83VcrA2iF1314N/fIALNyU
jbspqTm/x2tP5f6yIZH86m/z3eTl1Hj5oQUsq9tdVSh2GUrXK+1OjApdSnkCdF9d07elAPEX95NN
3DFIKX8LQNkvyYHbJUH/RHOe87TMD8zaPB+s67HAhK3X1i7Z233QiYsflwDZgrNwKNfx037ApFP3
jn8VR1+1zHy8FgBX3wCWc6o+saTIe1TRr4MzfbVVWvspB0DtaEXC65jTrKgepQGGLBikmB3Wme+b
aYqMP8+BYLwToft/Dgfp8tKtpd2rYvSdnZk/bF3X/uDyGNNosM5+GoeAplU6jdylreQKQFh/UPPB
e7U2Lh0Vvz+pnyTT1PxxUEdHH1TqlBGALFa6V86oA+vm4JlK1y0iLgLjAyQG9VWeHb2Un2SiXQHk
y7tibPVKqPzf2FLc92FuQe7WNIDvsTSYNSBJVKMu9oF3NR9bb5XVOYEL1bSe++MaWWrAmaqC65qs
jPfmMpf8/T1Ob8soIjQNqAqYaIBeNw5z78lUdFvvAbavtXwgeytitLrzg5KBiES60XMbTXAPnRQ/
UvRSayYXYECDWDKh3aBaHICbYne98BnfzXsprNRlJv7G3El1mE2VXpNCUiZzI8hWnLXV5h3C5q8u
GqGtUbqsL7SSBaSHIajDr6O56zv+Ijr49nnweeEZw9/7RUvvGFGPfUbfLQm4OuWM1sZsJMwxICgF
YTMgaUNdLZiKeSZLHfQPzeT0shyHx9C7DXPwNaS5i7OAyv2GxEElFk5qOxWERca00qNRpPOwdFYT
b0qfd/GfM8BnWQ28UOJmkJ5hN6zYVQip3GCneHvQVezTweNBFIKre0Jsn/XtWJky25hiJT9mjKTC
022P3zeNSAYbvlAYmkpxVhq9iT2llg1OOLZzYEDD82BPR5tyIVpGiur/RvpmD93WNI4P8Pvbfkwh
lhXdW9vMt7/0sRkI56ccv28buM1B1iTOgphEtKHOL47tazqyZI8kG6XEYgOK64L5Lon/wcBoX/DV
McjELAm8r5wrbw3tTLgr/CV1v/heDuY7mqdY6zkY0w+CVmI2qjXqo8+9uEBM9edosZ5XEdd5Sg6r
Z42i8lOfPxGq+Ylwu7RG2gbeiyrq7zDAInBllku2/pm0tzMBMV0ZC7h1bG+TK6ZH3DTl1mh3L8XJ
Tu7RvMEnIJEaHbeD9pVZ/9tGAr6tphv3BGgsvpxcF4MiK0na3GkFjngbQCurdHtISSkDk6LXF9PJ
e21yNF3RsahRoZOdFrE1ZJ7V26e8hbe3Q2Aq99HPb8s+G4nximkBjzQQZfECc40b1xpcnmknyh2G
1416gdvilKUq3pJGIlP3MU+13TD+5n98JKSrdVdbA/JcjCsd7XEImbwer1LW0fH3lFnuue6g3YWq
GVkkMe5dBiozD8ehUiYNtVUiBkVjEAUWuo+zz1IRZYgcmxSWuhum5x0pzB75VkF0CewEtl5MvI0J
QXQtINlSWC15MAZgI8ACsDoHsWMcKudAeUWopVUOeehAg7lGFqSOW77DHDKQ/s8toOHa0/63+eM4
GcZgxmppQ1FqAv4nx3yOfP1MOi7xQ6IjAqS7pL6YYvFNnUcFbxXFYBMoDcI2LEEcFWbPGu6x5X2Z
jExqQRsB7Vo/cLLKcC0kHgi9P9nEH2HWGR2CTVo8HUFRNkXUul0f25XmszBeHN3Lylak+8gQPDjq
+lf9aVOF4VfFdlczJyFQa23t2uG6AW29YYgBt3FNwmgyW/nPjaTDylGTSYLbLYk1a78OZiNNSEfg
1GbQDBTH1yqmL6SM9B0ExLKqCpMbLTXsUeHXOAuJpqVYg0MwmNrh+aUHyU9T0ymVqdU0GXqKzpvC
+QwsqkDijQv+Y7VR4kEMSFvIz4ybMkfPpzgyWwsrNYQdXiVkfrXRQBIWXOs1RLjCSGzxG332Lw9Y
oUn+TdaRQuuebw9mGU0+UNtjtHEkJSP5enwncNbxoHjAQdKNHG4aBhCV6WNnK2zrUIll/d2YHnn2
zjMM8FINa2bKPBP/Gdk3DKDJIOXtXcrxmx+ZdMD2qDh4wfjYALMbiHzYGuNL9vp6Fn8/PSp9ytfD
G0W22KmbFlV1PO5JwLaAK+oZJ4ilQVIe1H7v7HXipDIbqg2F4rLrgricC59N7nqbpkOk+MiofNHC
FGNIg+3JC1+LnJo3U9r2g55hIsIVqibeyzIk+FZBGaC0N0zQ6BVB0ljH/MEb78bP0Jm8ZhQLowBV
O/STHXBm6BQ1XKEOHcOX211O7sBq+TUb72PAMn/JPLi0wDMCp4hM2uPQJe3h3qeyI7dj4IvJOO63
0mXQAtIdAPEtBRdnoPwvmnMGYWyv5/xLHPa3ls8Ep6+bXLMwZ9bYI8UHM/z6WyUOc1vzgt/SH52E
80T27DlIjVb0/bAqGPqDtJ8g0VXGZcdVtMnJLsYF/MoOWVH/PoFoX4V17Cmmgl0oqXiSW2Nhmr1a
kMdq2S6TLKOSkEPl2px5aYI9fpMfmBN4G0Xkg/7FRKhLoQmrIz2aMcqJBIsZIk/aAEZBBZLAksh1
IA3WPkWjfhJwJvJ0kRHRQRt56nMRryLCqrlJW/zT56F1Tlfjk/4Ru/N275VtjL2QLUdTymlLR/kx
hLZlS1vBVunL2SiSfWHARC9n72j2rWPIQqXUBFZPzLL8gbQ1lMC+rWE7hSFxLOJMey2JK3m2AeG/
zWiIeZDrsUAiJ5/7/46zN0tJKc26By0orC/7eAOWmVclNw6ew7ylcKwPsGWCzl7fS4NilwCXwemQ
St081+YeTSuNB90Tu5TJ/QLrj2hhYp63bROMBEbMjcJUHZQWZNOVAYFdI+FufWewtNwt0PEWt0e8
/7wyC99biCiZZfkr16jCZgxqOOk06Ay6+Hl3497ws4+ThgJVG7dEYhc/kGy0XgbNVCh2aoi0LuD3
MuPQSWo+xU2FA/hO/hNq9wnEFTDmYe+t9ZYTGZkNQnw98flPVirjzAT7g+yY0mRmzsAmNgCdnuPt
/RGDazIJCCiYrR4cUfZd0s0QWye5TGdhOGShJDVRmgifDB7DGxGGHgdyu9EDHlXpSMCKtWgvkR/h
brACUoMB4skvY+tJweKNOLk0epCGZBdGU4T2AIoel1T5zpe+Gcn0JhlDbtnovLBjB90t7T/6J9ps
D7A9VsX997ass4durZzvFs7OShRO/fPXRuwCA0Mvlhp23K1920pmkDqHVV3b4pOiu/APpsSALOFN
kaK4h1Wun5bklc2hSzfIQsQx1FFcOBGkLwksk48YS+E3E0sstyqwCkHo52neVFM4rAacshonYDuP
n6tkn/iaPRl9iA034xAxqmtQvXrOWFInhZvtMGsUlmquSDhTIAQtJDZHNKLoIyXM0QMXkOGcY8IV
qzo+Z7+MXNnSJnF2rXZTFEC4F7KdXaHivCgofA5+a4zwcfg1naTLoAIz1ZCEZ+LoRdXi4FPTSSX8
FPCwvk6zT+nWIPNHZOK25eE/jxIPRR6L4b4K27T154G+Q9f5G+UcVMcCbLQDEmzHP/AcqhEFLxMx
bnB3GwIDdFhLdkRtp+O7a9tqgAZl4/bPhNaCFIWA5L9gRdmXK0bBcL/mxnezXf5ODHUlmMctun8m
qD2wDiwxoFyOISvB2BOMazzYv3jXywUiCC+F98SKTQM9VPNarNED6UEdW+dESavreav4KzSiXU/Z
2tYCJRZ1A25ElOhq8/F4E+bPucSYPh2h7msbluIsCH1bdxb0LeYrHvPtFDlgiPABjCVsVKEKRyJ0
Xqx3+IAB3x5Bc+KKFawihkOrNcYritKVf6Z3q3j20NjrIyPfdivyj/Z2gtkM77KyQHKed37Pekxy
zyhC3J0YtVYggolyKP7k/Qe+pq1kyZ9syjFoul8PlXXH3WTu2zssLytG+neUa0eMq7cvFDVBIic2
dw71qHEp0PGhs7tFIrHXly8BeTpB+lyq8aD/Q5rs1dnB+zPu683SPnKy2e6DGgZtncfi50m/oL6p
996dWTQnd70EKc9jpmihxc0Fy91u4KVK1ZfnBgnyf+maIF/PWbMvtY7XCUfIl3gHlo1CZXZeYCj/
TTaO7s4ZEecdoJycX+zl6SIVp3iVOug0zGN9Xdi2TfCxh74Cf6c773zTNd5v3W6b/CShmWTsdDPG
pc9JpCDbADFyJva9uh2WYcQaVTvlTPViUpRBiDV3/olbV6aDSMaq+ZLYwUYtf4YGHN/iTqMFLnFi
VI8q7iS4fa9xxShOnNYKb5pjTi5ESzf78IRdf/LZPfqo46zdSorABivjRvWkxzIWiALxM0PmQYUP
KiAmC9ZFD2LvVOOZgx+3DzYRDExjq+PVcuLEiKKbq83oOoVAENVt09AnwnxeWfx852BuMh/HLnMx
lg5rylOHZzZpvnpMJjzpE9JwDy8YUXRXUf+0uGScNo6Xf24j1dXRwHEB0aBTzi9HonaBL7dN4X7L
dkMA0J2TIxI8gKtG3zOOJsGTagM3sEzeiwlRCaDjFW1ZpM7XA9inKFoPnm2C3CsKiI7UMzk6gYsO
x6gj0lyr0NnPs0O7zSSdcTlDqoXgqw9RIhfCmjsXFCAEyw2EkXlfVdBCKoWFobNPM6E9Tzj2ieR6
wShfaNHr459k2h1po+LvcNEw78JCWweORSh5UmCv6ZUX+xOZq0ZhEC8FPt14IpRiaFrGrsdYtQN1
v7WyHeK/Ry8gQAyjWksXhO9Gx/HF+QOZaEkfLttoyXunk1J90bmkeL70ewbuwO26tdevvHmT3wlv
zJ8QWrt8hLYMOTLJ7M3TsnHOoKX3nMzW0i5EE5Uf/WNrY+oHihOpwONrDs/E7z64l5zVEBi5Q5g4
WVkYDK+EW2wRvZEN11DBUjMV9hg4nDhZsMkCeSDOK5suxvxPAclMzQ4O+A8fgtAchN/KP7F/ig9b
KMs4vE8Y/OQ0XbLoxXJtj3wTx/wAaAro5C15iTxD7Sdy2sXWAOyNAZGu9cZc6EK/rMD4iIgkgEQ1
CeKjAPpgoCaxcLmJYj8UmqdzJGBI7bAn4X3vpp1g+tSVztGZ0ufde9FbOYqUlM/W6M0PjDRTtkdk
yr01LTNct3z/txBwA/kDPV1I799HUIwvq8AQ6rAWxf/QPuvIsmY/u6CG3C8ig2QYDe09zAaDxcil
3eXIjKhAqe3Hizrv13CNHdbF8x3Z98uIhq5KOSCNYqkN/HmyhuEP2zDe8UP41ZoPS4ThKde0d0Z7
rH7YcH8EuDik+3ZVY6MhuTHvcY5FDigiS5/ktnjzq6oh37/YQkpZXFh0eqPVHqrHFul7PTq7a01K
uE3XdBfhWUCVyCW6djNspKMAiJT39mm8DP5n+MPVQyu4wKHenoy1q7WCZg/e8lCqJn4ABNQxtB8G
XHllFLZY2UVvSGeLmJCRDJuZuXWUUgWePwsWB6bEOaRWEZ+3WdtSRxnudX7Pja9yx8aH5xaBNtr1
oAlQAMOY1E9ZAfUxEahLCNjceClnlPAxgi53+K7ZzzNfvVM14ZxUx+q72ekAFWpgGvZzT95ogm+g
G0DODlEMPtRKxcu4l2iLiqxTL4q/GAAfDqXeRctyn4iC4FhWyX7GUEw/RvSTHrhstT7UyRgGeCN6
+f8Jy/csIO9ZBglYK8DDHKo1oGhoQqMARnrrTMOOxTzNbqCOCIDM5o73vMQNjGpqxtgmY1Xs/OXs
1RMiHqAYuNlhVY5Jupc2YdgLNxzIkAHimjqVq4g0Zws/YHIfS1ALkT/06hfRZq4B/m9jS99X+Yjd
66IAq9ctBcXaPJR/067fbFnvYcIATiD56sZQxOF/tLEtbNNUl4sLS60SVgczlrW7tcWZTXJacD+H
UFzDiDhhvkzfyh6PMu10zvbY3AAklt93twylvcqoQlIqlmEjUULIxdlxHiS5Ot8tMNyN2GwTi/+G
v3aMw0JRnn8iziFbfYvmM8E/snhGyYphbMibcP/1GxAbobb9Zf624SXKpc6WVJhxrPgq3AhDhoKQ
8FVNphs+jIHJ5yEnEG3UF5jSjL0WePJA1gGNwTeY5IRroAEjoB4nxYhvUX6hXtsOlm8oe+6a///q
vs8u14igux3ok6iaJHPChpxxtN4hkeKr9D0qIwJ1axlGCD7F1KNFSypCPgibQ/+djEm/hmDQM18q
5hf8EBSO3IK74oiMlnfwJsFAaxQ3d1d7QBicrCbFqEIn7NVhsSr6MzwzYMdVnUY17d7JIFTY3rNQ
c8bOpKasgb08PTLg6awRR4nFi2MYQMaLqkJbDWUBYGh1kVrHDpQJJHBMVmpsqOqPHxh9J94mSPYF
2noK5LHyAaVCiKdZ/tdG57TlRAKuB0jdhEvM2bP/7S2Gdri/leeUF1Ae0Y887nnZQSDlo0kQlRRv
3kst2eheJCz13OEfVOWbqZOhHI7jSbKe3aQjBY7JR0iAFPDoseFFkN69jMx5OMKplmNYtk+PPmwW
C1z96wkf2nPxL5W3p9S5+e/gn1ZrGi3tAOmm6O4bgqOxe8s/Tpg8KgxSfcAM1BKYTenQdFNdEE1d
1B78FLjqG+Gm/0nhrwuMcr8Yg4lEtS9Y7tzwL3jieGN+GwePwUsP8H87bU1lrMaUJr8oWRZfW5jU
KL4Bjq38vUNsFKLBnxVgW/tDeDSZZVk8tBNYxr3dwgbnRy5hHHoNri50QPrwXCC0SYUh9ebJj04e
TQ/kOsKqS9VyMLuuR7jhaNPw8SK/qJ03X7ZZFG9WaWCkjGkyjsH9CqYV8RFnONy4uyYNEnIs6x21
n4yREPTWxvnVnIkr44M/n8De6zxKYNTfxCggEhqQ/WkftbOZS8VPcuhj9mbAlc2xjsX5Rtkhqm4r
BV8Orl7Y28C5+xVBWa2nYNIMkBeXcVZsawCL9i15qFgpig3jmM71FOIT/PxyuAQZ/eg17m0P28rg
QKcwSwCQm3oW1UbBmqgWMRQNhpnYZ8Km4/bHIIuTd0oVShq6oNSTelKx8eCj7PXJlhH9WPfhSt+A
SXDOI8UM06sw947kGhMetTVMZd9h2+VBUt/Q7pSnuECz/PnGSa/ge2n0GBJTfbaCLOX2hj5ylgcM
n0jpzfGEbkHGO9MKjXa4v8oBRKC+Anrr4NSfjLGtX9NUB0VObktGACCGRj05Y0A2xMQ+ztAnH/qR
d+TYsR5gandsz2fA7wsQjShxyumyMh8yB67zTn3Z7d0jkyJfEPZkoSz8dmwII/QQX8bvB0rGLVMg
Z61GlOxYxJYwpu/dx6NvcTIVCoG5n1NcVkynElZr9zsMotnSpAl46YpJfSEMzpmi6+EfsWHK4noj
cPNd2BFHFwFYZolI8iGLaTS/IjLJ1bPm56HPt/9U05Fki8m1H/jlMzh7BX+sk9eU3hO7lnpBQ2Xd
ESz2CH0SD1ObTUF8Df4j20y4QUaA63vhlxqVIbMIeMoEAIJpqvZo4SyPzotBnRgpSPGnPuTX35NS
rDoZNDmIbRDR/BcYBJoT9P5udGwPbziYCGgCYeA1lc8RaWFiwmh8FPQJR/KuickoRttdzYMoiYER
dMr/qA8cegj33fq4fHqmBPY6q/AS/WTwzEW54LTx7gigqdcTLr4YYLkm0lK+UvZMqPd4eWkT3VmA
ZFlj+1uq3RljQ9NiI791NlkX+TghYuMohPwvzfhiRh9r9f5mHJWW+oUlBpunMZ0uR9FBrHiiwFYj
RM9szDBc7a2vQI7MI6JmKfz0cQ2d3gO3u6Xc2ZBoX2PS9E8+iFzZFt5ECjiL0MSqzUe74DOcnm56
uUGXGEXfCl9vj82FEv3bsFFcKLyWQi5a13MZLM4SnYKADVD0TW3T8B1LYjrEJCzVPU27KN6KCHFj
qHzaaW/EL5zIl3zMDKZhBAYpet2CmGCGHqgf4nU1LieWEnj0fw+VkSy8Rlw9QnsZZcr87TulqaB5
zXYZM2W1MylyyJo+0kRsn9By8Kf+lEakriluYPYhZn3dQgEUL5fLv4mNFHeN/jBOVVZ4XvYUNj6z
zGh9jqRgKvv+RkrUoBKb7msqUR1usMu3371sAtGElCoWsTNM10FOCbYhyig48DsEpaJkBJHH/wOl
8hfaUbnCaLTdGYueuDSq/Kyfgjxbw+qYE+Zs/Buwb/EQcH9PN88xj5zctMVF11+rmEdZ9Rbi44aL
zEnJZOS7On3kTm/Hl3f99hhppa4Hg5J7XaKJpBC8fFDQnAe7D6t5NWIszSsIKhzvP5f0H+pEOY9J
vbFdjJdtfCJnvBB3MUA3SsJNSl8OXy38/KiOUz4GQIS2DPGWK2H4qCkeWdiptRgMgTNJHVl/9j6W
lAI9VhbRhZ6Z9cjZ4hROdIMy5haQMXJJ5Eyh6NW17jD6iQ6f1Y2/BwATEluJOh7F8n6foFnhGlMG
xXl30FxT4aAHtSM6E0Hd2pfxI1yHZfoWuI3GTSRvEmZr1eUIBdSvQlIgbSlvXvyFATdF9kU4cF/J
mFPDsO2/Gv3Q/cc8ytAoiDBV8YVQ0uQUXxOYcxy99WIbbYziARyouRZlLsPXcL8x0CFqpUTb9Y6F
NrFPscP6Ckk6WTodYETPX0H4gPOMiBCqVmJLcCW8hRPB/xF7NrsodBhOsEgTN5p20Yyqbs61mOgP
MshdW3121oiA56aqAUitxbIJ7fnxWaUoAusF3Z7yn2VzS7/ydPHYIXGm+MRfdIK8YU9A5kYighZX
kHnAyqzTsSpmB/6g46HEStSjQUZC3c3C7bUynz/UX9CYxPM3/K0t6+0Qo0s7bAtgd1DLk5MK83fj
CTlAKyO+BjS17oVOsRnW5UqIARpIbXJ3UU1ecyehp+ryEnWF/M729F4W6WD4iTMhon4fuEHK5f4/
hJnxb0XtQ6+AdIAdOGYoatDXkGRott5dhFOvXGPeND4veKJ04Jbb2jW5fWGlGo118W7K0pvucwB2
jaL9Bi039yAkDnVRceUxj1HJWy9n0KvqUxwlCM+NcaZ3czQX285zgX0gkFPL+oJpz1h+GD93Fu1w
4RNrMt65DRZ31csGMhzDEfgArbTkvvW3HJntWb1EGYQ4S6t1ztXp1zp+70xzj90JWP7lYRHjnQ/g
aEF5PU+MP+53dhCNkQ5RmPkaPR3S8/1AtET+UKdvrS6FqlBVE3m+FPc5FabSERePkUnrBriEyX/F
OejVfVBFJ55k/jVx3u6hswIelixaYXXMZuCZr7S7AWSFpR3eljXIBoJ4hd2crysx162qfW6pl5eb
lOWYFNq9qjwd/aDChOLYvhUKmo5hoVpEKpwptczYmba1HQO1JZESiFuVp1Z+Bx7ZECcpIIkb+ODL
kDfk93PTvI89isURld7PgxzFuCWZ5xhFYieqH7/QBPodfFVJzgiHme+6kQPZKF0YuMkGzX/yoQKa
Spb/MiqL2GtuTQktVcZ7bLJ+9MBVOrAVs7fFqd2c+z0vrIl0AIX6tWgEAruXSrZPbz8YUw2twwP3
4gZLdhUfpaZQaYeQpSC26Jhp2cCTchaX7q2oOv7I2Tw/hxucmfkAyfNTjdIKO2dHkxbAxKxTaBj/
vxzPESjnuiXB+LxPACJGvfefmxh5frjs4yJ/sBxIHRzSxCtmkyLVktt567aesOaKMsOExfW+3U8l
trTfBDjf9shSXhePz0fRxYsqUX5A72EnoLAq6LTxD0iT1ComARWnU3vgnHV8urtAVmXaeZcbCh4c
1ej7+PXz+BKq7ZQPOivjkTm56YlQwlTTrcv6DPOReRod9CgW0KGwqt49ghT3GJhrHUki4LKjiwwy
w8si3wPv0CdLYKiZYylka63lZ6sCtZ1BF1PlthP9Q23hkq0DLqitvT0z1vPUucQSasep0sT6TyFd
kIuJMb67EhpluRV4tG9InDlkFPEkFLNuo2l7iobt4Zqgdsv9wAYwIZPZN4aiEvcAhoLr0o8FpE0c
3SDIh7SBud6REA4fWzKFeu4tcrM1FfvZWRnkCFGEcjRsceUec7ZOCqjEvMGGVvZzHYvuO1brvuiY
C4TJgqtXIz4tDhg414aoPe/0wLqkWjXPyTt4u4mXY0PP9k99CzS2w2Hs3aqkaaI8zHLb4wpYpvFB
kI35TNSKIib5YT+3hwv9oEfPgyZuV58fSm5xiPt/XrcO9QDk4T8K1QHj6HPhrUb1Vj8VI3lydjP6
Ng9t8e73MikK5D6amxRkrbT7WZE38hL9IzbnPmGVhznMLXn5KfneSYY7cals28/WFCyLZukVlrOr
ChT7rzaCw/Iq1KSOlv2xdoRkRZmN/+uPP5EzPUNfGKjr2EKKngtjV+rUGfRz9j5YB2KkA8tuEfte
9Bej7TOPY87uQciddKjTI77IimslwkPASfkZdLmIArFID9wHU6qs8wZ8ENfax/tY1KnJFpWDrGt5
Wm700FMu8B16EHSISi1LofQYQVDdLW3gLhiGZqWp7zwKKsD2Qu7P9lzyyRHObtB4vdvvi/ZsziyD
EHsUfIIgrwZkUJgIEael5pHfr4SyVdPbTZXToV+J5jwUjjP1tpj8gEAIK2amiiaNod6SkNuEntPt
rRX5VKccIKkL9l2jir084fYkIw+l8a0PsQpncjuyLqDTNuvqUP//Jd0idrLKtU3yvcpwommzutgo
u+j7XAh9jfnnv6DiEG5IWIRhfQmb4N2ZCfAvgqOee5Ld+/8wFrircmD2If6Gqam1i4vI6+PO5xHg
LqeoiTzDpICoFQjF2GEQcCz9MUgiBKUmTqIBck7AVm57mIpmZt78cS7PEbI4OwwenEn6l69P/wJ6
fPfDBDZkJKlvNtv83n9jGFys0imJnKGJqoqbKX8NczZEXPgMmoVNLSMzSqWFojpJGjJNF6C5ly+L
7TPODJNkD2PkSlX08Sh9+dYlPCDQmq9qNupBifMi1LsSFKVGdkMdZuAtsiTSEq/qQfZJTAbtXnAH
qOPh25bOOSGoRtbRGBL0zaUwZcWL97ZBihCUhaN8AGp56YPQn07yekSsJw4jbXh4G9uapUHUnCKW
T/deLCfmITe1Crj3sNqXXoJh2C8jtVsYbcCzVH5UlWvj30CWR6ZUURKTu8Z9IYpD+JLpwGmsd9FE
0g54TFtvcbQ+1ndXDcfvY9p03vzsORKldY8GhbNYTnLbfAOmQ4MXgYCj7VKHg63ITq0QBh9hzog3
D7d4AuKzF/BuT8Use0FeiO2r4yaeAQYd48V2kMPF6unluKctzm8jM03Rj4cr+moWsW3tc/4JbT8T
7UNJ7ZiagVC0eAkxb39ktDVixTIyN5uRay/c7xcrtD57pWtioXd7Qy9li6giQhlD7qnrMsRD+YBK
brbjlZ/dMds7ewZd0pr7P+6qaDUe1Udebh797YBTLWaILoL+nAh7XEnBODgWoNIjYffmYnaGGNcF
yVAB+Ob5wVhVub3S5CsIB9wzBFDjDXu2Ax4ZbiZ+K6Pxla6llC/wZaEr8X2Q+Mh3TuqGOvvAJkJ8
iYEnQ0e6x1Tj3AWIa/qkysl+gXQ9NbAMrxL4oyMMqDDsMOmFXOrL5fwj57orUvZh8gJUyKOFP8Dc
qUMF1PfKPwyLXFdytXzs12kZVEAem4YjE0sZ+dR4+eW0u//iAEfHdeXFngo3D6PbTl8Gq5yIWLXJ
lRUuYpMcuIC1r0Wv8cn91nPpJtcqn1xA5al0eEErDJ0cfqhC1Hqgn0JUFykPcaqveVbnlAZd+H4z
YMImjoEl8ThmHVcJ+EZUuNHooHCmtMVJlAIYT12R5kCDqaQgOTHcXUVxbwjAslAaCaxXTgQaYgyF
mCZpxteMKaxa8autDmafW5TRzIs7UkRrx7XjSfRh5T3TLwFcWYCX8yH4sBNP5uCKdj1UCxBAkgWw
hGg4oDSjLjDeFpcLIEQw98PILt67Dtw7xYPaEjp5vtkLcCV8ohEDIUkck3qDnd1CXrhJRQ+xhilw
GC3JjDEDWsPhwyCK3y0XcJ+J/ZtrI7kJDXztmIIZf6d2GsEy39XDBgZ3AB2dCZ0+UrCvU/R04yaN
ytrFspZ4W8D4STCsWZ0k/075+L01LLfP8j77iYsjJ544vwWhFmCW9qrW/yC340e403eY7TmVgHSv
JTXBoIixharu7RfiMmQlM1Vjg50UiwWaXyVaNTTmJVLWqNiq8j4elwLTQIkFr7KwZQAywy+acDYO
00zvAE5k3UQe+9YuR6YI61cnv0C3eONnvKJINBd91hN1dNXe+HLm0E5mTKX3yC5q4+NmIdj4lgnQ
hr8LzNmSxHydoa8gtN7Whbsh1e7lqMp920yFnweTSaEfoiayA1qH6sbzXYcK+Qc17IZ8jPc7np8N
/uZzWHVJSf33KRwVX5W3uK2IsLjxrzdedplSCdBz75uCZi6CmGkTHNXynol5aTIbA9/KgrGUvpo4
XDIGM7r+PhPKjMIrmvvXzanIBmx4Z8vBtCePu4/jEYVsxk3Ks4eX//fwghZNp8vdXwpjbfSKMQVx
k/bu4RZkSUAEA2YLpscZVmUkuFz/xryFpZgsCFYrUV+b1TVjhcOPyidTltY/CLDvPK28/CHokyJI
xsSBL4vNhXV/yVoqopwUTKOKEeYAucaLHTpzNlBiwNKQR6gpcnQujFdrju98wouW5oh6yYu2ML+c
dSliA/pMJ1O2KPLIv4VhYH2HdFSAqLGZhx15qBPjzxDTBdWfkF2PVyrFHvzS6hnh6gRNs6phIbkg
lNAuGqzKb4t7xxF0izOuLzeyVKOxnvG+cq2SEEDGAwSajz6W98gWSgk9vVOg6sZ1de39EzGlRXjg
3tc4+uILW7As1F3hzKSjplOnFAsVJ9zm1xQ1Bl/FBL5NyPmCmuE/Cv9vzpt5/O97d+Q5ScMfYN4k
oxsNaNOxnMSrFOaqjYJBwSTsshTPFThPhbD4wQMrXUodtihpoSLsHkTXJu6hJO6bz3iOm/BmgKHH
s3ZlQFySss4/sPrFLtvjcektGaue9Lrmcm3iL4KVcZB0qdS2RtBsjax56LECmyz2oYy08yc+4G4p
DNKxUrKPuPX9sEu6rUgj+2LvhiEc/N9HgmkgfRc3pNeUI2ihf0uu2ZydBm1gy+zYviJFWFNSgcLf
bkaJEwE2gEJUCkJAodUXhvmxW7KC5QGQYm6vMKhgI6pB4VLJRkc/ciXuSyvj75BqF0HJpIs5nIq2
sr3J3VPZAI0oKisZJz1ksd/79EO5Zc3hEX7+mZ6BGWzYm/MUNF7C3DF9xe0yypbO9A+HNcIYmdSy
TIu1kBcJ5cKJyIkVvoVtV9c+sl4lA4ol6WwGkzaUkeBjp2RW/QRmBfjJ8cehDyLk+GIJp1DJ7Ly6
yH8cJ9IoGrzVfuKG9JK+EtyZ6G3FdNunQeQZUKuPLV4bzXX/vCrTKlrCKj0U9A5xm5tfB0Qr+9XA
GZdutnGh1H0Cri8op2mV+2EhpEyc3Oo6XjrG52ZKW7dV0VCevw3cja0e0jB3e/s1d+OERaGBhjsS
/bv/kwooTtXJ7YZ7ogslGWttTSemFbd1cfo1YYbLICRwJpxSprmbzQGtqC0rXajMwbt9C/5l5zaW
MCR5XGkf7EYbx3N8X82B1YYeSwSOZwDSTQw0JOPhmvIWlL54LZNxWPqbpeCToyUDmciMKMOC4ccG
m0dpgB6ic2WNrkR3tHrGQaLX8AQtzIyXBBCGcFYOUP3+yIsW6erdh7opgSBwIOOLg1/FXdxHJ7cV
RAVWfn31CJ+KW2k2a8tLdSz3LRR8tw4Ad5Ip5YrbVWGkxBQKJTzIuo2G1tVRwxmtueRMMFNbTHiW
7s1SR+reuMLjZzh1+ndLq1vCDapqCCTfq0kgtletvqh/dLJiF20RD0gT6dLBF6E1/4v8rAYiJHcW
9744Rj+6rZzTJIs0M90BkyKr+ySByEfbJfuQq5x6W02EADp4bWDSwA9YI7ZK3f6/dNULgKsBjWkX
8XJjII6tBtbTOmHW4puSWENyXaz9av/3XXNdccTEK+ZtgR8ubi8glpNX2CYNwpS7CvL2dHuql7hV
SWOalAhDJuw/HidSt5/Qo+stPw8gEHDQs0kRGDN3tcYvqOQ4sEk5ok/jg25oi93Edj7NMFFSwsE8
++dAwj9pBaGglSGFpX02IxAaZaUP7Ce9/d2R6WhlKNIHj7iL8KhNzsp6Rjr3cktAg2m91Rpjksc8
9ysnWGKvmlgTrcAUjR+pSHuLbWKxlsNqmqdL3IBW+8fFks/IeFLWKJH6aSe2dw/EVgj0R1hgMgjT
QTNOBcI7UaKjAjtNEsCPnmmX60dYB0PgM92jAtKb6B3DuSB2VriTXZYeimcqG/Zuw4b+vEYB6spc
trgNVjuRFQ12QQ4ank323CXuaqNbO5Ha5UMVeDszZjGW0zqpnk4S4BdLyVh3SXVTdZ5BN2LU3G9E
J8Ri98267QHwhnFruXel3fid4kVPCFY7FLoQix+9I4anZoNhcdzGbWn1WsZKBsCkuS8VoKQWcUYR
18fKBe64h2/7VaR82DD7u//ZioLs+bcn3M1nF5lcDJrayhn+7yB4PELbXDSqKptFBNhHorR9tC+W
e+nWZmQBljivYgtbDvMNQ39n9QGbfaeUG45k6KqiPB68zZx9Gqx1OJhUnWvuqdQk3ySpUoblZ47s
xsTORn6nSjl+VP5aqegQzYNdohYS9luktlvF2lZRSOHre+D5CVJywArS/un0p0A76I5PR/GLjN9X
PW0IM9nRoFOP/SEwtr9NpJiix4/A/UsoueMILnO7Ihfbv/Y0bAy9n8xMMWbJIe6uy1dxZ3sv0iKX
T+grmYfRjGCIYuIMVbbHkz13QqlYkSh28ZTvn+Klc0tVb3rhAViNWtAr69pWpgOaJM4KeUwTjAwh
c8hypM9unSHW+axARghHWe3xDhMlu26xrwtagp4LejQGdwvGrUMCPA6oP/B0C+U6xEuT0JN+l+W9
E7q59T4uijl2C4kfGRLnaYzB6wP0HQ4Wn60QHC94d3DqFjXi86k8wSMGFSK0Y4MVk9m+3UEs3NnQ
9p99DunTBQTeVKhOErpcGt5NIbjmk7TWWUeX/yvXI4jQOuhBQys5D9RE/E+y4aiseQM6qSFqNDRU
/KfevZq5hOOiOgDyKHLOt91569GQQpGDJoM18N2JyuHb4odX7n6hlw28AoHUP48AlceT8260H4om
Y2LNXpVgENEwEpGXrvGbd21uuZ/I1IiioOyxTGoI8NPS5InnSTXwS7y6lDOGuw/PaUolC6qMKElT
JuM+nKh7leI/oSH7MCW0unqffLlzY5qljzuJ9/EXOmVTScTq/H+5rOjZlN2kxejCpIrNrdKF6u3K
orMoWEbg0U6NI8SxYyYwO9WyLP1kPfqEIGQr1jO34GQxeCXCvIAgb/zuri2MFBj5B9h41NJJunjC
uYXtVR3G1rwU7HSZ/R97BHKvgPKmUjp4KfaSZjZUUgGHdXe98eI4GxaqVAdbZ6EGoOx73hlUfBjz
mk5dfqXPRVMxZAHNUv/0iYmwDk3YeEvqPLJhnS9tAxe2d5H1V2ZCtaA+1kJaOtto+aYxr3VshUnX
l7T0AaloELtkDPL5I08q3sMUlR60RGw5+ETcyvZ1ryqbCKElMg/uNl2V9VjI1ce9iNK/XL+dMzBS
9EIo9tNCulkARcX9AitGBvx3sTnFEmrLo7hgVgsed5H9ZOG1reJkdH0N2oBX0RiQ67WPKDrx9SMK
QyjiuEJamZWYA8KPnSkZJ1yuWg28lwe1V3jcplVcDpsOAlHyJ3LNJVgPutdb4Dmaa12lmSFGLGK5
oNak7Db7JZHcP4m+q/SVQss/sUFqO9lHZSpDqqn4DoNfYTZpG+rReqceW1ODQORkegZsNyFo9Rjx
c4G5syFIUyGrH0vk9CJ2DxUubwFd4TuiSjoraB4tZb9JqnqF012F2T5Tb9S0f4YUx0XQ8WFQtvTw
ytFo87LpwrRXISAVjClHzyjrA/LbdKh0OBfPJDE8soOiqdQ+lvG+fb2cmRYpPFCxGuUmpnfu3ME5
R8N80lKhuBWq9F4OXTZ1aIjSi0rlhoahqo7NSIOtBzxWKQ7l0SOxGi4AoVTfOgTW5VPhbW7vv9W9
rLNBxqD3zDjQDHGrxdiWfYie2JNbhp0bJu6YUiFNqXK9uzCluN0e0T7JPSQEBVg1kRpVb6VOd3kk
qq4/urN7BckxggXa+bsa6VkCLJXLPR9X0l0We2dkwoVdY/UvTokKKrkTsmValx6/58xIAkLzFlFT
t1+KdWwAWpqm+QuOPARlrbprBS+DG/HPXkgvzJfCS2Zhb1f8RGHuIsUKoFh2t1O+eCjTC3jbd8JA
FqzuWxBEzCW296NgKZ9vaG5kGcz9IrwJsjmnsalRaCUEmODz4ujEU5g3dUGWLo1zJNzFIY0MiK8o
37szX1UZP3x0iERjvEGGZBNLiqMzbA0XZ/CEg43OUnzqsZjxnPESId3CZtGMQSGtlQ7VQidr+Ny0
mH5lSLv/e6i2c3jSks8LAjBmxSMEEkv0grRpVfLixJPgQz93z0XdtK8WbCQUzCibhqF3nnNRlCAR
v4Qsz63mPdIgHghqtOOiQwPPGeCM3pibgjemgrQtIkke1xHy6LZjmlVlaJWJkJizBQAiQEQqlpDN
VWaqVpyqWYqfXoFHpOMlFW2RFiJK+kheivX/QOnxxLMVBKADNQl2lgx+viAK8Thb5LGh7ygYnPCf
8jR62DN7/61U+Bmk+U5W09WSSn8Osd46eifefMHN+oFqJTrgdjgvIrThQMmmYc86DO6dDbgGKXhA
QnuFrvoK+icaFBdtEMOtfgEF43pXXJgld00SV8+PAe78Cu6vOHaS4cj4WQD2JByXt7RBJOyWp9kS
BjUVk2b3f4KQAZVdGcK/2rWB+KMrr0K9XWp58ceHDZvtiNO9IDS4zS7aP3n2/W8wNEjdkBsGp/9q
arIW6ZJNhqPNmdk88lMjboRL25Upx/sEi43pRNMUvklVpyqfGFB6bIyR55rIwnbQz8OJxnX/S+kU
+bGlcRGlPIDR1AGUArHytQpd+oyigQLzDvbrTr13nBfClFL3eX7AWNSfe55IKH5oN58fsKhdia8y
dqkwJ9g0mY0mJuvml0jRTdX1zbwmW/pDsJW3IuteEZEqrVWQO5BmUSMBETsc0Oz3xYphdboJ+a9Y
Fa+KZL42D1iovA8i8JELsPOkvaV+OpUkxRYEUIAVIfKQdd1QYgYDKCn0kuWkfrFBz2buv8ytReMW
LFWVUJr3GozebwGVNXJ7mWeN2lggYPKlmsssWEAR7WzBEqDu0V9zaIc4Q0tLt66VYuGbEODRWYMq
RslSOcrobFB5583kf6C2Xzq4sBJi/ICvNQUYSdNgjl0+jx+ggWt0WE+3XafsOUZh7YTGaeOvfzcd
zvukN6I4uKJHlWTIpdwHqbyfCBDqRQoARKtPj/6yOJhc4+re+04qIbULHBZ203+QEQ8hKCZASiJp
hXoHW1IrDH+QwD/XjBddOgct6TNxPOl8/1BXSl+P+5qAUYCwEjCKgJRDDR4ixslzS3TwyfUlWH4V
gxgBKsSdrKBC1hiHcYwssOojcZ8WeKWmDjanNDLijjCJ9Rv3Jl4HBRAIPd65SCch+qDRn8L1Xt1K
ZbqPw1+zaGXiALisIL0+UfSJf02ZyRiP6ifqe30X+wwsrM0xcqxdogrNLNypoHpGVfSHESBr/UtZ
/rhAP+ZfeoycASsSkG05dssq2KHEbUFOZJ1oUQmQQYuV440HEtwTHuyrUmFh5HZR6NhUD9haKnlE
O+SERHjkkBOoTRZg+NJoBnSIr/iOvN75vFub6aZtGBOrZzv3NFdRo9Oh4A4ynkY0oJ5QGEOD4VuO
/3fayhFO+Cm1s98sVJDTNTaWV2ViMQdQllXcNiOxt2Tn1eLmtZQwbX1BHeHoJfnpaCQU61MlrrXh
ZIqVN30Oh9aeG91RgD056+KW6lWG3CTO2F1Kx90MIQv+5fn5ajp31jYenHYeOaAIca+R+BFQM14D
BNRkcnAA+gkBJz+3UfhUxXk9vhUeRD7rueBqYlBKNyL39UaZN/zKJhTaNz/4NXQ84IQKhVhKjwGK
BWjvrOo71XBg3BiHsWh/o7JiNYRjEn4+D0cbfdkI4ECG4nvIJ4TED5c3chYMyIc6q+r/et0sgwNY
xAKKYYnY3PdBiDop8fzSDDNCtMhgTE1S9z+0OPsve0N4GsueXgfWUaeZk1hbHGwwW22p55JxcBl7
7EmlxifR292b36zfPKVHKQTFo/MB8EoJ4P5h23FnWpsSYMaKqwJrWqaDxF2BEvukYLJpCpHJ8Hye
37vzypM1488u9ghSqVLZwIHxh6/eOTg3NJMYyDeYiLSw9QCr5MCVgL1ejsktbSqUe0p9L3hWNHmy
P32+iOuh0gdvYQR1vpgJUQ0ZQO4KMR03895tzmqoyOb0YPl4u+G6pY4nNSKGA9+C3QZZaUpM02Pj
Z8Mc7dAmysqPWJiQtn8uoGd/bxqrPFRCfrB9D8CGMkIIPsfe2M7WwzWz2crfYVCW9JAhG3bBVzvu
sZwjeqad8MToSo1eBC6+KT2+LEM52in2vLCay987FxjZINpZNX/jNbumCMz8VXlcMkSr3auvINeG
8ny6tj8Yx12Bs2FeSZj47bUa0NYfjJrHCHGdyM5tN7C2uTc2uo7ZurIgrIdEvDronfYI357ttdj9
odRFaV4nILUtrxcmjmlp4GY1+g8g6VMIYj82GUMb/OhWQolqufPEbigcw+z1bRnH3q3wmJHWL2jc
mJgpIlKBswfAUiCZE9E9hS/g6Lsm7DwcD0MJX41Ft8A3ymBoz14nlMC7WdC7zACdwqG3nayiRIVD
GWsI8mpZQXs+qRDtOTJABhED5Em1L2GeJMCR3QRqfsxigeYM19pDAF/xmVIqy04FHdnhEU7y9C0F
YttDMwBi3b4NYJu5Ic+eEhFX0UbLF6132RYXytmTN2F21rZM3oGYPHsbtRQkte/ijtYeQAwhAyxT
AGyWKTqjn6FF4ej5jhM8eevGpwOP3xrKgzTrv7tmHAz0ggpyNuHcv2VBuMb1kPdjxCfMbHqN6vkT
9c/XOsE+lyzfUc6eUrAvPWjzRyzcaz+kcIpsHcOugkotF+W6Q3QMbnTnptkE6Ft+UW58QAvroBa7
yJ2JWVI/t+klj9sOP7a4ElmKQFmCsuwF3sWdPYpJneXRpK/bDpTIw5/bUY9yaAlhlCmQdCe4p8DZ
BXZIlqlH5KjOf5kHUzxOFN/feYAshoMao1Sptu7iPV7CoL/4WkMr8s7JvH8VmbJp+/0OPBd+3TpF
2NgP4V1sNR3PNHUVSFAWVgJdHYMc0wXWT9kNV61vFFMEuYxzGjssWCUPLVFXASYLhGMNy1mZklg5
wG2wmdlY9iLH59mft5GsDzQQM7vSQMt+42ihLyCWVpf3DTx8xE9/n9HL4AInd+1idXiLxje4DF0+
zwode5/7/oIY9UQDD/tpV0SdXhSdYUFlQ4W0qc6z3q/7afzyZqMErqv/QKSfgGY/i95eQm52xfLH
H//np9qmySJOXb4flTjCqEs0xBZfo1NFOOOXlDwZb+qDoubzNCY0C13NfQeZQHPmJzUoUfX8oQie
ENaClz7iHxMbGXvW6AQ3XXfQejz1q13wUXlf4srzFSDIoJyLQ7od0AkjS6IBpNcShDUx3Xspo+l2
afoYgmSyJcnrWLgs00RKPWMGDly6gDV7ZSncfL6Knf/ebwHDR9BZQS+o8qMTxzP98cuxQJ7RoxOq
8Ir+qgHxzn7a3uPW4KfDdUxADe1aaYPh6dFfF+vG6k97G4/KGhL1YmCMNo+kD9hbpjq30ltOdft6
KVB9kABSvxfBjDq7FpLh+jTEDVAUDFBF4H2j7inQiUrYYNDk1p8SGLjPDUUYhGU+QFplcCm7HRmz
xRfq7Nzm+gr0oInzf5XYuW5+4J9ON/P6FH6uysIktSjV7E2KYDCDQgcEv3Xtqkb+Jt5FMRqqyxJL
h/Qc7Opg8OVfUjJgK9J3jPBFidMA4f1HRbQwD9eP2670C24ENW7F6delzRq7GE6G2BX8gMD3Ztan
pE9Mp7IgOcoi9Weii/oRRKLtbN61Ta6Jxsjo7HQPKcAi/yHogfEI0hXmxBIRt5xIxjcM5UJ/JO0Q
M1JozspNxCmZJRKh9OUrnztO1gLqBqlcp1Zsb6aG9ge1Q8ScG4y5I1fNk6XXCNOWDnuovhLFogYC
v6b3qtasaTtr+nKg9CrfEIZNpAApTx25cqlpkknE3mQYCpB2iaT+BTHdB1Myy0BDyBmHoCAx1tKX
z4VmxvMxmKNwhvIwRNGxFzh6qLLKcD0+NmZDN+3yqNQwSnfXuAylQLmcAIdoTzgJRS3r+ke1RJqd
TJt5baSIfgGR3JI7BE+V1cdEre+7jlq216FXFBN3o+KOifxb/C8hYAXX3VgwUvGe9AOutTL95MdS
nFwXZkSNepLc+SeV1BYKwX9T4IorX3d4hOMWp6bhMyXpf6RE9uFCyTlXPIzPJXXjyrYvCHN/I4e2
EPGlrfdTCIBFKRBv3yMf8Qg4nR8zWO71Z4hJ/AVWRwP35q+Tn4fbeuaxRDlrVg3NmdIe+qZI/zBn
z4+MmO3NvYc0r6W/ITlI5lfKQ55BD0rl67Rh/y0CLyzv+SpSEsjA5ablrrlycOtNWdYPRdiRradX
MyluCnuhT8xKRYoiXaRKvxCdT4vQPr4D68sHid0RWVa/zSF0PYXsek4NhuX3xIL8IuqQ4rl5zVV0
STfA4hgPRElhBXxFZxTAaKRaexLUX+rLLaDt5gNqgbc2DD2kIbRLnTWsLrle/Nt9+TgrpW3pEyUM
6GSfPHf1Rv33x7vhcONePZB8NWhAnFUirupCUYhVH33UZ7T30jvOdVogZuisDeLC5VGz9YW2RW+u
lyQsz6h+Q8HxPffYStKTG3faSvuyPXpKbp+0lvBmU23xrY0jqSYuK8g9j39Z16QSMapMhWHmqJG/
aOfFRzZzzIJhT+dSFSOA2ZBBb6RYf81d2MwLNH4sC54IqdtS8YV9B87mng2jf+vy2da0EzHxtGAf
Yn1gAzduZBcycyrafkuUV6ReQDyHKX4LuOpha17E0IYBbUjQVP/fR1iupanhf6onke1Fg+vOzTPw
ZtZll+CnLp/hZGj5tYkKCXJowERzhxVwjh1hRmylL8Oj2ubd9r8IVzWctj58JKsZ76U8DmZx6WLA
N+4/FLTcYHB68utfUU1PeheW9mN7r9AMfWB63SZa7e/jz/ZDSn0lyeZohtwYJ8BzQ6vuC0djhrts
tBSfGd90Ttw66WOJKzzKU5jQZ6qnEW9V+zOjKwU3pn8fMmu1iK1R+/89Jdlb0yuL1mS5Z+mZ5HRX
rKcsDIoOUiSxRmwnkIs7Mu72GeyTU9+tCVzRcli1lY//fXt5zlHUdi59X37VdZ7BWpL0ztjOl/z7
KOndKHYMJ0VXwsStoRXDSnvEiIbNavNkG3sdF3CDF79APWzCu6tSYKaA0NVTTqBCig6WLU9KRNr9
q2wDtiM5GihX7APzAmY7TEsyf26EsaMwFEbb73UqDktjrW1/MeFdWG1GkglhsH8iACxPtLtAcHtG
jri71LiVeS7MqCiMIwgHrQBIV2L83fMamwH3cqR7rBtNcDLryi+mu1una35pz2Ix33GgperH5moa
GkeUHDaVpYGr3pzbOOnWHa1FE/BHKjP8A66b0s0//hzzJN1qHibZeCAZPMQQVdfX/QJQWrbIQolS
9Oy2RlxXDRUAtAzvf66mYlEJLr3+jiwqtdTX+BO7bxxJt23PAdU6+cJ4iJA2eUBvA/2EX+F+CP/Z
yRgjUMbJ74LhZHaI0KhZQOZxkQwG9G2wmLyLR19MF7+wwkfF4koD5Y9wXNKB83KBoKG2mhbYeR4O
040dgeq5uBylioNMdUYz969d0fxaDj8St0VzM3L647OZCwftX1imYMlU7OAzJiuEdg/fWn4tYTtq
GTHOSaa2KcjUn83OPsaWlFUjCHv+EFb2YMAZ9YFDSK5DvLbEccnMjEz59hr8cewmuwZV8ENexT9u
O98ing4R6ZcymZjVEJ0AjoxMokHE9v7XhFQJcz9gX1pUylXFBbsxElDkGavia1V17016CWr5ORV1
RewpVVJOkICfl2y2QWTdbObXlNiDHRStSB3lE17NKxI5L/VPj21O+7KTu8CqHJT6I0pJKmsvoIJC
IFqKAncq82CdglH6d5mzx6/a7bK62CCjr/xv7/8XFcUdKs8gkCJcTtod0lNEZcVw9zksrzSZU37F
9IOXgBReqmb/1eXwUeBlhqczblDYzmaMb+6piaYcK6B26OuKs//eRh09OyOynBJvg3t6Y7fnt5TO
ZpLpWadkjhlNQARr89c7VFtN4nFpHDF9Ge7Z96kFi9CBtilLMlrw11ht/QYl1kX75VhgthX0E+j4
bWvMDXuoSlxoKQYLTbuflmxYh97h819oxqX5oq1KxJ/rxp2Hlm6fGP/iPxGeBbgD+kWLFwZQt3a0
x+Cj9gTem3Gj6+yFWRvEvpjbcFqEGqzAMFDg0qPzPZ9n+GvkaSoeCEH28OdPVkfB4uShXw9NXV8j
3M6Bx9ktwZEm99YnsQBQquyzz19cF4SPy3sBtzdvIQpEnK/lqogWylLwG9ds/xPOH7BEVCkGiMoa
NHMKLat5toDzOFctk3+hVp81IAkTdVfqmpPeepeGxuO1yXpZLplfbfyJPIcNqXdL6byc8qFa4J1K
4TsgBFcjHsYhr8W8dOCeq5+3emljGmJniyzmeWiwMaH8ZSYm/rp1CXEpnfZ9aXo06lQDbhWdtgVX
bjw5EcgWpjKJDvLlYQjVxVmdCe2gef0hTi+Ziazh8sEpDUFVi4lWJLvRGlEdgwXAirjorSSLctBP
mMGzKVEWVFlkU33zMWVDunJrlBZPVeoJzMSiXFjLNL9USdepXv+BTVC6CJHidBLxN1HcWBa/BlIg
MP2un/HA4FnPP2nRFbiT5CodfFLdBbdHtwy23irGkxuYkAGvNwBiwYT0V44THFnvD41q+grtedEu
mB7zCiGis1QJNAtmUIfjuuyJitic2vBfsb8SIGTtUyLyQl9gnjtz9FFxtOZkCbJgJfVM3Wpe6p3h
Ggs6aMi1/bqHnE3tSi44ip0BmOwg3Vkjp0sDG+UevT6nP3Zalrv646U8EdolRJpG7rZ3prETwnWx
OqRDgFF4nAU1ZP1MiZ/TDSPLDstjFrnKNiRUjs3S/GsNUx2xH5iEtqp/P4MKjqU/0k9ko7HCqLV2
2sDVQ5+DCmzJ0auJi4ifu4nTTGRdeRdyaWgr5Dm6Bj1SrNEH2ZPbhESGtNPqwq+fq2eQV7GtczrG
DoKteIIJak4R/vbGVlSWnjvg7tEOXVtz5QQfYCkJdyTdf4tH/oTU5R0wQ2IWZvuEbFki1QsPPCR2
d39xks2yFPXAL+A/aCobzSDSm4pbnxb//Ja2d3OaLg3NGEvKuPuEbipsNOk/FObQ8ZdPnt6EmD0h
6z0NtuGUDrPqQSC5L3gaXAz7t5tVetWUOgOG6T0BXGWJ/GTjhi09+xeo95lEtpkJG2gjdGiPeQTI
T7GzSQPbtjtyhf97mXMonOVCRR7T3TxGa1DBrvee+CTcrcmO3DndmJjqLEI6TTqlcpZZ0/mMoSL9
KtFYbMbZ+ODYvcaMs3BBPhkzed564Abb0euMRcCtovBT0dNC/inm4DeGWK7gnzAos7bxH3lXUV4/
h54BUuWX+dsFJxVuujI4z9UxYE4R+tk0FWNKIRzAvFynGJhiDb0kCDiyHFmGbjgGy5vWxXP5veTi
YJveN4fj+E9vMlAcNtszsl8czhTlmcpAcpuptaAxluc8nIVuACsetunh1Qvrff7iaoP3pVdOb0KE
EMTthDvv902UDlt6HRdiUs01VB9F5A1qm54mNMtbMeRZJtJGiizEV8A12LJNsqJhBlyowY/jXZxn
uCLrupS7aZA2Vji52cjeZBY5CYyA594Wd42AgwhF0pr14ip09MXd6oIc8fxyndha+teQ34sbUb+h
TjvRmR3n1jptnFtNqxCord8xzXyWV/wxVLm8eVfqxWWvqUkTGfGwy7ubYrcWUA47XB+Iphm8N3SH
vbB53UDkSbfMfC170ZFYS/iPp5iQrRaZmZCSfbw/epbKneU/18Lj6XvW38o5Yh+X3aLpfjsy/R7c
PzNxlubBdSV4KjYogstvMDKNiuIw3MYy6N3a/UqW6X3ruu0I+cyLNATCh+FqtndBHWvFGX7bgy2T
leMIJGK/cHpKRg+SF7chGbH9a5FciB2t16cKapKZBFyVQuiMaNJHnKgtVtiZIbA+yUWKEHzTqBzf
N7sxMRew/0Mc5Eq0pe+xokkSC97HebT49WnWricwm5TF+K/BrMFGGjFhOosSqkDGFXTA1iis4Ocd
X4cTbPXpFeDgtbvzEISn9FfApwKNu7xeoe5lRl8RDiuRFwPkF/gpAkXaj/AVuJcRZw9AMePUGlt0
kvZeQMqrCif72gxKmmD4agkIiZ2T7BRGN2Hk3+Sws/C0HafpnP468GXkYhWM3mVAOq98IoyLFWyq
htKOdzE00sVDSVqmIT7qdN3pyLlu1pI9YmetcW5zKO932p2h2IixFWvDfAxbq4VOCrvuVlfzirIx
CIN9wu304pcujH0xXRLgpRSHdDnCUYPsT88Y8fwEYcKf6FGuFB1ckZUwog2VTckkmP6UYs0u2ZTf
VjudOkaM6r90YtRFlthZGdBLRfsCAdspF2QHfUuoDHN7CZCdyUySabKakpkor6Sm8S6db7EUgB4o
TjOWHO30oRGTg1CNZEpjjCqhobnAiIeagnaVr2ImlVn95q3Zq9YCgPuu474G6TTg7glzip/S651d
mEMtZ/kQ4qDTOvlBj8vOcQr/cH+N/P45LBINaK0wHVNL/pc7PPsYRs9XVRk5t3Ecdz1fR1SXWXRQ
LR80yGTETx2UmQpNLHo+tqSYdnzj2cBOr5AOO6nZzz0mc955bNjWZGMwkp1nXy3jNl2kO5ogxTuW
hicei45zn7VTMFi1mgORk8+R9O9xJhNtJc1mxfjGgG9k4y7LDyeL2VAEHCOZMdnWCoNRRJynF4B7
xqil17xibWuPPcQ+e6yNgbtgrlEURIWyD64RW2/ZK0KjoCYoZT5GDk3bgMDgKT3kryfETWZnDYwx
TUP3Z4dRdKNm9q5H048Nke0hA2H7zZvxCuD6mAUj8rcno2CjFL9wHqNxhd7SuZNga99QKwIQPXiR
KVxnKZ2rSTgixTbh+SQXaIgBfq3m+RnQXdnYeawPgQwe4ZP2mLuxGF/mZHJIUlKiTCqJ4lhEAn0g
0tkbmj3LstsmEJ1it+1XDrgHrVgowQSGVZwvHMGqd4LCV1M23YhC+vd+HX5j8yjgjK7tm8Ck9ES+
bmZEll5OrhAldV2DVcHef+VXaEg+3cfXgux0sY2kU9eeE8nvXWYGq6oDb/MRRM6G84T0ElFfG/Gq
zbMq7tNVkxcsdd/xyn2EnfMvKmXJaSj8y6HjW/SnpJ6UfChjqVWnNJBAOZ85PVK1Ruzx8P1kyzo9
UbTi2Wn2K6N+8SNaa4QB3xUE6vWqFEmkY8N1UCn2pfTPsDKIJJ9uPxDmT428/xZuF71kw0GSNE7W
H2Qq2mn0gl/WoP0wKJ/8E8ICg3v8rFJMto/5qMvSsuSrH5cBrGPCkZBLB9Ykreq+nMKu5krBOuiJ
D4u5bYf+KCCUZ044zzWYuf0rQwNTcevotUoJuEnybChyYaV6YVaIXLQZy/PDZWZn34WTzG5OiFV4
x1nooAfen1E22ydRbWiDfQWxKRQE6pKg0RO7k1LVtQPDfzlmPf9ePyjwzFdmzP1enK4E3OmptUci
GpjlMdxpOEuC7mUMq958yfRYVXUDYFjSG75wSO0/y+XAsxFCVV21H7X8w7u6B3Do+0lOIdhA8tkc
cyEG1nBef5uWzTEmdEdJUk3sNYMY2LZAcnw7c0hU2l+9DjPRHmXLyCU8WkXNkdJBlzL0L05ooNBf
PtBmRAWG87M0gwr52Gn9b7/YByEvGAbHH756GQynNI7Exd7X6aiPiJ2LW5F9EGRAOkJ5bpH/mdyz
ZDDnuhxOCI6DWRlERWwzC24HLikHzzTnRdooGUZutLkXuSjY4iH4+exxFC4xicPzZuhIXyXTloku
WoaWF/Kc04rrNWz1AP5mqdgM4clcD15JqB6nWsNdmzt6O9j3tTU+I/4LyIYWkgiw6GVcc/ke+sdp
s+7vtYYKoOnDrp+hXEsEJNCTbAMJpuOh2tPx6/e9jP32N0PGRDWfYIlAulQV1eFiUPMopWhHxTQY
yb8LP1CejPvaO5TyTUSRyfJ0jMn+YtOGjGUa/Fqtr5SUScJfleMDLd+RoQUVLLd5R36qNixIDGD3
Rt6u0PKJk1JcirZ9ikd7j1Zvo84WNJUKbjrJ4jE4T4DvcYU+YA2HMlCTqbxLJHmFGCwHWjikaVTc
PmTwXAL4jb13Hau4s1u+oj3IJ2DJkYbiWPEznBp+LNWcn+kSPSnYBoRw1GeN6zfNz6IJLuBNQ5d7
oSdSHQ2z+Gp30LHisOvVNatMPq/11bRdDGwIXZq/QqixmqBdSdnDoL1EYWs5GEvDrdODBWw0W5/R
I8bFUNXa4M3uq+nd6invXqvZUgzwxVf0x0jjMliFXaXfi+a1C1Db2Onq61tND8x5RtqhofK9LtuO
qeLVbtp8HsL6KmaWIHUZVwNDsoUPpzSjMJ/fQ1yzg0+RvFHGvdFHioOeQNpC0j4yXOLHvAHbyVYs
Wmz/fI9yQBeAqjVAiIstmWX0g97S/VciQ+1rSEYcl0Ptk1e0XHSTxdnsMZkVBfkkZZcEa7fDKbxZ
tqta6sHg9q3JgnjuvAk1zJbcAM0bQsIj+nGZJmWTSLP49xtIfgyeAMXksHZAsiFGvM+hBdCt8ffV
bTQbKNrh31fl2Mpafv3rNJUlXwhYQekpoO3bVDDn8joZcu8VY8eewppZKIc5blvQ0XiT9B4hEjNr
jMZ8PiDpGAsMufBynjxzX5We8r4Tsfi3fg5I5r4QqNyiE6FeY38qzGXs1FFwOlCVl4KpLfjg0V65
cb1R5dz3DBDYCjcGxgXrC7QW4rjZLitACARJjPZTYjq0e9NXZLYs5gYV2Rs62IRuF6yLczLy7BJC
xE44rPlxyIO4+3/I4RrqZPhYCsjkpR/gJabChcpKVmIRuFqmAxwOgnVlH9jp0DSOJVjmbNYjXrnk
vHu5Lp7YkN8O8/Id4opqCFPu8FRp3vgKemYP3DBPy35Q7jUuqjBEM4ba3kLEZGlQtUkjYlFckQ5U
t4pWhujyxBtRWIJ1JtScW7EcgrnP6JNe1X1/3utKceyTWtnTpPvs4XQgRpUX0e2xCj9MyR40M6wN
6QmN3/511n4I0Yz36BU2vVgYr8JOevnNdDamDuWpJ4TGn9agA9GDO+KP4dVSgjJ9nwjYZNYLH+jv
1S9IPZ96to7/BvZz5lJVkjFaYt7uDEduzQLSxswPxwgUXB96b/GXcWNKc/Ym0SF1EZrPnYzZmyyn
Ser+NIRc/Di7pL8gNIPjXImwhCayI2OveNNHmfslKVlUBbrdvkQMO4ILwkSh09vCvx3Hi0mYm6Ry
1zextlRCBjrilxBo9mTnpNcdMuMglk8W/evvu+nvDStTommTSXRJpGBHCj/fznCR5XEx0/CLG3ZJ
ZV0lO5c7u/UEgSoC3qXhDHS+ppIi8pM9Ay4XytrlbdnROGvbrW077ssdF4X22NUXBcva8StLsc8M
k+0j2yOVHQwZ3tPkVObHjIW8m6GKtTMCxkR+l1fESY2zRDhvco4skbL6/ytQ9yZ12TvMlrig/P+d
Pu10iGZ1wImH1GkimMj32MksGbbuzTzZQaA/MuHwzpMNgmPsCbRPhUcUbO5i7RGP6TGncVeGMsF0
1ykcMznGxMx1iRkaYhJtKOQB2iI7jClXROgdQYSDJOFpn51krWp02nBdngoGWR2yvbglvSWkVzQh
ASHmunm5nmi18sTxDZm0QVyvuRlLW8IVZahVhofcBkGONuRdUzupnGem6bXYIb7F5uDE5ayoBcIh
++qSd/k1P8IoKy4TjlVezZCEPD2GFEYoF3vsZIDm1wKI1TwESg7E5h28gk6R02z3sIqifA3OPSzy
z65MPo3yjcPusUeVIxwYvxVVSJtv91mip8WgOPN4IPK6MHCkH756WmjMZBIv16srosC/NHO0lFbp
094mf4iSOMXFCmPtEV5qtkA7/XKjHaVm/FN3IE/McVQhu21W7cLvVHh+vOnuwiY7re2E2gaoddDm
WAQmyweKDQ4jIN9rLt3xPNg/BW0PRocIZxapMt438AarhoVZx3Xu+e509Jln+yvyxRLXTYCLXWIB
blp/p6DKjdgQJ39oihMB/Vgvh3zmex50+CAcMVpSClK704AKquVb2ZXV3fAdGedIRcOfcIFBtopl
iq+HpFHFSWS4BCnsxR2DiGBhR/bBYesvNQDxci/ewfkmE7QyzidR2FsplIaESwcJvaEKRniaAufX
W6Dpntk5+WR1o1Bw3YasmfEQ7EGfwZqUzWSjH1i8EHVgbdPhXvF1gkSN/1j9ru6nEAhxIVY1ATWV
O4EuGxdKO62W+WvjVedQxsNtGJolN9P/7R4FgTAzmPHle7Wq4U4SkWwZLYiGiBVcytWC3EmN9xqd
aoBLFxhzyuRNUF/+qEFERuAjPzd5MMqyqKb/23nOGWRSvMeatqhy1roNlwBv7GHqpU+8HJk8/jr4
dQm3iFQgvMh6JfHP7VqgrYJCCIgK3+TQb48pPWazpIaMMS92CilFvc5t2PNgeJ8bD6J9MdX/RPsP
zGp9E8icjxue5ouo2g6lH+Vku0qDH1M1SndFERbn70+gxx9sSzTr9t62qc1KlK+W7HBPHrky7Ias
BZL/bxOK5tWhkhd/PhHADmkRN/jWvtYfgEbt9tyl2tuVeWZ8uc1WQ8VINOnEHHc3WDeKRvW7sFx/
jsI/4pjiiC2PiDO+cr4OKz5fXmkSqfRJoh/szxZmCJYMBoKZuJvD3CTpaZhJ8VBclIlBuq4pgfpI
bHwl1OyITbwYL0Xa/2ne6cl7Lg7gygcunsToswgqUxQ7J8Vaz/PVSCFd0jd70Q5INsmUD6UEcmoR
h9ZjNvZPnZSIjuB09aEEaXInD3KeWweZxeNQO+iuLng0hiEfOxXT0pntFg4ioie6saL5c1jAMmkF
+wbaUhlokooPvR+sgHUfRN9NudG2Q3ObrzDPVaVcXG7/DONz2kqkUs0kMlZr5/d8xX2kfrUq3+M6
3vuC8P5eBaLemjjELxD5N5xKfRCc0vb15dJK2GyV0La6Leoy+sNJ4wmv7HLeDDTW6fpwsxEIGvSs
ZMpr3TsXJJ1OgY3IBsSrrsJSlZaQKnz4pZdKZXOnsyqnpYIXRaIoEZ1/SC+vzR/MipegEpTqPl6f
6/eNzZSG93qk9p2Pkr+n0Sml8LGyBb96iBKCNGiNll9kxKD/Ke7V+Pv8MQbbzP0MQrt+7CXdUQaa
R89jGbD0NkmkX+u33thDMzELZO2noSslgfDjX5Eoe48TA9q8JY4bfdzmrxxwhLHcsPrn2gCYH3V9
lqMHvACzHAEIrFVoZbeRwEI+56pgsCSJXKhgw9mTM4QnI7q+ViMO3W7kAbTPOmbjdeBLI1iMAO/t
hg53xf3RVDYjau2g9GYD+doYuY4j74yFXgRIzL+s+ruxfyM5zSRHRcbIJRmyQbGG8m1DsKA+fZRl
16mrFFp4qOXrRl0ARZQPARJLl7K1Tkoel0oE9S3DTd020gy+VnOevJ5rhakSlXcM4VOfePl/LM13
kMvtxKNifpRy14b4tqCDCEzjxbjXIkinrg+ltdE5YhLRPDvakWniSxjeglasnKIqhzKvPvwxsIPc
pmbDJZEGLt/G/6oPdXvBs5ElUAMCBeSwXvKIUeFMdLAE3hCF5RWXVDQAg9697V6FcJvO9UDkVz+1
rnU2VCtZn1k5h6agUVmzV3QzXJNuh3+EcPUB5JkLsfhHw9XhcZDrVtOZ2Rb3EMKUDmvonWDyp8ul
wuWSuAsC8Li3CqAXJVDHXlQLBf6EVVHBgrO1K6Z7CyFANShBkBNb72+kh5inlxdKWJE5B132P4FX
8Se4Gfp+Or50mKxBJWr3zZh2Db/50kwsHcaZ+Q/qn7RHJQc1McYatofDMWEe4YE+XcFtVNL8i6vs
kmMxuGlalrHCxGmIJ4XsLGBz3SqFbenUNCjvcKJ/ymTS5Sf2M66hY1kQ8Qs/zRYqYg+lsfJl8Pv2
yIYRBEIEyUyue1l7DPTgLX2xQHCTg4Tiuh8hDIaTKNaLq7KA/Ph9GfUwNWFK0UmJhuqS7cIDr0Vu
Ly7P9QGL/ZJA1NY/1JWclByYC66Hl94w6j1dIJa4km1JW8rhSnuyx1Z7iQvT4/N9EfhaBY+eSHez
q1d3EWepKiZzD3PotfcuU2SS0MPE7KA+HebUxi3eBZRfTpt+bQlH5PgoxolKku1GcKp/oh7XPIPB
IwyhND1J9eZSq20PX7DgvmNmk82o/riV4ohXJY4TjR24hzP3NsqXGy9B1puLORnmRAAbU47r/Cea
XtLfjXI9WM1ZsoZh1qaBXJ0Z9ezFbrEPi5GDzz5nmjv1O2icuzVeLQbhveWK5X1qvzuVjYjJ2rHe
Ni19E0pPD77EyGoJFrcDFzGRHXLOrilD1MKYbzkK3HwpUZ/TIy1Jai1yvjX0U3u4Qle3ZKwtyQzp
a4iBgQJ9Zn2c4s89p+smBAsNjKgvTOJg3MKLQwhm3Gs6z7YOAumXmQX/CVRri46q6u7PpLdrDqWx
KvrTckO+BU1wjE/uxbhjGW3p/tXEo8GpWmzlhf+oYiD2QUh8TvbQ1Sewkg0zQJOUGxMtRf9TuYLg
7hMH2VOoP6GHcQffXrw8HNhyicWyFZlkjmYxA0mxl26C/nTVUiEUUmu1pBhJKEKO2HrKcZmkj35T
tf25n+8SG4FOdoZ0m1nIbX9KSBWl7qngd3U1G8SUBQ9BxNVQXv36nvk6gcl4Ek+5x/8tkol8DX/p
af6Lk0pbQ+ESdcnbMwq2sMxaT5RSgrpxZGB4dYkid/mlNibxfwQx0XORBveIPJYclYbPuSsqOlAG
MdHP7xXOryG4FbnbkPtuBef4dEX1KvCdHREcoyqafFQ/cHqFeamMfbrm27kq9P55WV0SlZ8YH5qA
hUduYtYYH6ScSb0df2cz+X9TObtaBYhP/c8eIJLu+0Cfyi5hytIUBACAefHhgeUToybBoGT4h8Dh
W09h7TSEc52pg5QdTnzziXhXRio7gausCxgnIGtHOKRZ0jGEa6zm0qVCcgzW90GjznXr6pDqruYz
O17Q25eedfJtfaFRhaQLSW5sxQA9viTzsxO/wKspgPSOXb5vOB3dOXGoio00UaI47fergvgMePll
BOdR43SVHK6hnCSpaYwtOqC7A9SLM1xgRV5kvtFJ0Ot3ozHOfzglZDsKwURhhoSL/+9DDIVfyoBs
x8q5mZJAf60ywxE5ga8yx7dUc3PrHW0fSb8ScdNSgg80FZsGNtB/vp+95faJLhppGC+oETytVe3b
wrvJ/W9fKEkcJQEV015KYoT4Ee/dn4duxK4zqvAA/s3YNZS7E9oNCud942WaDaXAyucwKbr2Uwkq
/QkJ9apUMInuPz2Ylqxfe8IfIUCvvpMfK/p4W32mL9jo3nS3K11ZWlWtV3mH/NbnBE/bp7/JdthH
InoSFTRu3tQa1mlKt6DJ30dtgWlDF+e9FRb83RS4Eg44ImqKlN04td1k2j6NxYyX9wHrbXZQNiGr
h659K5LPmJv3NpWBe9+ejdfru00tiFn1WQnZt24V2FxJDwn1dCN1xpmiMbY5smojfnyVQaw3l9/2
62Zdy5YSlaJzgdYWAcE9Hma0QFcknuOT2wtm+yiSCofA0VLK4LsruTkg7FJrsj7I+RqZqyJiOWir
nt0zB4mOToDr+2KnXbX1s7Ttgs1clCcM82fnW2afqv3SYDhVjt+41bT1QQuqH8MMT21HeoI1SJvZ
Wh/KFZyUJVT2dU1R/Z8NWeFE7kbHB4eO1mKBC9yfDpnewWmy3zLNrvqIxjXRKxS+JtEa1diO1JEk
3wtW3nSI9dNqm8uwcVn+joDbNPA3NwSTqwnCZWZ3yjy3W+pdKod9BIqvpNBNixkXolCz2jZAJM+k
HgEtQ/cPxYfCZ17Kxo9l5oOpL+iUdSBFR8ztqD0asWwLnKiSrSaK5f9jy6Y1gyk++SuNV9s+A+/8
Q83FIajv/vVxjfLiRETrEt260Lq8U6tHEDy65hpg/3NynVaI74oLOP9ZqdfYxQuGB8bniJpI35KZ
FRbVHM67PWgF30vyd2tLS/+QFx31QaPRqBM6/oyGEOZvHGtK6f92mPpMa6J4VI9l38TbiPP1MDAV
6ousSStzix+IB3elDI30yVz4mo358dNnfbzABnvKe3bl4RRpMF2bs+iDvYcuet1B9JHDSMqGJdTA
gFILSDC6T4gA2sOfV0mMYlNM6BhnIK66h8diQgalI/q36RsocT+JiKvhDpLzZf8lRQnoU8EB1uwF
oyKVjl/DLaCFvnOLVi0MKjr1UTPdReDjVWVqIb8MvSvWoxe+8vhRNJgoxgo5Q+eapfGiWh11B02f
dlVUoKiGw3oydwQxTwLG7wnOW5VS2l3Bp/ohPAO+kBsCyi0ft1k4Q+kQg343GTtAGgEL7h/nCfxp
wo+leFDAEfmlUZqhIXO+oCnCFigoLE9lTJSs8kLDRJdGK0wRYXLt6PHsGWxG5W9YsaI50+sI5PJL
yHvTDgrGfj+ONcWNjeIx1y6m7H1Glx3ud3IL4TrynyDHjdyuyMjOtawv0o3TvGI7aKl6TK1L41I6
q676uhCwn+66vW2MacfzWltd1NxulDVFwVgU/+IeQU2p8udxv3hUln+CYMrq4xs4l19+gQi8z1aJ
YYRhUT4mv/6hFHvOd9T48Rs2dZcVZPYEV2SeyXhdIZGnj7YfHY/uTRtCoyvd9QhPqTXgXD3tCHiC
5G61lmCy3ybJaF/k0QlpIsI35c+pjY8uDc6Mj4Cx78iYVnKbdbnpgMCYKzWje5lAMeJrgDnqXSL2
7tiqZ6C1QcFX57VN77K8mUda/NEEAg5ghDZ80N3Df7kTpxS7aPCbOfo7vz9fcUyYThNxVtkFpOBX
np8l/IZqwOUa7lMu9eymKrV0+pSy1sgLZT3K6C2gt/FEvb4H2Es5ztXCvFDH7TSAoaOEgYop5TWn
tMorFxjdXlF6g1R3NtuzBMEbT9ww3Kw/CnOqDQB54QoEerODonCpTpA9LzWoKdVoe9D6dzcs4eJD
MDcDzVGOcWhIEPiTo3hjF/CFYNII2oTHIiKXwxaSJ11i8GkYHbRsMSvZbwusHxS6MhB7uRO42neu
3ihc/QxcdL3WcmitDgeiWooZs5shK5dYQFI6kZrR16ojPWIIb2lDCh3YBijPxkwZ3HJV7K98yMce
ChyAVJijnKK2htYEG9Av7H7R+uPtj4+rh7+G0kPrg2YQOISCVI9tZw7tl2lmrxK/nHYSVDiUbEUI
2qntQnlmfJMhSb8GOMny2lSqGUUc0yUy7+tUTtWJg1D4Lj6HCl13ac/m9QgbF7j7XQMlvo3+e2oP
Dmbx0Dyh3qifb+tk5NV3KVaWf+NTXXyv39dl0QGhPz723QA+TGapl44TtMz8A1e0Q2G8jhC3/CJo
sHlSqQliiuzvvzCQZAilTes2Sm2vV0OTIDJH7C3t2/+CbNDptTyhA7SIyYPjKJ3pY3v6T1chSX/n
pbkJ6i61jgVISb5j3rQKkO1qGNjtKnHlo0Etw6uE5QhwIv2gzbjCjLC33RMeke8ahWjaoQetOEaP
ze5E7PqkZkOoSILEyJi0WvdFEHyUcQJsK5K0HWD5kMWRBXfCYApKONMxQX9fz6Dr0IXpfR4N2EzO
3Jx/8x7er59FGofg0Nyx84heix6zADbUVpa5wyEybjytoZdqW/o2UcaseTPLSx+DmIQgzN14RIpl
l8yIl8zKi4PVboDKVgNWyALWdgxWeLD2yWp05XWrG51Ei8IYLjWbcCQ2tLaIu5K8uwLUruei1aSO
+ybGSwQNyj5uPA9x3KS5rTmhQLiOZ3OFyjrBkCJJlylt5hLtj7Mw0HDTWGyHgtBq5LfWLqJKFCTC
kKOGFKa0l8vC4DOCVutzX3lEDVG+fmuPSwliBwtduWOEBxURDxvfTgP998w+xK64Nj+cUPX3rkMd
SgeIhoGCGwZkxfCjCchtTlY2AkewDKYsDvX6i13u7WzVkiTKRXHJ7MLu7N/U4BNdZmPqEmlYAI6P
bvoFMxZbyH0s215jsPWP+SK7obieCGcSN18EtMlNYEl5JAB1z8ZRKiJ+gKtPlGgxgflNb9O86Rq6
3NKdi6iUX42GO3d3m8MbRr1S3SWE9212tdW4KK3tRLwYHn7+Ve1/OYeofgFeCGJiOD2GPXL/cjKm
UFk6wHIH9TiPjbmXpHsTi13cjFDO5thGvaoAHTTTztackvlCrbTBNtp0yXwlWN23r2Gwp7XS20Bv
KZ/yZChG2fHkJApGq6OZd4+jnmdcIkiZF4F7UhduyKXAFydK5zIzoIXV2I/NHu/G/d8uB9cBpS1W
Mnk/x3LtUGLyq73TFz5NXckEwaO/qottLOeF/enEla2z4FSOGnD06xEpfgK6Bn7mjFRJulNXtITQ
474kaeXCSic2zDQCHliKNsQRvjrRKr4euQ4np8wN7WwKbR99mN4O7mrM1Egc1Y0rGYoBGow6fN+T
dwWvv9Ku6vHXXTnXnwMPRYgu+HDRnrC035yDGzJYjDteCxoAZZlCL8t9y3D9toiBRx00LSwdjvKk
h7CAldUV0eokcR7q0BhG4ykteEFTK3guu357cU5fQeQzAls7XhU5B0do7E8LQWKDFVy8YB2tE34L
ff5EDNGqLudFKauQlWPjQK4TW2SXXyaXHqLj3zrkM/lb0z7PTuRRX6ZkJsqqE1Rys7EObP72vpt0
Wpjf7/CrO9BzUBWomCZp1ChAlVxVUWh6pmppRoxSdc4CrhWQXOEd64QKFZRNxRTKq/6a9A2RHGiP
+XTbmj8ZTdkprbEDl5ooigVjNLq961iNaOOZALvg81iLZsJno7LcIvdlYNcQS1AQOa3QbhrHwxe1
l7WRtLMSi/uiCoi5SQvgUFazq5npW/Hz9ZWG2XqcLV2ja732+HR6ZtmIOA8IEJu5FTBIJ9LzXiuo
ciLE31w6h0qZss0RDCphZ6KC49kdrMBSfZOkDbH5i/jpEh3AaEOavOgC20h9BpUr8DhT/WLGMKfv
W2oGCDuPQOfbsCgn5krmJuUeUCkN+9LRs84bPpoIxJCdVJpFGC9JvlHQzTkGBWspuAfOubQnfiWN
7LctbyCQyim5U2jXGlbSuw4jugfrpiAVC92iylDYR8N4MJDFF5k4mVVRh7OfzH+ArSSn4tLtZt15
3YCiE4ZVmrBRHNWU5CKHl8QKHPnn+0ZroXkusWvFDDVe8bxHpaGgdt8Tsih7Wytcjsh8e9wonjgu
FhjtWJiputuPwvcXJqsHhLPfiK+pFCB6B1IDhnQ5ttlF/vDDCZ/hvEu+Lj/dRVkEwmq3Y+GmkLtN
M1FfMf5sdBN+sifE5AnSH06ESYImCuczkUfBdBkokoumBoZ1X+f6XDw3fOa1ALfrYOZECbQZlwYH
M+GQXdk+gkT9VzhU1kxrQaV9y7d7YwnRL1Z+NkmqNnl2R/X7Gjfamt8NA8TMS7kkwYvwBojxDYQ2
SFnngm1LBIFBtCATtAnOjqg7YNkj0Nc4JN6OVvohb9LoYQJ4c2eczfGIIvSOK2Ou7bog0wjgBv+D
aOr6zhUSCCyXspgle3b2KsupfnsKj2o6y2v1iorZOEemVc+ii1S8cli3UVJawDkzIa32N1D7RKNY
cNkL5O1Hdd/oss4vCTEON2Cw1e8Mc2qAM82b0+o7Vd5Nok56ivkAbsoc7JbyKh8DHa+C8IODc3SE
M1Noe94fRR+XEHzDPm011riD6aYQ2LB18WmgxV2zq1zLf7YpzUKErhV27jcTxBxz7aMYiLwvNGiH
aXkyPhmR7BwlXlkm/tGu+6Gl5wCdYsHr63jO1zjkFYjVKzE7DM3SJDnmSOTqfftjKy5A1ttE0kou
dLleQaCaa9rLNmemiotw/BlsU8u6aY+wCcbpFLEYy/ai8qLXYFuaVR121K5JPuKPXwvAhDN2xUxA
6Hq8ieomm/fOv/+g6X69aYsN9oKLJB4uH0h3LN0l+NRK83rjqjPf+6RjZLSNVInkI2UU+tsJFqwT
WmkovTQDnKVpu/66Z/grzmbTa77+1kd4Sb79Wu0R2HatlSQMr91Td1KoCrpR1xMBNch+cIViMM5u
2GzGaE/cFZ5CIUEAQBRsjKOG13O/soOCytlmDuB0MLCIknxtX/VcybavVMRxm9NxFXnySXbyge+d
zrJ3hrvxsSUgHo6Jz+xHZ//rJFH4vEUooHgeEAMcKkhGcgge2fcRjk59MXbQy3A5b5o2OeRpdEl6
zuixmNRn/gL2TxGM60p5M/NiAiT3rah58iBwc6oxpToPbSBJzwSjHJUcgAs71R3faQaiso8u2W5c
bk55WVoN8RE9xS13Chf/QY/W9TU60Qfo8Yq0rLURNub/YwPU/Ka+AuM3+lRMECzcsl4ws+B9ZNKq
ZAJuHWfJ4L3rIyBOSoyxlYaaITYYgiFiX07cR4hiiySdb7sTkKXVsONn66oj63MRu2bNtk/zcwZu
1csTsoC33k3BEKPSi+odpzf/pNhjjeTNEgKvGlKHSKoJj9Z/E/KloS8yUNdERsB9Hme0oaL4eM72
0G92ipFV+yvVdyMWw2Xi0I71yW7/F/KXaMe2Cmdkz6bMi53OuvUa+DhEbhaXdrc4d7R8gh5MmSj0
9lWCe3fccwdICG7lzwdM8qmClk9bHDoSFj/2wIzIXHrzxe1nHd0ln7jQtNGqJCyRTowCh3CQCpMM
xh7W+871Qm7A5FcAsShl/G0olFV/DrGdGbB5Rmyceu3mwjNp2tl3apcDIPmpT2kH15j+UGpRBwqx
iNZrPXIgLx1dQwMtRBJ5b/hczH2HZhi7aimyEtVbZ50gmAqhPu7FWK4TlJZmNh834KIYSsMwtHfl
oLAiq60eVmmJDLTIh8ciEMM9b4C/+O/C7IWrwgVBvFbctVIVRXv1QckaBEENmKtRQYZcxuTOcUt5
t0s6sFmznA2QySJ1ELwiPi4vtoH50kfK56VHxU1FdjPsPccgP7TFYo3od4X1POnV+bhioORGpeCb
7S1LBq0M7MIusXJN9whZMwJIokDW0d8Zx1v7CxgwlD94vOJK3WESdVtaD0ILxwtVTPDD9DConkef
E6x2+VVe0bj0xkfXx/H/mNizgQRvekUbFrbUiz3W4d5kW59lSb8o5CfEBAK+FHC6IAQQAeJzAUO6
j1LSEFeX4GmatIQQi9AsOn4hsQAyL1TcseviT50r+XzZzSnfjcV69RHibLC+3bIG9tE1u8FFSrF8
vVSHtFaUDHOtc7zu4TiGtrd7/k8xZJTZPU90h4lMwviIVcK9ZyPpq7wpqLIp9W+QaWmvuOM7+dzd
PWivi4kT4jsQwrCWojSJx4Fwdnzjquhf+cjcrV+RLGr8CsDIj2PWF9l71xxvjKRnmg619fl/i4hW
u4+hPBvqzYFfN4QK/SdMzzyhHvLPVXR3747AEZHyamV0GBWEXTtJ5WK7WTRXhbF2fY+EYPK06pGp
gx6lo05dDPaLJclRkb3Dk8l/nsvW//KZREVOuQW85fQ+Fg5/Psrtjkk+NSfpdZbUF50UcJVSOg2E
KYcqnPNgmNpWbSenny9QWdlyuy3VHKob31Is8qDGP8+97iACvWU/gxIefiCUZfJSk9AetkbZoGjw
Avs3abKnMgqwXZZbiJUxkcwNnzV+S1vRjzdkJCljL5BKL09i/03hG4AV/W5APQY6WYDpaNoFtLde
KjxvgQbGAcqhn6/sj8PCIUgwpzera4pBff7eWmY4sfwLpLA60+wlLgR8iclQvp3/7AW2qXHAUWEq
izOrFhzXh6oAg5eDFaI5ngJp3/4CgjscA1WTTaev+V+HXl8Do0KHxfOt7yaXuTLwpfnVZiH0cdlY
x321/wr50SRi4d0sujp690h4PcSn/Zh9VJtnHp4cTK4RPEOQvRDHKA9puh5kOvFj8IC358DjPNVO
TuCk4dWgEKDG6yQya4oZp57+N9i2yCXMNvFIHcSrFEeCX7aEuexMalLicy6Oj+2ip7EsqrXqFR1o
ozBM4ZMVuHXM9yUkO5nLu7cEug23cF2Zo92jhkJ5YySo4DDs6wEurAHt/JVKfaWr0cTtneViH8uN
Tf0jcxTe3t2mkl9vpnSrQAMcu7g7+qe91extxLr4Fj7j19WxhQenOvJmg9hcUK0sOJg/3xE5RVpm
+w9hijVrsvQiN/ya6aEEtcZC8wJGzivDbxWEooVpLyU9E/VS0+Yg/WrYwJaHQjSF4coN6w2aSacX
mW9x10/IJXyUPiy7s7MOTnpiZrFVC4mwIkiSv9f3X2oNiR/zr8eF4rXdFPFKC5V1+SdiPeRnXYLe
1RICGPFPcYL52xRY5mxKOg45D8XGrMwbw50mKpd8yqnK1u7KvAZeJveBMIy3JUYqA8/tLQpvra6T
rC7FMfqyjWM3KnB3spqJM9sAUuWEHs+fbipvhWBPZPr7Feov5cpmMTZIc/Oz7MkC7BEDovTlYPsE
cyhTPGq9HCUelckJte+dOvfdvvPtRfPS13E00z11HKjASK9y+dwZcfhYGcBwJ0VZoj0gT8F9yMLD
UFMnp2cXuZYEouC//iYOtmfZdH8x2mw18CwyXu2MqaaZgrX3JWE7l+3irkXPUQur7Stxp88GeiaY
bkY6OXsgaNRpZynPyizC8WoKh3Mb169/MIrM8PJjmDbHKH1+D70seVCYrKibryxWSTKpmxgEXTYJ
D9nnbOY1ohn6FC68DujEkP/GFfM4z3rxK2lK9cLD25XVM/LbHRpA1O3MzvEZWAnMaw8CwvWspHY0
Olfr2dc/RrIUI+tkwZ+x9BhUtrVc8a6QEfLKK6wrBP3xPLLOhm+fwm4tbp93Ro9FGXjkq1yaKHFW
CdFk/x2tqY+4m4xfTxx1hjgfa9CCyWw7v2LXDMJZhMOs6N3eGmmMKoQQga2MIohJSVyvOBgYsZV0
V65+/WhyOxm9xKdjc1q2lv6aVx2qEyycWjVFnV1Bh+jC7BXjxMm34smzVVlgfOO2qJHfeuRgj/Dy
bRF4FbTBLRFoSt6QZtICKjffC513JB3UhfG87ShQ+LE1mnrd4guIfPIQPG8H7FocUcv+fsUeAz6s
yU0nvQURcnJT4BGUFPt6pOHbfuU0/yiP3g5FfOe7r+6E2xj0/2fVKOAoClMMKxigYO7Dbi1YXb4m
gbRH8ULJo4RAVsf9NugGnpQGVgHbK+Xu8VXI2whzI7oeoQ9dx2rQ1+0L6yTCHmmYQEoXb5WZcPUb
hgfU+x46PyKnJFiyrIZI1BF3xN7YC6wKag4dBt68u9D3gBG3/dhT+MeOYrQHwiUuVRSO7c0/vKVd
MzToGijmSkiLq7h+qm2b/Fq6Kg9AsFIYH+vJalX8kqzgkcthEMlg7Xkg2p+wT/YRPPnUdr9kA+yf
qHTeBMBwpwjGKtUz8L6CE5D6dUrijOQNi5VgsCyBTbITcH+xtMyYQONwFwzBYjvRb70nTrXvBwYA
mSNVLdjK6c//OESlAeM/Xc8b8iJ4GsXELS8/fP4L0nFi004WbFNUDRlXIU6zp4Xo/PE1qZe+JLi5
anEf5pMxoLnETWz+8Gg6KSnfNuqyZenButFEXTo72RJ0B//8WD94rNhtaU2mYNEzqG5qJlO1HpxZ
u+u20eD1aHQ1cJfEdySfktKOW4yzliFG3fbb9AECiAZzmrs9PJMISInBiT3FkKtd2lrURgUscijA
aGIe3gsiGPL1qConzJJC2NED1bXj/cdhMETpHUsoKg61ABUEY1cl+MipmZ6iftwYnf7iits+uu6T
aiJPP9gwzv9iCOywQ+czr/xxiAPNANi4ZoZduTDiKAxLL/l3ojwPb8nB6oeHfLxco/Nkbu2P82ST
BKoRkqNlwhKLytOP+sYr9Kc2PC0fDc05jio9MAGQHEVtVGZ6CNlOc+PzDLyEhGDY11R3InopZG+R
ksnRW9Bngn8JoZQU2rETQaGknYJJa0Sq/V1NGeeuvdq4FPqad80CZNRMcjwnIe5zGy4wEq/JGKFB
VBwZ8gOgSgG59RrsEZWoce2ffxM1lfWnWl+Zd4qYhM/JPqGidoFOznZYdriHCT+aj/0kIBP1X+N3
xgtYRjfVmr5ohv0+edWAVSr1TuXj81WUauEu+nKlm7X2TkboQT/j5KibW87pBGWqTGH3a9feE/9o
SbdcNDp1/G359x9jy7L7XKcRGn7rOCDrdCdUv/3DLf1vWhVzHZtMYq2dfEy+3w6lov7tJCM18arS
fbpVBNHFenf8gHu/bvB2ZQiphkx6id+eivM8D7sbva+f/NTrTpLA3zx2Ue+eFAa/V1rhhSFczjvK
v3lgUriTR2NmzF3S+8igwRT2KcNbOtK3yVAOn0bHWceoYYWO6OOVE7QLOb1fBPk/3TqzscuO83x+
l0rgPTP0jEDJT+LOY3ga/3hTs567TgLsKl1J6t6BtEk9w2k6YxYyIocWRlslebNcmIXGCx+eQ9M4
RYa90srgLzFEfjmofI/jbiMxcX958yKVWEDVUQb4On9WEwz+oI34ATOunPtuXM3uu8tb2enMPCi6
d/UxllYIWCgtMtlVmmPmO2Imw0cEvMRQy7UWa8j8nu5WVbOooOEybT4clWxpaBO6z71gbPM2fi0H
KIZI4bxb535+43tV1Lu49KDNSSc5UZ9hCkdYI3q1SgY6yzJul8dk21YbyT+TysfBPvTt/NKFKknR
f++25zcD057FF65JyGuf2O+uOoQWZlbF3tVazZD6R6b5l2kqgBrlw34tDzWgu7QsDXGNqFwHuFyx
wtc+XcHRZXFoTVuROrFnZY18xVrg8OWZf/oj2+C1lbpJvEJiqBBA3fLDx7Fq12UfRIL924L6iKcA
DSqXkhNStAVn3Ma/KqWFUAU6WsBHkvCeokG+1n+4wS9MdXGKw/g8XdRDHuXbxoETWa6VNyq7BUdR
S76DYiz4GSXyyowkwYcaVQvw+aTPSksaU3zKLADnvo2pNPln2k6MybUX2Pl65UsnQBGbRqhxiMXQ
6nC/NutqnqaEITdz4Np2fPJZVU8G47WMPoPeQCDyFbfKleaLPyzlTL96lHimuYKTMQnoWjQObpo8
BQqnOQcGD5ZuS7AQUGnepGfIGc4NZOoxbk35qwdHwAh271q3OvBMoq4gLdN4r/MLnWUXHpwNXmtS
I5b3ahDqRm6Bwdrx4eEfLS6iwtoqXFof8ijPtz/pPzKI3mgjdRrtoujI6YnQTTxKsEmkWGC9mbcX
ZxhNzZNNQ6syJNFnqMzLcO/XOcAbAiQk+MQxvENCNqu4kWop7KJJMeQn4w98/VFrRFVV7ozKE26/
f/gc1Ss/gfJMBom7wdPVojnmbeylPZClAupOmmrcQssxCsqnMDwusZiw34iVyHT0FE5iHNlgRYNL
xEnNF6y416Jx34Brq1s0WaLIEQUclsDIRrIanfVNs9D7vTC7OUvmzrXBcESGlzDW892ZuMVnI29K
dElPtcweuh2SdyA/9AhzbhpFTjkGGKFVifssG4giVN9wSsOF/o8WRp0JP0aOUY1rWOO6EKNj8CFA
S73DmEVvSHSFyBRsGdVYF2jdzK7RnGElnu/MYEBGJqTHdg9wrefbs7YQwT8CHJjZXq/RaXjB10Qx
q1F/MG3XF+Jd2o2waKZnDKpmoY3GiPUbTJ1GO56FVdMTMCVBJR7CLWPuLcNrMFadeF6o7hbe3BZh
wbxCEJq1Xl4AjHdFugS45T58Q0nHyQG9KouISwGygq4Y0oSsTVHf1X5g5VVWY5tWTA4+3OzLRWj1
9fcqzhNnE3psaZNq4/ZBz8j4tLuGIbF8MbAtohjyJvQB06n9ghjVyIkJE/KfB4i0EPaYfWjZKtUg
WV5qJJy4YN/87w1NGB8VkolyHj8X6cqBvQyQbbSUefDoKDuL8GvcQWaIwaD4Z5CQuxH6kVo4D7Z5
a0/T4toA0RC9D25dNRyKJstanUjxRBk4+vorGjnhmFczdsw4iOQPpOu1P7+aFwN3azJRVR1VnUWj
nQdkPJT9sAInHyArHgbEJw27AKl92ZjzjG3ZHfujo9wlM/u9xQcAEsi64eLJZwE320PyUpk0p7Lw
C18Waa8QvxQt2HD6VEGMt1H+tmJH7/lW450pLcSPqNd7kaJdHxYQtMo1oIBR0elzb7QlMsEeDbOJ
upkN81cEyR3S02QiSXkCNCV+xC4DVdnKQZKKXLYSIkVIjw/RX+//+Nv37TzNGWzS0/Y/f1qSNCCt
rj3sE44+D/5neW1+STrGFybP8Y87wZMcHonl1LFwWNkdUJYad0Qcinv31XcHlUVqmpzzo7llgXmj
M4v5r8In/dnAKNng/wt0Mvf0+1XDILgwGaUZz5qtJsgZuEVGSyWZ6gVez2vU4hiLvZ1tRQKZ702p
PQ0ZFm7NZY3NDluwnt0BXsKa92254+RusVOmRai18pH5ogrXbpZPG08Yx38qbtTg+FdKr12eml3s
/zqdeu6G8nhirGVjtNI7vnfip251DlIUOXOKFzYOZwq2aXKJhfm/VOtYK8gR0PpgcWjpyOi5Y1tw
0NxwTX6pvmCjWvdF0Q8O8hKVMWOesU1K79NKyNuFsbIOjPvUyYAiILCezQvgrzNDrhXmyDm0Vmzd
MFCB9WQq4gdscOnHAVW771ugRwCY8RlaYfG+j6zAi+s5Tnlcn2eJ8GOMUIjR6jsSJ56DZELCioIY
FdrPvGcez93+gc2uXc76tkCv+lqpnv//uBZgh95UEvnKKOBPiJRFeOfOsxq0d/S1DD2bVdoBo4Gl
zO3AIWRS4t/kT8erqWbL0Twk252ue9aueyysb3vGMBbVs4eI6aiwJaMnS7yMcS7rRRmpfcVifNDg
3Y13CCZCoREWS0xciN7Nx4sIzX8/hmN0xISOkgXC9YyrAk5fRuAdLIOWs9mJllDgiCPnNFb+dkpn
CM4Q0OLADAmw1GRdaMQVhIifXt7H8Wn3qgby0LPJ4ZZpopyqo7CvKe1TsM1zYEY9Gkb/MVFroRT9
PTaVYFYeFVqwzc54ivyLCT3jqPtNNZ5OZwl6szbuUYyhdMu/1AEQOnD9SyXlQ+R6ZzeSXmXhsacV
ZyEzyIBT3DMG1pHM4KNzrKxs1p9+WJH5YkhCTd0a8Hf+z4/5ObkIjLYc8aiUCYLakijgGgMtZNvP
3OBTcR8mBPGmnMQJmA8y6LGqLe1cttpxHKcMQgJKbluVNCsmuXwlayfp/BRX868z5d+mc+GLrUYc
vpVkTmt55/TKrjt7sY1m0fnjhuwYQ9lqRjMRcNQcSwtPIsxFnIs57uHFsh5+KaP2EH8Yj6hMeH0C
U+GOis95xjA35l5mzlGQVkuNitaTdr/awRQ57JxDtrIjX0ulPGA1d0nS0k76IBqTmsYUwXwkJ7iv
0NN6lWouxdp4LT/DVBNl71YwDOWI+LXX9uS13xU9stbJ9AqCsEi3R3G1e4wg59LrrvpAeRh8ZL5K
C8cFPDukyR71s7Z2GddvRXq3DnU6NedMfOpDANuasuaD2tTuU6Q/fkeJ8bHZRmkwZsOfPVGZFsJs
/QkzWPu3pE1lG6kFkyv0i/ynCxO8zcMywiBbmsCTsXv+P9L6An5QXq0QwAi12p+J0WW0I55QZgwJ
3PEB/Uh9y83XczCz2r7cQETwPHR5ivseg9ZzvkjRIo8wwQqiKC+Kt6PlmPUKEd+UxFNJvX5jz6jL
SSeHk44oFzKlxF8erOHOtc+Wu/3ZAsi+c+nBJqcDz+m91U5x3sMg94qEAZMOcOFjwSqzgVjkCixM
u/1hM6/Wv4zhIySlqn6YjO8li3U7unERhOE9zG9tnx0UYwbRerIBOLCBrmqECdJ8k1r32fuyAzPQ
+6okKgMA6Bqh8AQnYw23zaSEYSFWJRnsj6uEJOWT8n8Nlk5BmSNAhV0GaPGEIruTVqUERZ/HQtYn
b+k0XfcitRs2FjsbZBnedwO++fZXPS6zH/A0NiZXWfDdzKo/XylfxOxViLD1dZrxcaaR+JFMnFlC
UDzeTDk5Rnulxt1eK/wRROG7EkNdrzrRICcoyQwaw0uxg4CB9yyr/vQk64b+fVLHegnScYmfEklC
gUfRFaka3NNkW7qMbGJFv+70sxzjmQ8lUvaL0hK/AzxSbT6r/XH2PE2/FKM8DvW65D8r0dethavk
BJ+ndQfAtKH8QMPP2rdRJx7eLfkOBB30mQF39Pp4xPnMRuoEwGW/DzUogTApY2HcD38mM439oDo2
mbpqvcxo94drDsCRbiM8usVsiLVeMOJ3znd24I6Od339C+IecgSH8SgW0e4aHNTHWFgmVjELwH05
wQdGNRzmDyDeDr9DB/+YrUKSj9t2qdsf7jdSBAuno32zsBDTg6H3g8iUp+3Oe7Y9aqW5C7wMXRzI
tS8Rap8t7dANGIREVvJKsXYOSAzuqvcYO7MN5Qi0mpU9cLMv8dvPqsIQnRFW6b0vKsc6DnR96Y23
Y2QfAoFBDam05ntK1v6CoUVi5A5t0E0LI5REr7Oi+k31gLNH+PxBs1HfWPf8em1EcRRO/rGZgPEz
ASejZ2qnecoXGD1C8bc/KEYJnpnHwv07S1Ov0E4G6IDJvJIO1DfmFYgYGlaVl5GbixKtSb6f+Lts
EHyedtnzdTdUDERu6AoHvMj8wsbtpVLKtGSQK4Y/QTbzymdeq9gCA9bUbvmDSy7Z63rYd+1GvOKi
AE+LHSQZIHCmWHwe/327uqF+Y7xCUk/Z7X2MmkfLqt6GKGdIOTc/5TzyLeFSyqesHGBY5YPTDjXR
yB8TL3GgdeVWrFx4THlGop5ygv7O4D6P/AzlgD8DzNlVn7hIpVYuJCZEVMTOqF/X4Xz6ujhoeneG
BlZIrL1vqKzCOtAd57sA4hR2PVpCStMVtHwJheF09q7EikfSmPJf5Huf7w4CGslbXdG1e9lYDGm6
/9rKF2+p5ZKp9Os26Yqfl2Qw9NPBOSZXqFQcKdhHPGpOz2IrkMNrG0FNex70zYLGCzIIDeFBJEtr
9fQ8CUw3q5InsL8KnzAzxX7b2kZA96r5kaop239NU5UkOO9Dz3fDzFnNjSQaOKdIqHfF6jNsaenm
h71LbTk6VBhpthOrGkHS4uyzoArgSKCuxSmLKAnbwnRTrOzJG0T0OL1K2Em655qV1+UxCkYL6dKf
i95l8m7AUY5b5InGTBD1IwToZfwND3Eb45N5esB5dvgbHLqEuDytckCUfQVT+jsQgKSXQvn5w9M8
N3YLvOisVfwwKq/HtHtTTAXxuh4YtD5u9hMArBEwltWwDT8zhrvRfNGtK1nKscBXarHdZmWKISu+
u31Td/IAPTtQBunq8sad4HTPL/bgrzLXTcIKlSwyOmt+kSSDXYPiyR9PvmSaWCk5YaRgGwrfXJzi
SJ9JpN7iDOc3Sd9e71ed4ZlmsZxY9tchsNa8LJTv1HuL0Ikqjcc6A8VtwcClTGABfbruDg2QI0Rd
ieqSYjGAgssIUE7wsvZ+yyIQyoENdVK+Uj3Qc9Zr/Z+PT7JvI/X8krkQt9KVqDYl9IrYNYGr4rRo
9OGFkzGb+mzJjajY4sr60f301CxKK9CEmk0kdM5SwqExoM1FIECznjP/9ETsjD1fp+3Ni3QhZTh9
jNckh55gIn8Q381jf97moFYWXUxap7SSHaKRBlAxA+bou5uhq6h9iclbdzS93pnlpBkmSVLlxcOQ
8ENvIL5hKiw7RVDjZl2dO9Xu7to0WagpsZhI51wBk/SKetrBa66I+YxwQr9MMiOOLpDksEo6U5+2
7rjPf9oA5Kj3Rf/FBa4keY9Kdbxla/ukm88pgDG7wplWdXJX+LEVHdfeysNX5oy4nE48U2kUODCg
HmPpmHMjX8GxSbFDI2vqhDhwtnZ5Kg0DIymC3Un+doGlH/IymnLegQLKdh4t424h8csb+kGbC69l
cBAhBu1SDtNER8MZSsbzqVlSbXW8S94QC4Gz55SnUedBeG3x74ys0K3yyvfnw+vfkNRkDQg89d9F
jU//F15iLk4nLVC8abUpVnJ4wX0VkVQK14EOsydkOV0k1nnMgqI7DTeUgycU2G17uGorof91ONA6
+laLkA49bcaljETiKiLxMlRl4I0Rb5xkcuJbDALltDVsPOXP9QBhaIjS9VEO9MhUm/uPdz35mU47
PMbf93gqEXefU3ZWLJQNpei5S6hJNQVCFksVhfPkoSlZp9Q50uZrjf1NfNRalRuwh0BxbCuePzOJ
1QHJJhA8mnAHa+2x0Te35QCtObxRWWbdd+jt8NIiisLfGe3dsdskjHFZaDe2cXsP9x150R2Dfdgn
JGbiMoXJgQEXJ9x60br8//+XdIocgykw8LhmtIIeC3G6HiFTE8y7EgY5xQn3QQI+isqqEcOjudDM
ly+gPkyPvii2KWnHbMa7KW2IktYEYvOouxfjbA/sykfN2oXvh+2G6rInymC+a+wlhlX77cHm10h0
BhWUXG+Bv68DHMj2/11c41kBm6LX55OL87kSKESuHWS+S38UWq0DTOWsqCa9bYHD9bjfpQRHdigH
HY/8A5uf3Znz2loyO/s97cQGO1C0NpS1rNbzdmbrHjbP1qY3hc7keOzIFsOVtrHC0Z8CIcsBAuAz
OTW8viXR9auFco7wzubNXU7X0v9QXt8TSOX635ENQsyq/pmjrYHhHH025dxL5fPPpkxYZiuyxB0B
w5QIBc7xsqncggkAiSHrVnC3umcpWTFunwGJzKHE6jMl3fEZYeGp9nBVV8tCTzEU1+RV5b9rpulj
wLRlBOYSOv5MHcRmQXpuIjZ/klNZzM0gx0MrRr9XPH/Q1SVUiMlCfV3SNPbYA/RqHLaaJusnS0hM
+q6m514P29CkpY4gQkIzW3dHZg//N/hoH+lR+TA8tt4tVssPJhcq4f/ql0FP33AJ1BNIkGSa7Ge2
e/fnMglkGSnzuOlRp4839FQ3ACyMBpQml7fSz842Ty+XqFh/DDTOWQbWL+4d0No4v9l0ksEFobPU
nCG8+WiHBz07Gcul4hcBj2bsyEuyUmB28uPDb2Iz004vuyeAggTfm4uzMRzt5NXOervaKev5uGSs
xzajv2NU3hqgZ35fWuL9J+TrcRghVA4NC6olrQa2QnJs//05aKECdqeF+1AgS3CjUoE59gTjg86i
Y4RkCS8NNK7CadyfWXCp4gRf5qeb+vQkfeMvjjucghVGMGm8yjX7U2b7l1/B7rriVBPuEB5ZD3WZ
ZWSHbL3YjTBoCSjXpU9h+034Hwy8ytKM39yLRw2AbCPyQ6MBlO8PB1lunDEzHrOpOgP454KCFsoX
ulHeMNoSpBfuqwjHKWli44vsMfV906pQbLvsLcf8KE8/v5oGjXFmbiIQCs2eDc/wSVwhzVxutZn3
qd+w6uQUZIh8rHH3dNdw/J18MU5/9eUlehQD+69jDLS3jze9Fq1NOI4IL6MnX29r5ToXEztvJWPG
hfS6PE/f0if23uHxWMdpzHVUhFvWu8qz6LI4FTWmLIFlnUfnXkptnPNe2rpKKxT5WMYyKT6bK/tF
LrHVqYWZBPXQBwIY0AaaC96Vfp6RYAPjN1MdGY8sbcM/De76UE+oQtLhC8i7QZxM8pca6PrZlFlN
iUhjwn+3nxHJLZH/OEpbQTJ7WVQNfZLUIhdgM26Qa2RLgEj9Lan4XzaVXoXDl0gYU709vpOUY+Q7
Co9WCqH5OAk2gtbAWV6tjPJ6Liw17486ByjN4ZTT5KQhoXBBmsCWBhPwcrzvxWzRuJQ4Q/KVfq27
3YYlKuFHR5+zdvr62y2swamc5/LODrXBPsBG2RsMSv+L8pW8LQDoyXYBlCiGNY5JyThGDJbUO0/c
H2aDsxL2z2+o1k6tCj8v5YX0jWz670VHhd2yOSLPG0QGpu/Se4RxXjNQr8LhlNdgXQU9osxzSH9G
+M356qvEvj7+F5ENJf1OV9l5/jxLcWkYtsjNtUUC7Bf/PHteaZvCHwJH4M20ZTz+lzMWOuKJivuu
Ut3pROTeirmqHZofQKfnC9yS2gqN/oX6ZxVkXdmf2J0IgoGu7dQlTPGKi35qDTreCWQOoOHbk3lc
n+zC2xqAdngEOEHij3pvCRxj5x07avhjXtVlxZZWg3jKfRQ7W/Bvp5UjRQkdYIjGdbDnyglEjaua
vUO/AK8ybZhZt6DBn2KFmNt7I9vnAuHbprdSbdpJDIxe0gdI4Rcmr50bTm0U5YRNxyHsO1c709Ou
AUrxZbEONGE2qGRhP3zZPZvWQpJohPn3nd4pl62wOB9rpucAhsFN79HCD5/gsr8ufMOJvKYmO4XQ
uSyGFZwR62Wx+/OCj8PgGV9PZmM25l1LeWbzHpKlumxpcKiPgt9inmOwW0YkqmK3FsK0ji8qmUwC
S+dJB/TGMH8SPfQ7gqPu86lOlUEqjjxxPM1Pgjcg/P3A+j/PTN2ApTgP35SCEGIgJ7BHVEVnEIiY
77Gi781dMkp4+HoyllqtsxfgUrLrnRUwY6A/EY2Na8YW0oXMSZxxZ89VgT5B3CHIshoKH+bEuSof
27xM61xasLvCR1qD84Ph0re3M3A986JNdIb5auhHLF2xBNn/KVpgo35/boOsTqrpmv+Np/ZTDOtJ
bvm8eCSuWkv1++Z0gp3WVkMRG6ZZm9vWXThep0xBVkizy5Nxg8xHhnrcvjJIyd0ifn7xp1LCSoac
UAk9vyMeHKSxvjQ4lZEu2noRKnA+yXRD2E2c7tIIZml+MLmzpLCSfyZu95+0YRnQ/2FsD84RXwgl
ME5bmYIC3sbjaDOT5bbOr3gWyguKGCjuOsAKLr2K+TnvEwrness0ZLhefMP/aamq0rDJp3un8jKf
Axh0AhTOdobx7Nk6xCgmJQ9OrCoaux9Z6haIxgEA6XzbpRSDJnOe080fX0m1jT3X1ZDqenALbKUS
XW+sOX4W9/jtyQxOV4VTDApuAFXuH5Kzj82PUbzIN7FnlcYsu0jMWDBTjgjl3SZeC7aDMTn2CkBW
jukx7j3qrxmiFTrguUiDX/arhFzTcLxjwZeCLFDUB+YNwe4dg4Ga7iSeXbtTlw9nb0S/r52i4uco
A6cQViSfuEGWwh3OfwtS+9m0L9lBoP/CWqtLlIhGQjLmWDY3TUo4suVtV0QCh5sm0rLyj+p3K7+V
+KLkKK+0Kv1M60ZZKd8FllqRX0ZD047dYuPTOdyllxkI06T43Lepd01nkMlBWnbxor8lOl1Mo2P+
wz4hIU/cfCPhv8OcuKbAS26zUcJsTJxCBDPoigmA+bG3SSLrbG4V6egPrK/2ONZqpZFVjUX44Gui
Od+qsyQiPK7HC4WpKyNArddCG3XXTF7L5ZoLbZJ5y0LwesTaKQHVmUBYHtBnCTrrnN+8cJWG78qK
A012WDSpbJWhnD2lVF6W4NGLiPH5lPg6Ll3vt5j4ZiAVkAJoOeVjvvz3pw8f0zb2azOKq/0LnPGh
MtNTeM9+ZWqy2/IF9SvQEOxqF5TyOnYOYZYxHdNCHpXRw3veity8/M7QWHbr/Fk7ZYMYgKpL4Ym7
IQxVS517PkPWBMEtKIqhtouqgkK8lk5JwFbUrBWeDgf4Znz5Ldrg75t1BAGlJwnhTRk/+2j9j1YC
gTWIj1drtASo0/dGd9trweyI+pRGZ0NZVtCC6EStvITn2FBtZ61NR+aJcqSz8TaEvGkEGkPo3BSh
DtzYrTG+e7N39ccN9j7ikA0qp8F/3ZcVKghVqm+Wv0SydwLrTYZ20ovTOHeeTKsD46beGwK3sOn6
dqKACXrpvyWYo2GgJcO62JNDR9sMgUphLNLRz7YGuMG+SoX59N1DvVldaO0gPdlJHH+poGcvIZm7
A41+xGSnQXODRszUtBj4ARo9vm6TgQLd0IObqAAgRtap521i82v3zhYdy+QuH6Y1bHaTWcJwJWjs
9/s1NR1tdJwoWuklLaprx1bzIcgoU3EV748FpmglnQBEuUHbykdH0HIOwU60JSpgfgGEqKK9BdJD
UHqUKPqAQfWy3J2fwciDvZL53odXZ+J3ba0bxpselvEOcoA9TuoQA5Tb5Q/bmEPK+aVauOXnHmHb
KTKsa0k+BOggLv3LX2gvBtHW9yAchtqOPVcXQXpHVkWxVy9jyNNBqYaeA9kJkE8tGXUSuD+sFKc/
7oL0ua+J7kn+c3sj2hw9C/FKXM6Fl7uHM2K1zndF4V08dY6U3F0fV6RpdQVj+VZ+ILmjYNUD1uUK
8Tmbz3cpxoa3Y/NL2CuuuS4Bams0i+hG7SdnHw1PY0nVrCFjPNN50RbegTP6i/mIzotdnecsf8MA
5y4xP5FUA5hjjsCThgJ2nSxIBSEISyCkvcoqZ76zXVw205j5C7m8958Aeh5rz2W83EKTqdk8a74z
pTrf/0xgD/Hs/FO8GQuS9nvfRXtYpfqP3RZMLqChcq+9LB2BvfDIwBCxsHIMVp0sqQcw09TQym0N
Xv75jRsvNNc7KQCXpqH/0Ei1+mqJQKQWPGg1X+79l/NAy7R+S0wy4sjpNDM2Gfag+rhWg3XMvAkV
6tQZXiIywyzKzGHXve6MiWT7e279QkJso+tr/Z/mKiMKjpmrHfPQamkR7bWJn2JjLS4OqCd2J8cx
4EUc0fpVmVDtDorwPAHN9U7zISeGtGzWNpV/MNy6DlnbBxXomM+IyyfqczXOtPKCSeJgAtCNtQyy
ffXasS5seEGGOxghyzTR5sQnlBlJTFQOSehsJ656yE4X2mR3H2II6zqg2k3N5jlWrBiDzI4fq2US
686RIdLi9fHMQztkcV7qjeJQkvdei0iTi9ohHW313wjveU1PG6Iyqx4iEvc1j8MD/GuTUp3xDCWU
gWqIJkQwCXHm9/c4N+iIQwBDdSusboGac4cfv+HnXsGdNzJd0RuFElmbFzCZjFH1PIA6KznE68ib
Anuf80jPWOg4qbXHnCYICzzDCaCZ2VkLvEoq+GhLpsjiMKOG5TL14ZsWn4B21PftfNHRGZGgFfm6
2LuyPISGdxipzw+9bwdJOES3q9tK0py9TxGsF3fpzoxWSr6Tp63hHb7FIBLm6dfJObJR97CY/7Af
Aii1TYsN2Ys3JioCn7OQg/RLbckfbYco2gsI2fzyt72Q3OdDmhCgkImt6xx54JcypwXiaOc3CDDP
eDJbPL9dgualxyS+jTkOJ25iXr5MlYQYaFMw8SRfCKd27eAfUILZvVK7syZReY7IjEhxhHhDJKmp
pC2nncpSBVCqEZDiMD4Utytbbe9uT+qlgais/bkdyAesXisSVUpi7bloE9ieFEnUyzr3wGFFTKjy
531hP0zMTJZjSnX9BKa6A1Et5bOadRaDlMJDWYCFyeF6nBDgViqs7R0huQSRKxCF9gQ7KQHjhd8U
bRm64bZPZih9MLCmPtc2Ib//VQ0J38Vh8cN5Q1a1CA8CRcigjQuTI1tMAPQx/FkJJhmk7yNRmwlw
TEgpYfhcD/G152bcD6HvWxmFtmfntifoWFdKcJTilbT06mJPRFzk9dsO/qgBaoaHjEG2OdvjQ5Vh
qkulOo5UpebHGt/xaMkRDYuTTTU/CUmrrPwtlF9YEOVHPLFJoXV9gnfZV1ZSHvd1+pT9ZUaxljSz
KZrUX+HK1NXIHWMap3QB3TOx2xm7xBFQYg1Z1p8/bqPDkLeAdELlLIIq7f22XuPUQvc6PPCd72Tk
Cqvg3Pwn1O/rOc2dyVCf15m7Lx0v4k96V/x0WopCi7Q8UIPVgPW7jNP5OK6HYxZWgcUKVKMc6Zap
jb4Y4hkZrtbZ/W9JL7NdAIRtwqBmShpSr0i5bv5XuJ+nB38g3T60afF8mDwgUNKnvejZWN6YqEnC
rqBXZcfjS3S+95Dm9T+7JRs0QhhN96JtRA/lVyLFCdIGzYVzkRMBCR9qdEO1gw5a19a6RGKREOaN
WJ16NYojmRdjiqSa++cfaZhFX+wsnVJJZORcRTuplHjIAxs08AMIotEv449FcisfHKwxTnGsH5uk
IrbNRf6dDgkkTVxfEwQaHpzq4o2fye3rxrnCbiqWpJUYXk2KHPEnpxfiPI2FJXfJNQi2pOp9Zs7M
I23WnHuCdKp7Uagl8Gi2+JVRrxeJtNWfcwLmmG2w8jcYmn6VYgyVnUVWX+3QEUtcmlL5enIAK+EH
mHULLEMrS5FJiGmHFNWs1d3oieWOMD2dSI/99htWNFfydDGd21B3Vqfi4FWXmpoj9jOMLUrLr0gB
6Vlb7Xj6O8yp3w87Q4vYuuqxkXS688fKOMEm9k4uHY31An1vzBkmPEXCeSEut1ut+nEXRw4vIDIp
WfSrXy6oHRYoMTbLSY6mXt9xsNC8F2JJyruzAbl05xE3zv/x2qJ1ArJSNjlwh2cYZd4P8MqoLELa
sTkRvmV4RB7dqbk+Y1GdDd0X8/2xfWuIdqMdvs1NUzz326CmIos4EjR/+52gPUbq0dt8DeB7LJr2
C+BRrdKaNnPSoU723omowiVP0EafFokhdnu5VB598FcBv/ww8LkTtnRg47EeuFRxAZWlFzP9DCYk
XjhuSr+xTNYaOkygd9RYKXTUMd2zU/A5HJ2Fe+Ba/KHC+IzLpcFeH2sXkwlPqwBRf6xWjE237dlP
PUa328oQF/G0DFTnMlqtliYY7WJzZUT15EA9DyWjWCROajTdbhmhPCqPuOjBcvqP36D4ZaO8qoj2
nmbL+lcVu0iVRwFZPMz2ErzDHXFlNxLudJ4HqxHCmai1f2lrwoz6lP79KbyStlm9RnW/G1TywFMm
kEr3DDyGCQBqWgNd/8nKzp6moD92BE2wKdTOZGrWh476SdZcmJrQpUcOqpc8yO0AEhqlkqaJ9N4h
C+4DF2Ghdn7J8aSE6KVDsnEAwPh88dx08X6IJ7VetQSsx72fMK4qax24Mr5YFaON4FbVDwV7wGxt
NDZUh0kOiH6HaMe2WgtkuKzJzJBmOjwVV3oTTwuiQIdQVcoYKvIX/ZyENrRr71cbGermr98Cf+bD
oOG/jDQo/QX4x/aj/HPJFKnvbjyNPUhxc1isacHrLZVD3Zh8YVkwvtasYIChyP0l5EFrnL4HNVw7
gMscAoHcReiNcRHbVm5enuT3fRRW7hRgUgMRadYa9TjLwh2yzpxtN+OzPZpuMph+WQnuPkh3ZWmw
H6eI5BfnAzJPegMXpVEjtnvS2G2HRikRZhtKJa+wtaD8FfI40jqseaPtpni2RmwwIGmV3q+ghHVB
BfM5J08TWsh5yFseyRi0Y2k6rZUTdiAHIVoW7V3W3Ey/vs/re/W7qx1YWWR2bOGrOodxQft+9ZuS
fGX0j+2eElg/EbCxOGlpF0B50iwcDwcLOWlu8LGrVwgHKwKG32pmnYriLb6RgH9xBBNoJhWJxZD4
NsHQq+GzYQBfReUY8CMI/rJ/of844E4D/NYoJgrK1zbn3u1rUDAP4zntKz0tHyx4dZOUVks8Jc5z
49vG95PKfOX8r6INGLzb4lmRXQLjaAWU5V67A4eVg9ocxujEmmAGGatfIet6YQ5QjyRLir9cm1U3
4L3g5Y224X7K/fUkSc+hhoj9RiC4jaJPPJQpdingeihvlqrjORqquyWRyy9yL0Spuk7exiIrMNNs
ePtDd64Qk+QuZOXw/Dt9M7GBIyVjwVyo9UMhhGm+QBRXjirKljshvX8MjeGMkZl656zB2F8hEHhf
0Y1F9vRSt8CdBn5jGICWA/k2wXISpmz2/lJTCXwpIaevrebBC0INeUNBtzM0M5wcSpamWVMTyKkm
UJimermVcQF/pARVoETJFoq4D2R/xSEc/MlGHfs1skBxMzYmhY5Sffg3WBed+1OLTjPtP/scEIBQ
Li4k+fe7VkekxUl7UCzdHgPKqn6IvhHYIVkZ8jMi+o6MJokNoIxKYZ3/FvgO9ThNh7wThJgRzaWP
CAbCP+cG0UIXUW2ox6rBRWPY6ZEzOzKLcW+ureRRfgvSGLMJMRbLA96y72vK7PftUAfKCqzeF7RT
zp7iAdoKajVqs6a8CNv9ttAA7fOX13OTUK3LKJmek7FceatTuGen1tQMo6iGq/Sn96vLVZrtLfrp
C490tyQKggMMhBpRAezZZOVHUa5yjd2XP/fAtirjA4agVIvDEiHP3PVPm8YXDijcLOACFMoFfKRY
2xXQNxCqC5jq5zld8C1738WZ7ZUAyJP0n6pj0UdLBijCsVgTe3T2P7mPflaLvnMv1eWgdLQnGt8c
e1oiwO+JDkKVKV+DBN/7jGvdUJQHlJrQ3GqlabYwIuNq1KrdT4CTcNfRER1XxTs/2aQcs9RhIN94
xg4tRX+XegvJeDDHsidBdzX/0dfMOqnFFG16LqsXockA0GAyFO4jFXbOgCaWWq4vJm9EITQ6BT1h
rdp/eNXvhH37shoB3qVxrlLkwhfp//MugI0yRjRy3wV1sQtb2YtXj5JDMLcaC3azJuBZzLYo5UaC
J64NeVliJ1DJsOz0Mk3rpGr64Pe2y64o7RDOh5RfifdYwiGQ8dQYdNLZYWnPSnCG4kt3Lmpi4TAk
wXXSrRopsAM1w6GxhsllDsKpzgMfI6kvL4BJGoLLgIhKZ6RFkiZ28s46Zlvhogq9sEQQ8tjPJ/24
edA3u44n6af+OzaXRXzljQB3/HzMVBZFNpd+djupBYIK0SE6fHvoFe7xUNQ9lTpLASUakEdyEC2/
Bf2islDFaAbX7ngnj46AaDOsdIu6Y49h3mSzZXcTAfvE+Cz4f4ui0oRoOh7Sw8YLDdep9ZkdEdYW
2A34TzW0M/7t7u0DFKv7O8whxwN80KcWrl+syWNDf0e6Vmjve9U6mKMHknH6ryU1zPAFedCB4tSx
ch7Pt9oekPs1EQMg07SA9EzfDdgtuKUvsCRPzEwRH77bWOAjhfTnrfKJeZb7iajthgeAKCCdRbni
t+uxPKeBy82017CxZRiDFS9CUYQYbyzOibg1CHHvS94GKKqFGfTO6d5wqpGcpJzH5mkykJqRiKm9
hRHKaZ1lzPAnF8D2NwbOtb/tVklTcZIY5UKqrZvkGaxr4uVGCsjCewdA9OGGjGIuJbre12eAafYa
0SREAaAqkIRQkNwq3B5NCQZe3/7AsOSJ/kYTkUWloBhpLpN+OjftQT1C7kNfQvHoEvurPaI52vnc
62okeqBsyNQRvLP+ceSbt+LPYpkLHhrNksbSJhDIId/Bh815eYzvXG+dAqf0MK4QHN/+TlkSkviH
nYmzRNGp+AS773ZdIVshQtSjE+ZuA0tk8HVy6Slpsppzv73YrHGmC7Y2rN4mMZz6Kt+hv6wiSSn4
HLpVT5u8uSjfwnSzGsvdZ8qdxPAaZMTGEsI8i9US9c0zLaP0vvwOpAEOmNTtBx32rmwz7SWEiW5J
xYDdAN5ZMNEGupUq9sJI877z1OmSuuSTDik37EWb7jREUpxuRfcus8c95Uptx0xt1dQhHO8WEDI+
XROg6k8UnhEk15utA8IKttuJwqM9KNsuMAumM0kdpjpzmygdzmG7E9Dn2Dt5OS/acdCJoFf/KFAE
sB3evG9tqKh7/+SCXTH5gpqZJ59dUPHILv02Q6k0NVYagBug9Q1WaaiCvqgMs0BTomeUUy0aJ0F6
Dc+oy82/IGCT1aR13+XCNNkesS9+QRrhP7y7FV5bcdykUlxmVLx20EpGIPsc9g/2KRhkD0UTrVra
H0ObRsuLqq15v4rN94Lzi6qSku293y8qt5Moa2odqYuH0CNQDN1ceLczHbGX4Q908Q4YPVQADf72
UommSOkvMwNhR/PUKCl02yjuCAG/pREs4YFd0kV561J9QcaSFSGVBdpqntaqTR+xdOwhWgi4bEhD
5U13kfUBNrOd81kpWlkywbCveblYO5BwCKIwRlWsLJDFHbrdLxZ0+zyhI6PzznJU9U3K6ptXjybB
44wnv0LoJCqv4U/pwPOewH+AyECTr6R0fDNEgy1KnJCLNi5/QjwT4ecRLnszjpvF9tWXj8rUWnD2
9ypTECIM4l0MDDGKJ3ayJCqRYxaMJlZqJub4fDR4Wb/YQ1wkImqSET3AbbqrvjN3xbEgrpFm/TB4
3Fw4rW5q7tepgLs1J0XhP7KNxpe/Io293taj3XWMhstqTgX62ARGz1LH4h/fZ3QIdRuswvdFMGE1
d+ki1QqdF6aLBF2IZTzX6Lj2qDZhi/CLEKcsac9AWHdAjGyljON/brgCUeyOoqdlP+8nQ1hTPTo1
sMs+i7XG2ciOuxKYFm1GOBa9KSPnAfMxe8oN3YiWhCygjKvV9RBKqMcu8iJ5eD5kCZeKN9SyyZIy
jxOqU6wFz1cloMNbYvfcl5lYbeA5I9dOruoxAw+NE6FRGtgaFQzuihUl6SXEAhyz1WgGslWyMpul
rwUhQCYFL07BJ0QgV5paVleSEJDRRc0b6RqTvh1U7PnY2hHQv1o95VCDl1om94yvrvDTIjN43k2F
lR1lNnBMRkygo52l+lEi7cbjLnMtuK+kKbGY6zDb1f7Ow2/taZPNPUG1GfcL2wZMm+iUb8He+sSb
GyMM6f1By/VlJUR1v4ynvs53/cqvv9hzV4cL5x741/NVPrt0QhhQW32gM+UY+aaIdYNL5Fu0zJSn
mXjeXlV+8sZMdVg4KhWbrxWAXH2v4ZrG4Z4d7pSaikrVfY/pGVoDdAU6XS1wE6nGDzCpOKMGFfiK
3x822xsh97L7ULAHoGlpmTAklr5VRL7wJuf9e/qo9tSpZrMaGOGbPnhWGMzuCi8Q7vj5tn6cB8Y4
kiJ95ufT22PB9SODnyeEt/PetTT5P6Ihy5+THuoDMhIG6gRVhlEpYhDryi1eRN8jAeXS2cROmYRj
xdRJz+ypU1NU1a2iBBdNUjURx1q+tu9ljT2X112eMeUV9zMgX4yZA4Fe5vR7Lxi5Jy0uukdiXaEd
tuSpSrnUFUaVHVdXDT/bmgDrPiPEoHRj8AqoSaX8Vsk2g/nEevXVkOMoufKy/EMESPUhYH0JC9fP
QRdE01wDgdZ5zpwazzrAe6WIpU7pMpylnn11OCEoT0i/D9Fb7EtryOvuXGoDQwwSNmEANfjlwZGk
/HSR8kCnQJW54HK1HCpdrpv59ZxiBVH4XVLzLaER89vKYU6wgDZUB+87y5kPG9xMMdx/41oO2qPJ
6/WW1X+SmfAq4U3FfeSSwXnadvMwcCNL4fuBc7dN+HlkmMBvOu1AJMzm80rpnIqxrDbEhUykIBaD
wxXdAkdAiwGWRo/HWB+Zb8opZn5Uzzkko4PKCJsOOpsizkxH/utK2JLjg47T5sKnrwjVo1BEzOT0
/XTqmTI6UtJqDVx08ygBEFO5J7wRUDvSsK4xAuGFGmD2SGdegZ0s6/ZFFXvrJL+k+zzpOLFrNuS9
naHCHtArFBMWGzHH89gvtViPInm3LbV3dN21EYSMbQZhG/591ZUXPmW0ACkUiqKmNeGvIytKamwR
uNr3FO3SguVbWcdKu9uWRGRi0llBXobU7BVNLVABhKGjQWTa2vmcXw/Cvhurhlk0HZGUcqvsuBAz
HTG0pvgKwtd3ba2drvIOffDJvSz1Ib0slJf/GLwZHT2TH4xUHnesanjAVmp3WI9MjRnAZb4yhEtY
IJRlY3GqmsAfC+xZuOYD0zeeBsm1rkDrChRRKdV4vMDIDE1dCtCpg2ll5AD928ByM/ifGQhGj5T4
eSxPw7yY76aLYnP/EU/I7n9jGh/olmISrUsOU7RlHaCvvBCbVwPCETUtk41Cdauw0Ov4rCT5uLWG
i0pNDddgAX2CTdaW9PIYNS5ujkItK+minfYW5zu293ToiqxIDhpEkvR1j+ZUqa2EA2tTu0SQFC9z
AKWC//X2pjW/4mxQRZlEvgs4orJN8c77WgNMC/lQyagUC8XVXrnF+wl1LW06UndLzCV5LZG5g7AK
FCHnEYoVO/PbQUZ8xWwm+KEK65vDhnz0ssR3XNcYc+5OyrY5tDUPq34tHS0fG6vx6X1niZJSR+Dg
7TaV4GpIOSuZuqr8JqPxbBEgnhf4AgadXKqIBmoo9bsmt98tNveuaWBeDmWfzMrkppxK8lgpR7FF
7Y/u54oaUQKun4LTm4PGkJChyZBpQu9CEKn6Unq9Z2Nbx038yK4evkfz1iwRMXdnqTzGHcuwIy6E
wJNS/g2YUl99w9QHJEwYg3YVG80Mn2Tv3CoSuCLCWZt/cyidwpDRb4/rgHW7JQurctPGl/mHdqKh
t/ayImCdr6zpHCUbhkPuA8z7xyfkYANuoj94FqUkAWvgTNgp3bo5yw+yzMDZKJHb1+GDEAbpLNac
JwoSF8t3lbyQjsgEI5pMx5CR+qlTKu1A3a4mqiPGKknIlT5sW0bn/DjLn10j7S9KFu4mTqbhoaNU
PRJ7fAD2g/n/7umlfmnR9PJNNJuss9fGa7qTrIU9Bb4MDaJu6mKq6qlIBmftAGLIiae8++2YsWYA
Mtdw/qvfCklAvlLE4HaGcvFYHH666ySRSJH7XQy2HPK6v2AcmIncVgZcsfywfh9c1ipzx7D/SqiJ
P2yl7kRz2k2bEhe6EhVKAkm9K/GbWBx9wn0KzDF+RtojyG3Y00NitiFQS03Ilp2HQgvoKCx1dHNH
0UBpFoJXYAHc3I8TvGb5HkS2XYTGtBaNihLsrZ4HdZKXrO6mrEVDT/RgHfkJngU7Z4b0EfHveOLa
Jlfc1QRKrDJPfgAAOSu45y1enuydhWQQ/wOx0WpB/nidnc4zHu5436vv4nbe0s/GBTRl1ERSzi5z
2cXS+lXKeKgiH3TA99bVG8z2yEWwG9vbq/+/T9a52A47rstVebi1gMjjhWx5uVXoG5Cg5DklvNgE
S2g6g3uZjvdj9CKtteKn3RBVon+wVEhHJq7bG3Y8quHd/xLRjJDZJpEpNzn6rv2bo9vlJw070WUq
uj/vkxCnJTQ6YL1ZX8u7sLgJpxXcxOOFdnNv+rNQhDadoyQt+crehdaGp0e3zyYXkDB9zmb0CMcf
ZcxagNDPKVuS960YHLTPShhpS5eT3to/JcehJGZ71X35/w/OVhRMDClDKU7s0OWXb1AzLBrgXh7U
CIaSpWs+shOsyEwcXPk5fpuz9q9g+P50QIaP31cEpKadG8lIQoTMRpiZd3vH0Coap52iMclmCvQl
6HMBzBNVI4IRZLECqDtoQqocIRgHNH9zWG4m9QylnwnwyUnfGr0hx7w0kj/3sy3lMdApG9LxqE4S
XKovbOHU4UR8avRxInL4k0aLvv7KBh5fwDUWzlf1o7cE+g4QXBWdJ7Em3c9zN9vzO4TDd/GV0rHm
qHI2Mjy+oN/8rCi3ABD9eYRUt6QBA92NuvEUJF/hH/igoekFTaa8MlEjHmB03cUEFpHKogmsHuAQ
SDoO1zBkRWkeVyv5nhl/ara2NrmFPt814QIwBz7x2M+ykqZZzGKL4ObbdsGE2XW0X5/XhgPO70Hw
Yuk8xIJTObBppUzyz8KMcIuFeF1Fk8NJqNUhM7luknIt9F9hEXamuEXAOxmNSPf7Y11S/M3rcq0I
KniCwZ4s6byGbfTdBnvM86QxoSO+vlqB9I4I02cWLH9MMpb3zO91On+oHtNxcG3Nzg6nhypS77B7
2M9lsAnuTVe7XTdIHuk3dYsQ2MwcUKpGajnoHdqXVY4VqXZeNjAXJAtZKxnDElwxru2j/oQbh1Oz
qvdHv+JleYWOZnQ3j2+kvFr/EQTy907kBuj7gvfFqrS/ll8rTF0GX6c3wC00ylyKtl+NCIzngFu1
bbxrPinK1cmgBzbWmIXWkKOWMNxjDYiRfUWutGFyPIAmpLkgOvgYsi2Wdichcs4v149aFXzgrW7z
wTEJ2gL1QvvArdfix34zJ0juUKMVSAzJ+v1wclSDMADUdOz1cblPWVC9XKZDw/d8p+WcZUqptXRc
Plrwrf+k11UuCETgDZvkTR0+tGyyBQGAlkCnUt+4lOJ7oEs8fOC5sVPqa/0gFt4uaK0CofWrtS+C
Ef3XHxMUh/Ed3uYCO5mePwbp12oNAAviUZERENHFZI1HKlkCyzIUSTkvIbVyDGiSN3XbiXuQLNO2
cUfvWoUbDif51d2MZoks7mAt1ZVvGxQUUFPYqF5Ax/fSDCIJ05BU1Zj7NToXANEpu5Esqt563vtM
M/1hnGa/ri3l/6XfSnQ1XzYZ7XTEuPwfBgI/u6Oe7VviQ9PYfzNHJt0ze1pvvxm1GmKIaxr2Sr2f
tfLruFxXJ7wY1iNcnni3+o7aa2Gi+DhCUzTIpVmgpQldmR/3XGPATFI50tzDnWTBupBv09e+50zm
OznxHBAlWR/j+3m3KYZXmSkQWyWtVIVv47HCkhWL1POS9ofSxlWjQD8SQSfRN553aFuXRtijY21e
T2p5giXatFWWUd2AzASYYW5OIzBhUV3fVxou9VKwWFcIMkschKue8FW4TSJdobQqKAmfCFVUKQ9x
kVkZeqBjwu18QMgunVlKsW/Vg/0WfI1AbMMpSdioD10lrxHTc0RaSASEw5w0R6y0IX2f/76Dgw9m
G14JT33wIegIG2QhaH0mLE9LT4RytRrr/0dMCkiZAI1sbJoORayMWCKH2KcXGLWAi3nnhkslTgo7
4B/VPbMvtzNsy9Bz9WJtM3NQ93F1RyY0/Uahx2Knmgf9/6mKwAZd5qOjoeR2VyXwxnSMZ8OgTvDJ
Cl9JiNCQTRh2adfmf4m59BOsrj1JQZAQFFSU0rjYg1YJah9TcLww0Lk3FfGy5e4sHQhE1PINFNgP
jNU15HgBViV/Q62ySFr/AmaBATvU7aY9qWLXD2YP33DblviW4TGC7iZD7suXyF9slElHs2st40BZ
OvXHA3L+cepsVj22b/Xtd9jYc8tVxA376HbpTXUDAgXJSvvbYy1OgHMF2nj2fCdvUWf1gJncGE9X
qZpsPhr8Fszw/OiCiStRtLzz12y4berO9iEtyGK0lrxDFBq9KKKjE8XwU2740Q0JmYYOSHPYehzy
9ezq3GWRgfksvAggChRgV3IlJ96EqORpl/NyiqoeScUhE5OnNABdbIge7T8ZuJ+8KsqRKaMJa2NX
y2JpFVjqpfYScv+MGLCeE97ZcYqDDs39tN859D0Vr4/ISeLoxOeP07scxHyIjh2xQ/zYduV4kDMl
gd6m8LWSCaohwryKr/Tv2K8J54MNxcczZEM1/3p1y7LTKOvGPhGmVIj8Oswq34m+kKKcvJmf4jzD
L6EOwq8G+ETXVQw32m4M9gKPjg4MQcIaIzz1PABvPr66K2SpetDbt611ZNYG/yz8F38v+d8+ruly
9OmypQxikE3gWGC64v1Dp/up2sPviINHGXJ1ozfC/7r6SCNsQs5Lv1zC3o/yskIL2L27bWMF4dZ1
QcuR6//yJZ+1rkMP5ZCTrTAmQAEiUaIfgnx+UgI75hUOn0GeA0vKyMv0RhwFg9UQv6LhJugOrtPm
yGa3OEaMv+KS0TJkJzVuAJVce2uhTFJKXh336Xu1WytUV9b6NEsBbK6pOnfyDsQArHBdLjMgKxvw
N8ZE5Jibxqg6zFvGZIyjQBtz8dEpn0RrV7KSN9FAO06R3TDhoh2gWAQvef03m+yNF7Nx8PigK5GO
YWVEzs52B07e/fy8nX98HmubCS0wguVofcqoUAeG0DVky1dTNC/9GhpGzKLgNplvy2+fv8BIORsk
zNNT5Xf4ONalHuUhcMYX2b7eSiwuRCmt4zUbA+FE+VytAVzNhDiag5MChPaic6Ejrnj2cvhx6tlp
8iS1jKLeMbfsgYFAAF+aWIoAGKNjq8L3/+brVzRI4vCCTOxdon66VGNRignSKqCWoZL1kN44LNjB
13gpKwBDnJvgr73M5Sn3fZUqnnzG5bEUaOe+VqI4O8iA1SSHXsfpBjhhYXHTO/YITxUitferhRy3
C2pcsfezwPNvra6IpV88x8gMQdHTPENlnX22nLWDELI7RJ0SE2VykydwLQdC38mtU2x6g0Oi6rbg
Ky7c47PYvVLbb+mkj3L2bwbhB7uRohjv/sYoVmbW/nD93N8ycR0zZyhRUSKY1GJHiEC+8vHAFJ+A
TkWy41sHFN9yYqFHtQEgS7r2fdTFp0K3Q3LOex1FfDLrvz2cFJIS5VRFGH26RZ4+4BtRcB1/SrNg
0lDqRGJ8D27wi7t4189yuj2UG6jE1Y6DguiV8185SZM42SRBF3oq1MurgPPGBcMXpkkH27RSNxfB
NZZUV55rbeTmBZhT6Cs2cXE6d/dGZZw8ZMxLjyRMkYaW65MryJfgPD/d6EJizgDMNOHAYTk67fSy
ogjQhRHApGzLCvDSZ8oHnlc68XjAoHHulNKx0DzBoCg00sKPBx4x1VN1zeS+4PmfTE/gJ0vIl3hv
rZr9sMQe6IxVxRaGnb9CVWpTonjueSual1NxEroCd6GW/1Rie0TlxSxu1P/cbGYphXLZaNEp0h/x
kgEX9EjfNJdnEYbRCa0Lf3afwdMyQfUeDa84QhPQZ69vr6+F2BgYqjL63CPH47/Xm0d2Dj1TJrVb
8pNxOwdBbQpYaAMdEmB+nUQz2ZAtbBlNAAKLHpX95uGcfkOQfyoK2ZV2IeRltC3Qhu/iUppz+g3d
2gYY6SrlzBl8hiksA1HKFOnjHjvgJ1Qo+h2afXETJDAgz1XcTpiLPnOJeS3IA5QlMsdKGeOLepbc
m/t+ypnTp4KylkyhIhSA9WkCH4i7VCncAbLAtKBT6+VLU5xSasMtLK9u91Oim/0SSsY7qNw4aZI3
OzzBPlugbDcz0viRXGmqGvUZZHozxfXDpjeGF12daNLYvsRyFmKavH4r82B0ZKDkTksWh2ijQoPC
GJM6ps+iSu7CI5wo0bPhmzc5P/eRwfYrVsOnEm+1KRBfWKWehTS9UScAY1SmCGJ+k1p3kQODyl73
PPcyQ4yW2f7DRpiQlZ9nZai0ayzvEcxY+dRJ6cKoSFxftbWPjRBpav4aiUtjbmaqbO9EKPKsw006
jVZfgOuuTByTsKhFG3VSBaibQnNdhVRdTzBCcvHs+rjaQgyggHdelrHGT3FVWkrOb/0SEJvfbB0J
7xQk7O6wD96sjK5JV9Rrfyjv8kDVHdjW4s+BvHPq71EIgSOIMEibL1m0m0APhkY8hajRL2r1JRaf
qy5dTtnHNIR/t/GQnntdpiG7briTef/OIIVjvwo84pKwPFIaHx8N/puGXT8KjJyqN23WQ9DXhuZF
ksrr780zlwcXOsHv9HO9ZytSArH9MtoxkUp6lEGB+VHGwNL65VQAeYRgWrasi4Ys+G3dwQI/CaIs
yVya4ifQ0S44HteNQz/aQbGagmmHKb2nWsRcsag+644dhlXrEH4xIF8mPhXtb8aO9J0own0RH/9B
FoSVS3LwPT+NBT/qtr6Gcefp4kyB5Iaz5nyCGM794UUtMBnEUYR1pbICDZUcMtIaMpcuR1FlWGke
/AVMj3AnbBFa7TspgPM4tA762O3uaKpn1LLP6j9Nuo2aXhvDLSnFheZSnT+6axupSQLQ6JA16+IN
OGugpDlawhm6m9p0rDSl1SwIQDEYfJzsaVDdc0U74SsRTyxx2dn04kW2YVOeeNXbvwXmDaFSAKF6
o2bKPOyrXKR6r89Ft1c9Sfa1mFNnrDf7N2Kt/W+BhM5MHOFn37uT3k/zcqCil790jRo2sRxTjQM2
WVbeN/HoOyoJ1tfMKroiZ5JFTod8wT5isw5e5VTkp+eBcZuhCb2uGkCu/TH6CjpIdOF3EdeER58b
ZSUX5fjMscr5sVRcIKSE4bvhPQ2azzrip2jegPKFHj1a5m6cmbKHDoLc92+cn37s+zaoKHP7044c
a8FkfjXq9/SVqyYE5MWxMZ9IG3bCBVsfm2j04kDkV/1wnsB7EhLAmL3LQPNVNltT2A9CpwmUgLgy
Q9Aymq2JXNBVyGx9ZlbYAb2w6lsztK/rwMCWz6zDvic1K1c+eJdrLESTsmDLpaXvrFB6UKE5NLjM
BpNzzuL4Geabt+/VDBX9je+Qeb6pM9p0PaAvaiKPsEK/CRhhDMVEb6qVgs/eLy+R4OdQQfh+p7uq
ZpRM7pdezAU9bjQhH6aq6GX18WgPLZiDqqFR94tW+REAjAeiMnlsbYAJfvvm7we6d4QMW3jWT56x
8+c7+2kmeQiKQjiDA7fwu4SA4y3Y+fas+LYsF2+uJkTSI0njn7wSBeNxVWVAwug5nozQm9/vkUef
ZOUfznuTFLHwe+t/PKXsMIOBQ7O7qajdPrLf7Z7MeI+kMZDsEIX6HeplC/Lrye15UBhpREiDoK7h
6W1H7vbq37rAJQIcAhV48Rh0/saBcGJz0VwlBLHOQv5F8YEfZXoaYPDIFbtUhcyBfbp3oLH0FhwS
TFpd1C5sT48LEGL89GjibJraf8p9NSBc6WPD9ZHrV/G2V+NM5QY4Cnyq/N8EecQwuw+swWKRhvnM
JWDadV9DKUCCSNoh0Ka1EbtxkIV1Hvf/G4TRpfKrNoy850KkWgxF+51tfmU1XHSwsRnFLXMMPvmc
BC8tXeiXQ9j+JGt8YCeE6Id2AtKB+G5VEI3SQ5zDb4BNHm2kN11JDg+P+EVA+dVRghc+XdflO1HK
DwugVjl1i5Dgwn6WC7WSxE7R35dT62E6SJ6Z/fMnjw9wVH8P6tqdKIkIZ5Lj9dLdTvx9L1kSOooV
clnDz2ChnnDJ96vUrbgSsuiFe6hxR0ZTU5EJHUy8Gi3LNslIl+GE3maYH/uRKkR4zuVV5Y8pkXHN
DQ1IXJpX/4dIi4UK1T66JHtYMW5z/HUoQvk8D+1eAldmL44SsApN8htI76wqBVPDfnFMaLa7gXHv
pYeDZ6EdmmH/5bnYRdJXkqBsHAlFAlUYPoQhu+TcwCVZb8cjfpjfIg1haE7R9SSiK3T5xh+SSj43
9uxrmSBRY7L19irvj5v+CkQaMWeq7xdHdyORYojAsVR6I7Nrt4qKNPIn5B2WUH0ZeLSkV2mdA76P
CTdm5pM5I12+W6SRqmK0wZSGdZHftQLoTh0kLYyuQ01CV1SYDarNGqysc2EF6txd7a6pWxtd/9MJ
ixYVs4smQyx1T4w52PN4ReP0pn+0l22qQ8gBHPwE8yAm9V85gPAfDoUKbGxW0otaQ32x0eUxH48p
NOkbGREZpF+aaz8qDEcyfmRz6hWSg7Y2DZtjj8ad4uf+Ly5CcNe49LUaT7XHTd7fM1ZeQbXGgoFy
C4r9P2GZ/pkQk1mJ7CW396h27vM21qjb57atg9axlEyXB9p2jTgFwvezY0X4lPvni8ACEzl+tpmm
wKPUjgxLJHKZlxwZbeXBiVFbMnghTmRDRlynQKmYWUXdNNTUcLYL86V+co09HraFNFeJ+waLELUK
DE3lX6/xRO6CZRTVGO0bCOvrdbelwz6lZEVfzIyBGKgxxXX7ApzvZIBmGbsOx8aS9Cm22yKC91CY
bC95Nsz6uaJgl7zVsw2vFbtSl7gpCngkCwWDWNt2jdmdmvRHfP8Dn6UxXodQGtlhmWk7JD7yl4oS
PTgr+oVWVcJPTgbBvp86Ulzz7uROC9oZrnsZiBDoeT3HPUm4f0g6UhVufwGGsbVdhPIGFcV89OFM
j3KrawG8zYdOWPkg9l3gxyJcvL6AEljQwHiAJBEmg2806pJ/tzRcv2H/CjV6B9Q0uJv/EFTfRLmW
LRYKcfNHAb6Fsm1e9jK7dEWSlZN3WIcXhqxw+704xDTEXeId0IDpHSAt+jnuY7PHjqF+MVewXufC
sZZ4dbDPDT1Zce/FoYlGsLiqmSqvKLEOCQu9aoOo5udMxG5QVHZ2jw6iRtmnF2Vzpu4o6cxOmi5U
NuuzGdIF8riochgwd7+qs/ivNO+ca5OpwdTm17o6X6UmsC8Uox4s39bqnqUc6jnefAhsYl2VlKo9
ANN2AIrZWiAodmmA8frjn7wAjFrc3f+Xzc4ZdDZ2gCnvbTjbXXHljS+YJESHt8IcyW8Fj9oBFhjT
ObsvyS8Y51mAZp7QEekmzvDsCfsOpbcLkhoIcObFQZEzgw34Y9DAeHo2g5S3uLYpIPs+oEpWrXMP
Di0tt6AWACydKgnL2OOPFcGc0eiJkY0+BeCQSo8e30Rz4HHyNHK543W8w5fTbEQv/OIMuF26YFlQ
oCv94djIMZQK9skjVrsh6mBpsfIWPflL+s9JtLYORf6qabjpMcsHfUasQR+qTIH9Nvx75VKYrRJV
FYAtHyXXSrnXqHWvNP4da7r2BdhIa7jdZL6sEOIP2H4iKsmhh86Le/fucBISyWjA1t9pzPnbpzJ0
CEA8MAtNI9KD79ndjTRKmUNyS8dmhc494s+l5SoIb7Jl85nqYHlFeEvKPb+YGCLrzx7Sk8qYL9b2
JMwTWKvbIpkYoaY1DgnlKuZAOsFlp70TWBFKMAIAhV95tzWBotl6ugUGPOsN9pgcIdyNVwBV2hem
GkJa2hV1+k96cYoHGkHOPhQ+3vArcd2hCJTuMGG2HsCPEZ+CT5WBmsMdaqEOREZrOTKOOntQlJ28
3Jj7fVNJNA+mECnk/XNYjjUmolzvi2LK1snuRPJY/pBuMXLsO2TIHEW3wYZa11TWnl2WHD58js1q
/4c5Q6fPdSNje52g63NTUUO0NZKJ/EBwbjPTZGwUxNbMb8+m/Wlas6YC1zudngxI5G2liYbMVHwT
EP2oMQkOHWNTHOCRCzuHaY3tHCYDtYe3XuslhxKBPVrlW2YCvWoYY9bN1VboD7JqxYSyNpy2p1bO
hinBx185lL6pdIMW3vcmXnUuKajOphYlFlQKjvT5nAaBp/cqwfqeNvja0+OyJWqNV3TiFa1wj08R
nEevm4GJ3jfkDKt0kGqlDcVsLOJchl85bmUciwf8xbmgljc3X+HEfLeypdfponbKF482oBavXdIv
lmeLako8PXpFZNdrx9vGfZlnuPLbj4CS6QwjZAeOsljk5b0YzCP1vqleu1gFDHhrn9elGn3K9vaD
MH8Wa6eiMuyj2bZL3E5g2l8TDGMOMHbMNmLA4tT5ipyRA5eblFKe6f5hGffnXPN+YSuk3CGq42h3
LaHhQfJ0V295QUToVzZjq2reEHUArtXJlKzY1TFpKCb2XuqOAT/5m3WhR1nAbe/MGvbjy68elqMG
EzQpe4PIrEkC1f2//CQ9XQ7saYTFypnT/baO34hJzk1pfXgTBIbtbY8KqshR6FzLPwsom7ptE3s8
Y2EviN47lB1uktMCbE4JpPoKGa0ctz2PZqcG0I7gvvZtpxMSAfVcNLay+kw1eXR7a9h5LFg0ugwX
R/sZ7nbf4ZKmYN2Gj84DfuQzO+dFkQr0TcU0UPN/ZtVU7pIw1+eVmRlADmEPB/t3prz8K4zewYyH
n2YB6hKtr9S7gnKtOMt5YZISfS2W4enzuSeXwKZE3V8jia+dS9g9aZRDAr8o4JtcGBSdHkh8Kmf+
uQh6UPjYxNo7Mn6jACIkhjEIKgzKH2J0ffet/5pIbBvvqe7vht76zoplEiavLzC8ZqThDDHK5rTv
AqbG0soDUnf7nRNbY5LkNsFV9mmDAdQcxqXoKKlT0pprEknfb+pOkITVpHEqkGa0H51KwG4bwqZ9
QlG7Z7iQBw1gJVLmcPGwu+ivtMKXGGPTROfroNj+bj8FBUfrCXyR7ALkeEA8SC0IZlYfZJdHHtk7
KBg4Fr4RYJJxtgNj55xBFsMxTdI9YHwdAASgQr/0XXun0VgrANc4kl/aH4uWuZLd4FLApUS0STiJ
OBYzVv5YqgawWLd20OdXg7paoAb8rVQMrn59pnhjhfPqq0aAfKPrDNGk91w6d56m5JYyn6yT5WtD
l+OVqQ6JquhECppI7+FjFM+EPqCfW0ecNShBczsd3b9CdYCne6dkG2bB0aQPyr7pz9CPcF3LL5/X
d5mhTds1HaSSlGMtsBqFLTD9TE2BvjwjjOVMENPLyFlVKCC8en9/N+G6qecDtSq206D1ZRfKdOop
CZuBxEEz3LZAlHEp5M/X8QoI6JLBG34ZXph6g9n7jPyAYkh3IKCfz9DfNg/wehPUrHDISfNRvMF7
SlRpLUMasmDvjgWLzfal3a1t6mIOnn0M/IaEzs59EhyUWh8TE6KjznnPeLBMv43fl8ACQKIKVGAd
griz/rJzcm4yn0wXPL4SbvKtmQQWieohVuFxMIkN7jZGV5Y69ArdRg5b8xBDHJMzvF8UhhPldbKd
4BFqkrTi/Dxv2+J7VIy1cojpVoUNgCiuSZqmuuD0XI6DVP4Z6Y+NwmSq1osOmImBAjGQgmA02ISL
Ww1bremYfFWf5TOAPbMFTYNla8bKmOhAE9i9O7qopKNB64mPt+BC58uSSMaUV36j0T/gPTvysn9n
JjmPga45434/qBjhbclw5OlMUDmtgKlz2xa8602x0rpvj/yF+VtJbmCitBxiurOtYrQbyyfal6MS
apo+4uvmbqPx+QoJdGdJcLV6GttV6FXZLa6+kMpLe3S3+XkZKs3SBESAukkSllRFoI6MpK8lZuzk
6NGDELAHtPuuQxYMeAw8V/NBX1mHpIBnFAlnERnSn4NK85lc9ssN3srDc05V3FLF/h/fI0lSPhiJ
/7J+LXddf4wDSnUYll3aWves3lrfnnlgtKcnmez3zUQyzoJAVjRnsbwZhbEr1ZX8rYfR9EWItAie
0kq4tLyv9JApfqhpcB2RnHbwo1oM/pO4O08yLNL8a9rvVxFebQCygPls5UOh6kRSANWD9Xa3b4m0
NxueE2PcbARDhInW2N4lUOeFHOqtz/oDOWbuZql3eXN0mvQ36EBCV85/nz1VYuGP/YhNBKucvook
KLIFs16ISHy3lyJo3XUwerneJ0zuxy9Jzi9NRiL0FO3OCyQqfVXXcZJEpGiVp0nkLhXB5MSxV9d8
CPzNoIotGNQSJgjxTMabY1nMZ5I9hE7efKD97C1WbCyNFg8KSuX+GJmkm0rqlHW1HPvM2k7bICQb
qDRdFaqUn3pXkpTkfxBjzANh8csSlqYsevRofsWPunzWnPqgLWfYLVMi7bgMqrMm9JBJkU5DF8H8
eLCY6MQ2MO3kjCqy++FQeC43oO19M2aVzJxQMDl/paqNdEzOSfkaRnBK6wWGEY7tGVjRJ7nT6uTX
NqzE3P3VNm9krvnc1qZRJresd4Sz421lmHo/HeJb73gzuA1FFVBK9HytMenDM+FJtIsz9WYSZPQ/
g64vLC7EtmJgOqbXyi72R2hYXp4vWXaC56ATtC1rHbSgFc/k/4HFqvDlBWb4e3NlPxhdniINS57B
J76QFwNpXyONvX5OBQo2xD2tH5pFk9otadVSYeMAukhV5Fah8L78hdpPWfKQAWUHIlDT+IqoC7LV
wzsviDrNnV41TXEl6poBAYSgiIHLzPDQlpLqJBVRVBmCsKHAdCj7PuYg7ikeCQFZENx99qv5y56S
Zd702Kd7zRx9uveckgoaO8VzrVcd1dkKjmalIYFGRx5KfGS/MK+Q4lekl0UwgesLBgBWpFrrKi4j
UGi9lmaO6xJJN726tKi+nNCFpiMImKNQru9evaUlUWMpNg60FezQBI4G7vOEG8muhFObAQjK6Qck
uqtrh1zFG5jNK35KMHHVVF8UUIJu5Iq6xNT8H/4DVIwG4oh4bGTW5Wo4aFANOeL0ct8rC+JML4Wc
ZikWfSLGtEJxutDZFwnmNobT30dHyIDCc4Us07Akjfr8O2CLGv6sSFPWdfAwgtJ3iHPySmd8in6Q
s1qJljF8f+knanIvjulGkhbvXuyK5P2U8O6lLtKyRuzM3qurrORoEwlOB53ZJ/C8jHoO9k52CB4o
3vVlSgc64AaHbfgtToKG+ytK41zLIgx7+bMg6Sgj3dgKUVH6YX9aeyxFpU8IaBNoPDqeH27PHchm
1EYHRYX1O0l6CeWEhdS/Dgr8hhCfWzhyq2zCBzVdl3aXSCZRFjmnkjpOiGNLK9a2yoBQcGfgODmW
2j3QWxJJWjgvNED9/ShYXY8lmqoG3m6IxeW/2BP+ncbg4s+uWu9MCrjqXHJ+9QTUl9M05rb071C8
wYdpcrck2U8CFUwLWhS9+u9hxy9m4gVI/YQmSYaMTC0h9/QDKWJtKuaP/RiI5jD2/Fd5WHIlgoN5
mBJCzHSbw/8IzadLJ0nFTpf9+6hNnlTO2E1PV0QsBFq7xgOuEb3a5y86LvDBzMgOyp9+QLMQKCw+
6cnC/ZfEipnxdKZ44dIo1M7s0+fHs8+DEl5naND1d0V3LXtPZtSfgbmZkoeVsGEQa7qJzR/V8Bl7
9nhx1wxVZ/E5CYRotFwr336arA0xJUXKgAoZ+PznIFhgQkycQspRoC4CxEoZLZuH6M4FLJSoUHoV
X54/DcRRsbtElMdcj35atykF/Mq4oBbjeCRpYYc3TQZGa9NuMpJT+0d/vurWO7v8g/bX2XVV6Tq9
6ihjVhSJnNDc3/plgf7G6RIIU99ScAIpnHvB99N1cYATgihjMJl5zGC27KYUfTJBIG7r/DtSCdCt
0MSAezA4oGtaVf5ygVwLMKlzbPacbLj1e27bNUGmKUpAdNi8SMTxDbKOs/IGQMdwZ8+sxuyFE7TB
epDHX14ZdpMLogzpRiSyPlRQUVdxKZG4LbqorbTRy/BXoQ2zjK9IYYndyhAzMJ6TBjka0F38G1sI
+CdbQVjNPP6PB95DOToYEMM7zy6POhWpz4RqqKnnPtZPsIZaCIHNrqeFy/EW7cdTV5+eV0dvKJp6
Z0NiAjc/UhSfjiOJv8p3l6t9OjjVTmSWfixXB1GZ3Y9ORUuQTCXEmuz6+XDbXAnHfdsppCu53jmV
2kAoDiC9Vgw1gb5Z6094aCvs/LoSCgabMTwSWznyu9RM1YQuBHwaVw0m1GYvVEaycW5SuPPL0kq4
mSMQq53RFU6MfbSAe9GZV+JTVJbuBEB3dq+xia6AKLnHaAl/k6x7MSDgWlzHeE69erajsEta34qv
XLkKpKciik63B/ioCiucGtq/phK2U2C1+q1YHuaqf9hTd1LNJChVDxCKBPMsJaQL/IIbFvQzhAha
wW1f6jrWGlfntkZyqTH4wXNN8JNzN1HnQUD2SwNOVvN8/7PZvP0tkA9JLn0gkP6ZO6FLRFW/hw9h
I1iGxq76XrHQkIXk/sSR0zSE4j2z2tU66BfpByM/UkfXpQBTwZjvoqesdbNguSVECe34vay/iATq
FuMacvJvlzIg43pISzL+ashbWtNYfOgdw4hcUcOk8S1ooNo4PzipiN4m27DTTj+U7Tea62QyN37U
c608aso4HwIKy9V/gMT4JQG/3JSLZ1MdHGYAd8tq7ZAuJ31Q6kFqS4XSgswJDmPyzkuucRHQcFHN
Pi+FI3BPVMGa1dxEwxPB4byYzd3AWl7c0voxmt57EJtxOhi8ZhQNW38rCEZLzTNA1Cw4xiEzfJmI
h62kCBjl6fJz7gS5WPy1X79SDPJCFEC4zvQODR05eHu1z+M9EtwziJH0Js6bDAAYGk17q0uFH5TL
J1qO8f/suLgGIftiImqP1Gx6Rbze/4FHRhygg4HJ97QyAFbsj8M4ulnudlSmcz84KAcR61OeTOpR
yF30iJsZj0DClKnXRBuQM+gZYj17h+lANU+aanQLu8SbfRW5FiSAlsDYW8ses313mh76bHR5MqWv
qt/6xi/LThY72mjgog2ul6vcI80Gte+79Ywj5uLsSnNXCyb40HNVT8dSB1i6fn6iX7q5piPnW7Ak
ttmC+YQA85Ehab5FzaDL1wFg5sam83T7Mt8tK3aBzlx0lOR/yiZYMwAAQsFJWMBxPmH6rfHHkd+w
8m3BDPmFrDfJ7/SOQtAm4q9ZzbqXJA0SB+kfHjLKPwZOsI8yFltSK1zezerLsm/jl4XBpZQJ9db1
FD5WtXILDbppuw/kEVp9HWtQi+6Fz0oHEQJMp8jE4zNDObN59DLAge12ZAM/VSTXvrb+ce0udKtS
DCWMVEaYFjzXQVxwaaDdb2F7yiSYqH3AsenHBHuuiOFoBGWpp9TLb3CA5+8LK/ttWUrpX4cYCWWQ
K962NKrlJZCwwHkXg4g6PJuAWFIRZq5PY+o5DUjTG9DjHgMKDgKtzA94rHSUYsEeoGLu4u81EQEC
g+cJw6oiuW2Z7AMMNTTNuyAsuL5/rNNF/KlKAFSj0mvKvZte0Ik+y3dSG9Nrp4O5rCerLCjt57AQ
PflC7ExkyK7IQDORoDQYtB9r6tSA7AlRVsSjrUI5IOZZ94+mm8+k9k5I2GVKkSB+7dOXh80Hy4O+
G0vPY8gKwFwYL5BAXBsvh/eRDD1ds1V+APoOmrLmdkSXWsbhP+orr8/StvzsDlF2Bgcbd2Sp4JzP
sLQ+a56DQ1IOIoPysWwbQZxv5/FW0Ef5dAFsAebWFQnn+UZp0ZN5MTegzBtkw4ecMGVOd5OAxeO1
k80fs/xMs6fhqFbmeohyZzTFyUNtMfpQCFLwrvMgs/fkZrQTi+Pw+NlDPq+rt8uB+lxfX25LDmR9
XyWGnTjL5cCbQbo74vJxRV88ZzuTSC8iVZgOvY+erB3LHTGMyC0osWaWHwOgC+zHDb2mBV0bNVab
3dtYvo1bsamf+FGSN0mnxFkAi+3WXf0xqAqzEaHsToAzn2RaLgCi+RA2Qo0q8ApDzpXq0497KOnd
cHQJBhyeimtd6RyfRavtsNTdFCnWMvZvI2FCAZNWG25fY30FZWvNxuQ3FsrtItTsAbcJNkHyRqc6
ylC2zmq29rC6Sq150I6NArtQz3kb6lDRglFCMSxt6FrW1FqE2ZCYJu3fOqEb6xBIoJeFro/7EpqX
lqIfgSFaepDNDa1lcUARXlYJU7XGxUtIwI47cjOVhciTePkkYE3nkO1ZfaHTRfnN+dLVLnVjOoAr
7reAaiW8x2PL16lkkAq0EEDPMpO5V3x9PlpbdmOJRU0kotLILoxQ0o5TlnI8f5sexGl/IMqPtHhf
txpnCohkTj2tn9VbLowocPsnQ1G00yRDQ8HY/IS9icF2nMyoD+6VgXKhAXPQ4B4pUgT/xypLshwz
twJGDtWunY+3JiDD6VY92Amc4+xhVvj7lM3cZ+H6i4BTYvxT7UDHf3CBai9uOp+1bR1TC1atdTwN
pY2Zd6eBerG6P76p6fd3Cc80sd3R/CxCOLEMTJ74YeQ7vQpEA4OcOiYkgVjmxkeSau3jjrffIbSF
z75iI8Oiohz8gu2WFuHFJxZ5tt6Hwr2xPs2+NWQNo6Dn+LJccTvTBLjj4tWCeOaPIW8utdLTpFYp
/4pVulz38OSwb3tFp5pePJIxXEX/D8Jxcz40mDtZ8kyuHY4ZQTGB+yLPoSq2NATTFh0xqVscK9iR
qjatjFKZh42fy6Q1WL/++GLNwILCD9YdPprIGuF3MxrvDcn5/TyT5jXWE2vjkzZ4k1onKe7XYL0j
PbbWwqyqx1QvVroYMFf/vcpht8p+LqOKQwwZa/9UrnfzoxKvB06M04eb9+wT9rzOcnAFWm8OvcaT
PfKyWrwtZf5EEpjkqyu/rwQ5A5NKAQFmqQ+OrDn+A5CUECHYY/Nc7uSstNXuUzcJi374WJA3yu+u
siQ5aNgkOBPXanTn2wB3aJyKgVCeA00z7K09jIluOwN2JIMvgFIxP1Wx94a4nvCDnAFB0XBRoKDp
HcrwQUiflOEPwv59rLceIFQi6Arc5eugK3Oxh0+8UhlYFZ2eiAf4EpfjKBj9OBfMFL9pndh2r26r
9k9Myorj3PUZqsemn0jzO8YN2Mo4XuhxrYXRSKpKI1BTD7J1QPjfTWmps5fe2JW193PtUqssijtV
5SlRSAg7NIdXI88mNznbsNi16EPBFqIANwKQt+dhNjS98E6RrnQfeNHoxdu08zpOCy8UM3FngWgG
2IIuFrKQiozQMsr/F3pHzW8wHb6yTN6mj4TeqXziYwtg++WNMx9d5jGpEgHWeUnqaVvmK3wtVjU1
dvh5RswZh3H0bhf3j26pQtkcmUv1yk+DCwOGQYC4/Mm9kuAhQkgBms4mix3OmL/LeTNdL282qPR2
vSAtiAiR5Ei9ZLiycZnw1NAaznR6z3IaBH+9/jtEVXw33V9oVHAEErMpXITulcNIP6RM+oVwxJ+j
D6deztqD/khx6UXcF8Fqz+ERKuPrmv9XJ327GYiprbUPxo6Ga/8t5/L4dScYc13DQ03IlbzukTH+
XSZ+7zH4z8q69h9NdjGOa7JZ+cizOovIMAy6/KT3MP/urPISLztbHOMG9+bUKiLk3sGCAOhYEdUn
ZSyxeDJzmAceMrFnothAJoES0jQUitPEpRaPsRhZmkvO4K85jfb65XQXUA+EgOV1NLyadqPm2WDm
pIcA1VMgw0bZrnyO0ClRDoz5VQR/j0ynsxVdmuNIFUXl+CyC6OCkIGkdVF1xFwCRdxAHFduKvvRu
pOLGYhti49UmO/RDPXonHJYqdkLhWfO2Oi26Vc1zn6mO0lRH2LNmiM83lO9sBSiqvQx5bDfcjZZD
HGuOcoES9q6+q4IcJbH4x4EHS8Uv6P28b7b2qsI4TVsSOeyzW/BTfUt1Z0koSSz3aFDaOjCi+l7W
4J/txrY0mj6eyhiUFwJfB7dDAnQXtAVAq2RCdR1f5ZH0TMog8VWIrhVOBqpTzK6hIEHYuoZdF9iB
QDA2ZY4aZCNu9vy4xuR1oxvZfP2lGK0vlTfC+NseqfjSg2/uHOIjiehSUlkbzQiW89D/rXJ8T/mn
hx48MCxqzD41weTndBV0k6YnAJxk5puzEZRZJrZVvMeSwM+xdM3KrYtkvFj+YjUQGnvnITQq1c2Y
g+yzupOxT9NTEMfcf2gKCQN6CoIYe3171TiMFTBer846a+FWCZM5c2ALi0WatzCjY/J88lzfhUG8
UO77G1+OY1G4B5qJ3eD+XNctD2CfJnYbu/nfrVwKLXuEd4IVO/hwhFoiTA00K0EoTu8Vt6QvywJC
AoA6fhuPZ+qMAuYIwh8BiFgq2XVsYA4IX7Ps4hUXtWrkz98Dl62xybQBjdCLTG/mn4SuZeOIKJC8
dDxJGn4PDsv2gwLETzzcUBt6Zwd9QAtDfM97dYaSyRltURrcS5jzt3KkkXYCnLKI7TSGJE+EaX3i
Xz5zGYDFRGd4GceRmTD3fcgowu77zwTqawr2H2/8EOnHYV4n1wKne9iz1aIFa84fdxGydO4wdLDw
BiLnr0pz5zWAGit546ovHid1zR+jdadvaLj4tvAvCq8JNhVjE5bdQQPJcsD84qAoSm7TVniS54R0
fyQjND+oyGVHsIt4+hxri/ciiuot5/Cig6+krXy+vvPvqqjxxJLVvk9H9eYX4yenja4pi0MZ84JK
MY3NmsB4c5Fm3EyzNj218Eg7rK3gapqUGB0RmEoTNF1MPeRDZwn9S8q93pspWlr9Nv8yHwX9Q+ZQ
x3PRt7QaKYCK+mpEu4hjE43OWtESKEq7k7RwoDWm5FNeaFHplh+xHTNAVHRME20urSxA3PE74d04
9aGRKyPM6lL3kVZ0woVjrF/k8xQePKYSuINOfxO+SWVkEXgbmxwyZtcJXrYIgITSuQk3DzAzOM34
DmWtTp2BPxnp6oSthnHG/+QTorBMvzdOEtb2A5BlJFNtr5kXobNFBrJl/ZoXDQHjrAOn0tQMDIwk
6dy2yU/9l8zz4e3EuuG6RhctR97C9UtHpUEVlttvjBpR+WQLPBjxreOvhWwtWOej2ArpDiSHe1rE
gQR132KFU70Rm0prUYVqs4AMiTMTTjaWD79N/ZHSyKu6hJLIETvTBIi//SXUEha2Tum9K8mI0f7Q
PCcRNVq/tMYQc5bstXthHUxepU/YlBk24o+jq6xXYKNZ7Q5i3U5fyJhiWyjeOdAmoa2nObzlopc9
ZOvHtvJyuUhzZs+9VSfM+hvSgF47hKpnOzkSIjeVJo57uAwnAJB4qaZkajmobvNs/5hznsf8kndI
dR84uoI3PqiKlUCLBGXv6JmzpfWogqcn3itwjqfQgKSP7pAmBEIUfpWB16qdQ8WryTirZHWzWL38
i3V54pgUGJEnG6eDZm8cCR3HcDgwj6YeKI3NZntKktjJzG84FkgJrxJ8AqHGrf4hbOIvL7m5793w
uiIapAfmjkaVktZmNduKF0nOH186j5l6rOCsfL7rx/0FXEgLEY69Ir6p1bhRDwuOkFkaHQk4g+Kr
GmMrnXZ1GPgM9lL+z33jGzNUG4EJoq5ORYB/pe8R/XNwfHItpTCEn0mzkLuTJGXYoAPN1UUmc7/9
KwGiEBKI6BK1qUp7mfgUmQ/yAYP1V4kE9X93N1imiJRPLug2NXhUadzdWu8OoY92YJDbu1bq8WCW
P1A7KEyg7kUKKBOu9Pwl46GYUoIunQ6W2sbjWjRLYtypQyxOlrg4lTl9zPsVoVskQ3/XA3H+Vh5N
mZLOyDfJFb6N1Qrwl90cWKcOWBxCcTGPxw1jUOGiyJRUdOnKpiZDiZNVZC+3OYlLX+H/ntGvJQRL
qCxTEFmgbfPRjscus18RzYwxQycVXLAXB3j/2gu1aAXNbCpy+jjG8S1wPPWRq602vMUQ8T6u7QGG
93lzqhRdhEkXPbNW5PQH9mpo+qLUskzPhC9905kEGLKxMNMJqzYOprkwjU1uFXr42uMGSm6ROgc1
bHKa8KiYPSznnAQKcl7nJ6xj6ZuObziHFzN5PDEUwo+1JioMY197iKz8FfGRPH18slckSOQizInx
LDNRhM9nMtKF5QmfEOCKAQupv9c35bexROwFOrb9iWWyyEjmqmNqR26XEcRmPLargiCKgzTFEKBv
BaskwAImnfwdJDJZXYxa9frCQUG2U//JI3XbqdiFKy1H3wPvCLOuGlmZfccV/8w7rgaF/UEehtfZ
10mbttqWHDdHFEnUWVp7kERKIlgtfIRPlkggR8kvmDJ3QLAX2ykexFW7ZKlYYcaNcorecv/fRKzS
a3ZWhWfMRDxfeWFJ/UaVPyxGfMPzrF2O+mhqsNIDvgq81NBPnTSjuxIpmcs9fXIIFI5xs3LHYGlk
D3Ex4/n6eXDdvP4HaY97G0rwgUPs3lLujh334wD7S9+nSjYQa7PWePbLHK7T3L1NTm/BfNQ73jOU
nrWviO+w40sb0eXdeoB6Nf8DiolGH7BUQAHQO9kaJG6fAOslGTfSOXbvuMHv475Ixt2NjRuGTD3J
azd6qwcBNe28sS2xQrRWQ3mI4T2S+NyqVcGBeTNMZSo9UP8Kg7c36YuPHESeLcXDEJ/JEwJ/L9Ws
O3IdeWSAwFVoFgMCLa9XIQHiG2g30EzTDTlhexyYQj3KEoUPeOKwLA3ZJxO1nPF8d8aXuxDIXKZ4
dl6RUl/+n1I+4QBRIlIKwjkhefapHc/Na/t/Q5lSlZjLxVm7SMwqJtiCceWIi+3hCaU6AtK3wM4y
VKNdAPlPrkQtp/AF9GUhBDnrECI0wPHWyK90H8rklq63/TFWcxuwws+85pv6QKizOk0QpjbkxGuA
O0KiKaV95bgXngbQ10ScnKch7eKTEGK1af2wO+c/IvXHV0XIQ3RYLtRDHiY1PsoEZ5Obyfhk1QIG
BnT3ZgKrfmhRxUPDo7cIbXZpCiwKSdbDviTr15TNIN8PWN2I3xHCUXIOXZhitiiGtugz5CJ4qhie
yJ1i2qhbD6FvQpOFJANWewLRqIq3VBeEdNAzYs1JMkWvxqY8dlXVyurqcuHYwwJe8NR3XJ8MWIzK
fbSOJ3wQnhXydmfn/vKF9Iw06PodPD/FB0dGdnvmFRvyfdbAahQ80xBVytma+iTpKdSd3c1cho0z
HMSBvqDS34L9Yt6chMkNRwF4r9W43t7ewjhz0eGZQ7f4Z4kyKvNAjJlD3llpQW1JscsagdHpHpRc
T9ISmcudM15NMa1dWl9Vi52IcH1bxO8962balfon6bvBXfvg4TlotK6Tlb9k5yq4GYBJwsVq5RBX
UA8zt6CRyui5xmk2ZTA3l9BXQ+JIJff71LvYCc8eskd8t9u7JxupNGdqEWUnaFmbKWTO8KnQqlAC
aaymZF/SapOeP/ZMEKTDYIU9oHDhIuWcF0QIxe4CmqfWpPOWXwILLfkLgEzK/dbPwpwUUfJXRwcV
RRyUYqaUWVdZHBGADlN36vnYTXWHmoxh5t9aacAq+1oBtksGaUxp8IyasoVSmn3pIUrybPd4WJk0
FbtUuXAt4j/Iwq/etTT52T3CdyGJkfrO6hU33YPrILB5cMxC5R58QflO0KZovvMRA/j3lQpf3Clx
yqFN/mkZvQ1oCIuC4zO5bwFgU+6tasVOOFZ3nf17Rr9/CuthnEp2d9l4HsPE7CemMD+zWXDapoiE
W1bSVFgdJlUUWwVnNPof6Hvqbka6m7v+WMpOOQuhgTl4ujAIqGm/jLCYPPZ2iJzzxvR81c49shwm
Bc9ISpMQUQ4sQwnKGQdOv0CKp4YXByG+an4ZU3JZkxDPSDlQu7ZjJgRRpyvhqDQnKLY6gv+b0fFv
bscGqGzsY4JuO0wmotjozrVI7hAIA2nLCygP34eP4lQmQU/ZOX026OCTHPPW9Dao/vNMlnbt2EeJ
TK1p2pvHhHbLKy4R0ZF87pU/rDwMwezBHQhvrLCQGGJF68Y1wGBiQvsvE1pjqx32Wrs7/yt3h14A
tf5SLZQkKcxMFkzGo7GP4yC066GuR6CgDzq4Elg8C+ljOHzQjjP3zlyodabytZwnAWlLZaEj8u8m
zOs8rbXFCR7moXr3tvPu5xKXVzm8/Q8I3U40LBVZERrqU96kLhG1ipyLzpBAtJ4vDEy6yrm+3XD7
nzF+l72r+P5xZSnEM/USfCaGI4isHS+FHHDntPri3ncWz764z+o7y9tFdcBJEUzI39FwSHVwfrFW
b3DggVG4hyqQUaXHq45mirNb1T7u0FhGOv1B+UQI2v8C9c9xZzKU3iuGk94VaxDDoKN/k8imNdQw
5KyRcnrEyTY2bopdpugwHjNpCEzgPG1rCMKVFqQgcZcR9du3jP/Eqoll4sIH5yDA1UDqEc5QDKRJ
5VPo2yw28OibRrO0pGJNggw8a20mylrtg7R5s5DU2QO9GXUlfKxCKOa51UFqRgwUoNy8F9VIMy9l
z1sj8/lYX3PVEm7hC7QbwJkWolnM8LHm7UfDgloMoreb9ih4dTaolXhWNSsY5dyOKaO1SDLK+snN
q4hGvH5s515DF+VduhNOC6l9m5N6SYFWwWRYGlRqZvxVBtlTkqz9+qJsiGU770PeBdBIUbb8Rr4x
r9BHZ49hJ+fOnJ3mR42e3lUUCJLVWKtfZEF/nTjr7onwbMC8fbCmFQf693X6yTfoLhbwV57llXME
JkaZ9Yz1JaAHksN2YANg0sFhZeYqigvvXE05ejFKinHYpSLtPTiZN7ZG7eflOfx+Gt1E1XIxmVOa
lWi4J/P6DBG/XCCkcJ3Khp5k1nqIK8Ah2qooqQEHY5z1g4sSUdzvqxH3ZE3qb0o2gqMwSip8i07g
N4v9cYci/j9GlhUOJKuYkzxojxXxn9vLxtu6CzY7lktv6XMJouElf+1m8xoXOck1yKZaEjaRdhFg
NzLqcwQOQY5EmrQtW89l/la0735q5f/V+nNqPx9DvPEIriFQOLH5xyCSWAgvJgPuPQP9ZdlWCD2Z
1rTaNa758A+IUDTeAAelQD7TtQVRRf6b/59Va6QwgIR2vzgYkgJaz/HeE6ACjqZpwKeTwECFb9G2
oqoGADNdQ742zHH1Gbto/8pBiqfSBrepV1BwXzJ2CEwfs7jcyBvVvY6vIdE5WQzZ55FtyiZLQn9A
8BStg1s9bX/s23EEPm0RBcIMtDAxtuI73T+pIh64v0ovpFbBdUOGzk0cmU/tNwCGVNipts7WTOmn
bqQQSi/6l1C1j2MB71e2/J0d8Db6W6XZo1OOmrKN3HNWeZS4MoAoU6toHTNOY8A1angi+t8dNaPV
giGkPu7dfXwf0F9YYqmY+gVNm65vamVj55ptapLNf4EgC/Nt1cEUbi7D01+/sQhRUkgduht4rdRR
7bqGCHwX+kBSBfIvfFht/PKKtgs+9ufi/O4EVAmPE8EVAFFgsBmMFL6Fjk1ooSeXqEJnu/E029I0
vy3BQ+IpWZWrPOpFyo+ypVIGUOA42YF05UP9pR3EbLAcnnHvuDTWmTXbMmYYT0sxaiz6WAu+hvNt
c0RyZ2oyqrYNmAn5X2K86xKFkHrvmdJN74Fn1+dT8COBPZpMZsY8HN6G6M0OQj+uk1hAM7LaBHat
zwUtJn9kxA72EAK9yF0Y1SKbYC+UmltAenvOWHyKsNi6x6ixQAVhoH0l3h51COVvDUtFm/y0IW+1
4aWno3T/LbaZAsAUE6CwUosp1nPLSiaF2hfyYGoTgOehBaUvt1t2TGUUzbsG29PbAKmQKHpwkH80
nyYojHlv/RMfa6tKm78EJTfMJsxQSc9MjCzxvn3trmwQXxHTaUQcJPFOSV18J2K2uKG5op7ypFz1
CJutX6BNnT6XRGvtpsPkP0atW9ypoQl2HzTXvQF03X2gkW/Lejggm9jWkXEUFlw4ik8rXXXU1een
Un2h2wAwHHX/XWSuYJB+/8Ml23kZGIJZRe8P38j5HZm5DQa26s8v1ypv5Rn+WgnJS6vJO3M2efYh
QjP1J1ztjUDn86XwfT9CNj5jyF/hG6/3AnxRZxAF6D5GLMMtyoyZYeGfniB4JT96xMgb2wpTyDbU
5CuPQp2IdcEG23T96lOnxcFkFxj1OJ/z+itup/j6Muq8D+1GKg8NWpE4ef8OmIR0M2kZI3JAmqhY
Cuvj94XkJgcoAZVpt+TcrMIn2dErzekLFnOkCCs3moj1M6VnLLrgQbY9X3Z1yvIxJ2S8uCdSa55d
tFMkxjPVD+RAZDzXVWW1DrkrwNRaJvPW0QRgxTtEil/HHnG+pcaIL6xLA5rTuB4v0BbwEuDk6Sns
zTXU2Fk28yC/zwPBB3RZAcWZNNGUmXcZjjJPsN7KIXsuMysS91kyJriqRYGZmerFHBHuruBCVh7C
MLAQdjyI73tpkWb3ORXm9cNAnitPDsEzX/6E1A0gTjP9P8xwvwIlu00s0+p4Bq5WZ4bmS7e9GCF4
BeMka15J/LwaIyQLB6AiaD8TrkWU42p7rn7ljuiR7L1BHz6WdT1dCO7YPVb2ZTo4OwylcIaRI5Ra
VdM0NmnhZsIMVCyKjzK3Oil38nY48KZeV+YTAII+OQ5ikBn/6reA56mhHBc605NdCvcrP4hDbRlQ
RXUW0YtNJndcJNR9sSK9lw4MhZNhdJi7DKSLun4qbY2jnu11rqkZdhNA7h5u5G55cFFQmU7B/r7l
tm9riBd5aBPTf1gnkUhXT6CyHiIqWNr5FRIujB++LMCrJXUlHpd4P6DSu2KsS61uuIk6Sy2ekRaQ
ObpMZMdvwjBAbS63Xn84MIXpI1y9jBGZJux4jW64LF3a2oZfwzsbALHRucBd1N/yeaUBMASfgGAY
fL55Ki6Ejt9ZTZzdh6U6/0QN2nE4Efmq4P1R8lCP9t1MtHiXrNOtWjbPEXJbEenlgiQ0I61phpzm
1rOXzzwGhzu3y54V2XDB9f51dujM3H/pWLD2O9YNa/AR0MZHAq7Hkbq3lX4+jbamYG/7FoKzhELL
1Q90g31nKZLYSYb2lkAW0M10x9OyA/iG3MNdLlpApEaoNtTxWxWYAB45l3g5KHv28rdsYUn3ADq8
tmE53Ki8NuIsqnwo1m46kyR6e8UbVbfbNLTMkMj59MLOzWBRMbWW0R+9QpQjyztdrx2SEFo0wjHk
NQWS1Y+6aXN7rg8xA7H/8zJ0C8r5MAqsw/ZFdpJw0hYJvncTUHt0hFPqnleJkg5IuBWez5QnGcor
5xOuSj9Mo1w4GZ3JcUOuWZNQKh9utxNMqU3oVH7im+MMbbLjCOM0JhaA/qH/hICFBi1E6DSxoSmG
qJS+OdzOPMqamax0G9x9ys2lE93aZCBkuL1sXs8FdbH+KVFfkbiEdTGnf5vSGanFhZ9qYvpZuUT6
fF6oWlLln5/smlDI6NeVsJcNZdtwbT6rJlhJR/8ZgCNozUwWKcOdaHAUl6RD7W4w/sW9dRLY/AOn
fN3nD0B+K7CMZP7E4vjX5b5kdv+aFGqW8WnHhBwB32VdT/8GItSum8cFkyTuUbZ5EM4d90t87ipd
Rlyspo9IKndJQG7uHrKjoQ5pZT2YjsOaNSCRmK7AwsSXV/TXaNwHlaRQyed7BlBkv1E2Frh2kDyL
l1eqPaXYLThP98daZpWRuJ/D5v3uyeG/p3W3T5+0CJPedJP4O1v4o+lU7kWENqlhfuAdIN02LSg0
9ConH2Q2LRPflweOnuh+ApBg+SG02QxncLjDMOg2gzPRdjoI5eWwX4ca9ckYsInHrH/5fL1iCEJM
uWXlqMLh9V33S+hjJn6jTf1jDv3Uqewth6m5cOHuMBZ0hTC0wEmRliCsm7S6TW+dvIsQ/XyS6978
YfIDFEbGQGeEK/mdVILRH3qshyDX7IBQLVTs3hpEScODuRBL2w/4naPAPBgoIDPGUxSrxYaZeXZR
qx8pE4d7MLBFxIwFtff4VdhV+89pZ483VGvDm/KluQDi0eyMx+TQhPKVrDUEG1mFo9MOYsMt3U/8
CdqndjZBU+PPkbT6FX2jSwft7tv9WyqdHeJo8PJFYoubsJ/DkYXwKN2/U+CrXkgZEE515ZtS0CDD
SRi9hkKqMD/TzpMgRd+vxXjGEmn48fGXQBrX4hw8C4w6bPL3Cp6mo++zLcrU/3kACpDSNeNWfb5L
rF8Zv8nBIgQjrBdeT9qEC/JiecoKwHo/45j0rWips6lPcMbsvBZ5nr6nyNWPR0IFhzqQi21yYYWC
2B6XBvMB2Hq4KCP1fkS3uqu0T6fPnXeUP0tMUG6KIdnkroj3iF6auS/6VWI7mAN6QqqXgE/1rHJw
HES3qhq1ODTAkFR1Jq5FVKW6mvFAA6KRBN3ojKybIv7F+XgCZYdwRAOoOCV7grbQNayxvl4DD3tk
paFrZ9TTzV+H1DJMNZMGDhFwOC1LsU9S55c0d8MIRJXrTXR3Gqs1v6UTDg7E6W3bHZzbhoqQCkBG
FuF9Qk8VivXRuf61AlkUBHZw/uheRpmpXriy2NxwPjs4p6CaVumM/iJpZaQX2ZQjp7jTzqXZk95J
RQ13JHeVl3rH/hyfrfJbHWzycKN1mOwUFOLqE0Fi889D8DBhoBNw/G7dSjmKRjw0CjeC5GIGMh8y
ZuSfRmEgtsI5TsJd/iqh7l6NnU6uUVs7IlIPTVxP5TZ+oOVJmfz0bEV53zBaLFW3IUUQXzR83I3P
kYUi0onzNFZavUvSlD0v/mmbyDnkjdVggbLA44cILAgHc3+WCvtKIQv8IDpMDJR/ex+LMYdiWFmm
IEzPCyJXUM3HjynBS0X8kby23pyBNjc7NeR/CRTBBid4XFYBthCOU0q1NJA2Q0WiqYu0z3NL5KFd
IbPESxn2R7zLzdEI7zUmDrpHSoSnF6wVovSt6bIEXdagLSM3u6RMPx5TnMYB9RhlJrq/qiQaNl9/
u0XhriHPXAIjp0MxjaGNsUCatIUf7t1sIre4RrFK1QbvnApbltt1Cwru04xtlcL0xRJxZuv3wcGN
bez/M8TiAzo6YvyM1JP63/1avGMfupb+pH3iUczAC66mP741Zk3NDSKLCS3g7uubo6RgG40R2fVA
149nlFUf1/n83GTUf06rhIQgtNA2xrSPSo3rY/OIdCjZOx0mCC6bv9IJmVGV50qHeZw0j2cvwR67
qzupIpBtdg+YPv5b+lCZO6E48kNaO6f0nYsPmh9j9pieq7fdxGfMFD2JY5Kqxu4TYworVglF1yjJ
/wgrcR5f6/a73RggDgsoY+c6Of0lDwMdTU0RriWpwmw9lcdSGw3GZWRCA+jIJNxlhkyRoM/ewFGq
CO/dNdTh+G9Ac0kCLbwCpGciZIFwTbnNVOY53pLeaeVBCEi3q06bgl2bokn/CInfKXSrUkMFMEhT
qXTqWqxo/f3Ji8fMIBJExFf3Mdcvpjt52tutvWcYEEQa2uSRGI95/Xvz1IT+VLgVusyguLhIMizp
kaQFlok6MRZ4OWRIzphDuZFYDZmBHOgNmd14t/g2JZ93GevNnR/sH6/BC00vyie1qFQeVwlgj9lY
GfkM8dfftM23SfQnKB0NjvvLhQL7hOTH4Fr27t3ts8jKW0+TU5gTIwRQtHzDH1dv/L0WQxpG34Jw
jSw+nOmkf2cJHBCW17sRGBCadfRhtBNJ95nNs1OWGs/VXN5xMy3i0MBpgyx67UV0J5uAx9XoFeE5
X0d9BYHvOSON8d8MQLJxsCxHeAh7zdyEcKrl5NIIs4lBAAPgVFQugjYXKVu9IHuwrAInsAinzyw/
D1J2HSwHYI1ZvRf/a8C2C76zQp+aHxhobMmkviiX23i6/GW9SBtl5fLVs3FgYe7a+UhgZyHcPhEI
6S4CzOUb3wrqiYbuD97cVBP1G2prG/rZlsInIPwoXGTeK+DqlpU7Ko/7mN87DEPmMWQAEVhh02wu
dPGi+8Ynp2AxzCAgm8sw5S3apY00B6n2IbBq9xaxoTcwE6LSaoycXT8zfjCzZn/0xMJ234vnmEYd
R8ytsPmIQQjG6sEs2sfxl5sXBDU3sUJ0+hKezajMoedFQN20TIXtH53MBZy/0FbvgRQ8gbU+2ecH
yUHE5nMhG8XEG7KoGWSm4ucTEeWlkQ4cCtGKHsvGiTq3WiuSxlBRoYmxmrtcEM37q7mDu17X4dXO
BBnnizMZ9n9EzKubgW7i5gUkFKTyuMO26GCeB44K9pgBhFUAJrxNZ1q41vQi9gRhDzajoXP1XtI9
iLSGjduJN+qOt8KOFxwjlljh0ArDhER/fB0gLYweo3vP3gJp0O6QD4Hw69HMUGR7qtrbHosfV2lo
286clXFBXIFNtC3HLfon/+TzJbNqdFrwCt7SJT+x1bf/Z/3Sor9uMa6bb8WbtVTVBPAVwjhG6msF
mZJYS6XCuSXuviugSZ/W/Tn3cxn3G2oWjfymWvjPYLtqvqToYpAFjWt8bu61IZYueT9qaJqPdmeI
Wgkioomh3skH9BwOQIM2QwhExjAsljUJYTFzxam4yA4xPIBbUBlV4XSuez4x1W481aCkLWLJr0+n
Aq7oUoCujHbSTyyJPZAizrToIjcKP8EuPcjlRxP4I7awQPZwdohwIt97reA+aBEvQYmgWZOcVdAj
KVkCS9VAyHUr2VoDbxtlX7j3HkDF0cfINtRGjWyQlhxbXmLEe54mRawRh5U9/NKjgFnu+t4jTkE9
DsmzK5nLRWA2IOPaKxXZGCOTkM6XD40JsoH/Fyd4NskR9Zpe1R2nPUM6gn5hS7wzgJ7aIGNJ5XPj
MNjRcKlxUVf75C+fgOpCtYV4ZMaxFe3s+FMROyktf1KMyZvwpbBFmZF2/Si2hU1Fmc43YGpOOK7u
nX3LptXw0Vr4FiZRUQzcnLI+dqx8H+8GsrVoW35o3+qd6emKGPJtCbsJACXDehCNTtDznL6ylBqT
ofdJHwNCzRc99qjmWt0SnJ3rC5V3zZ9ezm044F0Z0blf/ySW4e5rNGd3v10rPvKaRM1IT/g9i3KH
+LGp8dM4sbSeYpLcQwNgZD7yHOfIuyOru0BAieqhcMKuv6eZdjrYk5u+6d4Mobv4OTa5BhOdWqPT
DCjtFJcsnDNEHCSWJ2834lMuRzEIdroQdURBarw2cQpy1ujVIg9M76P+VQZ0847OgCqN5op9E03r
hszLUiwZXR2M0MNf8d9lyGz8yF7xl9RoOccnl7BLfkxL3CWiuXxYAEtxec/Oe0gZSPlPvcc4u4de
MHzXnBhDSXXoamZjzZ97pkR9XVvEokcgNqW7uX2zwM83pb4bO7rofpXJkzALJgs4RcEUFdgWEZ4V
/3HCQDIsMHifu94QojF/SB8voq1XNT0vbfpt6cnORpT3yETlmV17JDuFgU5Ld2Mw5QQ0R28iW1XJ
C0px4b7TQJTGowbsbS60BmVSmyKzMgIIp3W9hGxXspPQIad/cDdMRcvMA+DF4UWntbDQDhh2rpgK
MRBrciGufdPcPNo+a74YesiOLKYsdxMjYASB8p8aaeT893s7lXNbdod8+FW1sJ2qdhyYNy3p3CfC
2f1YYVZ4K9hByqS0MiDRmjoIFCwV1388ZFNsOep2/FXBNNgib/8fl5lkZG0itYozyNRiZS76EcKK
6FQecZy5MB9jM4+FtLvtJPCgzfb8ZnxsMOGAm93gp8Zs4Cy9XA9TcSW+BX4QrfhBY9gBgsY/1Gmt
AR0ePEdDmue1+3THaD8sdz1QvxZcv5JVQLKXRYBWJaJTF7MEnxsxfAl034+B2IlZJK4QIBPZbHm7
ZVmFmRT6Lj90Vh369lJSqMpIVqHegbz/IebgkzPzWYN/TRyIkmTO5y7aSRH5Oh0sGnzjEHPhL95J
6TkdD3GVExxm94vuoYlqy4eufsX1zZf++g5F5BASDdrCQKJ2H6GSg2sOKrgVgHnzvZW6+vn3/Br+
NjFFI2kbnNgTlkyx6+H4b87mw6e/CUo/bduBKA66Ev/N0k9AfF9rqNS8lw5VjzGSRSuaPilDrZec
0gjKtpXj+z8oBgPWCGm+c042rxdlk00Ur3kN0+xxRiyJAq1lnz2II+jioocVH2wOYFtLi+DYKRuj
yF3KA+gMcOlw8eBYXVv70xBmtVhi5h0T877xvgnJl213m/dbyY4U8agCwVQITC7bQ/ubAWrLJOsq
mn3+NMpekrGtJbyeqKmQsyfU+S/afTiL9MWHMZXvL2psvlxsMcMVeOq1CP5M0QyVd2wrcPj7Bdv0
dnhTvqKBH1ystLtrHIlhXsqkIRgB0Ly/b/X145MTqZeJ9566Co/0+wjqVobfIyRwZiTkVSKN6FOJ
cg0hg10QjigpZ3Ny+xPGB4E38LWY068pxu0DtfQ1QbG0MYMIGFXBCvYOE2tQ94zlQK8U1sC38iVL
1P6ZF04vFJjHQjJ1E4QXWlQyh6pN8Qs8eqD+9NrolumqlsvaHRI4a7r7qDdNoiyr/L+NmB9zbVcP
Q4+7g7Fn25yJnfbo7peGCG+VY3g+BwwND7FdrfwL22TCiKVEN/PenPoI2ixH8brjvnR3EP/NKj2/
Az517yiW+dXxHt5nIlYf4GBVlnB1tpWWW7wXEw3ac8ZWIFh6e4znwwxMxrlfAoMbv32Wwwtlcg+g
ByT4uEYCDCMPyxjVBtrIfmAPhhO+Zrbeiu9OpJeq1S/Azc9llyCvzcgxRKvaOabPCQkNnt/K5Fgc
+EmKyHX7GPCEUA2tVYst/u0mNNbtTsdS/WkZAUEw8OC8ivR8FeNFvFt/P1W8xSZFuBEvwawCqAt3
q/anmKZjHJje93xSw0bZve2t7H3bZIuW3Yxvocm/9Ug8to6DtizWF0NN1lW/X/b0cLgkBETnaERq
F6fRhQgkfWyAzuumFc0RrCYXSmgNBzdDRpdulRfBKlEj6IBM22+dXMMIDskjl4wrYVHtjoZx2KEs
iqrIPPDrgcdSlNFLxpyJzlUgX3nD5597mg5u5hDf8wJy0s9p1BlP0shRg0Q27U9Hpd9fDa9Y9owL
7Bolijx4sjwMyOLhv2I7sftT6aa/2+ws9fXXca+C8wQUW2g25vgrqDAKbxfdu0fKhOIRPM/6wLQX
zyR0rmJtLprQYGSMo+VuIawBMCyt9HiUfX+Biktfj2k6dZKXLK1zgS2x5n4nYwwDm6LGbig1kWNy
W2FPT/iAlIl19daZMbun+5Cn6HGjEEFvqVSjaxVLUwa8a5boN+ZAGYb7KbmlhU7DZ6Lsm/ewWmAc
2LKLR3gE79Yk8hQ5/VOFB/uPbIxmMCLJLEzHecLDM8GwOTKt3tCIU4xi6UqCmo1B5N60wHZRv2M1
8HP01aanK0hOSxjw05GDDYIgez+rnNlykf0BhLpPYtR+9hiWL1bQvFQJKIWQXOGL7lPizG69XWl6
ovHCTErQQzKyVuHjH31H+flJL5mPq4FI3+gAu3QiH6vNQNDjXjFHJ2h5Zhza/Ub3Eml1ZKSmKds6
FYhfIGpzE5qnshh2jwR4pIm3aJzdfKcWNMA56vivouwiWEDWCo1mgFh4VPJjQ4RinQY6XEMOxhb0
t8ygz1QUzp6DEcLSgPsTxb7LUg9M1wEeEe9Ghy0kwQyRy7PsA75kUc1qWZCwH3LVvXcUCP3/QS5H
hayTXKY99Jt9cLAAtUJ3xv78BWqctqy6zZJAoQiS4XptyKryQ2vFqcjdF+3viFK9gl9qdVlBGUWR
5SDddvuLhxsSrK5kX3CIBLCBxCKEO4W2WUPhTOqnBuy27A8uImGNITjFNDdU8sWOYCFDtJmBxa6Z
PoifPBebkbSuJSHDUdTpEhr6YJCxOAynX1cb3pi7X7VGfWX0tNmKDBEcTcPKC9539OKxZonoMJR8
AyrTPjMwLinlqs/yvVR4Bep4C8Kgz064Piih7/XKHk1nRmLzMO87QqlPPiMHMXMMoU8xctCWPoK1
Zrn6rF707eSP4Vs5YWu1uXSWvQYWcWlTvci2MAARv5+0g1b7ELCNpQNn32wQEapysZD8jDZEaMs/
gupQR1nXFmqon6la0AndldKTsr16YshlBoiY/mgdgW/WxzNyFswwFxSQBjdl6QfABgBhVlNove+C
/00FsWMsKAYdJbbcgNoBSKZUUDCvTYw2SpqCWVrMr0ML8eg+CkUxiXua2P2SpDYNnYCv71YD19lb
Gk+hukArvkL9AjGnUyhmaIkDGw3P3QHnnBiVM/SWOlLtccQImTzwJ8SvaU3rhUxKukEfonEug0M2
hoh/Q0ZftrSKqocU8nDb1GUmBL3FHZEVR1YSgpmjRpJ3SrWlS7mJ3jrEnObUVWkiAx2Y6Cc1PW/o
eZxjKOEcRXi0i/dOE7cUhGWj/ZP60XUZOX7FqV3I+/OyPSURhSmXKqbv7lV/F9RndPY8e9WJ4J0b
rl7CPJ/+NgkUxRTM0jxBaY6QMxANjyv7kyK1ywXkaUz/HTMLkVqntatuwxmRgAJdhhD0tFwU4jUc
y7MHJ86KUgr2+cLJLJTUFaP/ZwIbwfVMA1SnmPAz7RfQDcKsM243GB4SB70LhNgv5Qh8wAI+hVRT
Fso0IeeaWzuiaoxBMHzA9axiT3QIH/+hp+zPnzW+UffyAeBVNVsTKLgrAKx3OhZKpNmcbH9pR3tj
vefRcDKJ6sCwgLzYxkjahQUl9/g1zpKx2MSaXjCOB6ER8ptCZ1ZwZD4tsBRR37Es+j53dcPDVbMI
LJ+FtWmi4NyyAWQroudXwSORO7Pl5rQHTZz8E6Cspo8YxU2yfZjWm+GtT5wYwh2Lf070LMshvjHP
dJ8YqJrSpjaHsNsWW8G4Z92Crjqb5xAq61FaakiwnLi1OHyzyuIKQ02gvUxLea+0SNWWs7BNHmCk
yAZnaK/fxYL5VIKxWJKDs4R954rcFU3UdG9vhw6ikAsSY3G4oTKn7uZi4INB4XDjM5jmRFFGorpY
mYgOuTGMXtGpDDQYOUdSH4CDn6iqjs0xE2E0rYvWlmVURpGgPSqCCzuN6wVRcJXqzqt5eF9Vnska
dT3VfoQvuXSSSasaStI+LCrWTJZd4tRX2Rr+fus9NnE6Hib00H/iOBeRG/fKlG0iRdchEDsQvLus
V5XXuP+jQk/b4Baoj/3QLYT3e1c2v/wLkcyZoVxSDNIEwpkOiTfpzrBe75aHAlAWy7MepJOWmtKd
T2hF4qdB07XPMU0lofXnYsEqiluB6pg4DkkKv/Ou5BZxhzud7dQQfA4+SDyqXnVQR9fW4Aw1eJx4
yNjvOZTREzlJoeDgyqbKpyNXmmy9U2LO02DIG0HjALo8KOcXYS0joTNISxdUuvVQiy0zughoZ/Fo
EHXgseXOB2hwaAasg8Z9yBz5O4mT7CLtXvLNN0igeHKnZMqZ2aJts8SqQrTvxk1o0HW42g9fR4T4
p2ZR+hTcTNzD2xFBPw26H3jGVgdQr42bBlvckmasmKttjUukDoqDnnHb4mI3FewgzHx0kdQusUMB
69BnGXMW/lBw1fwd9w2VSqAWOYNHLTJgAnf9YvBYFIZhlNPcvjsbQUvxKLWlhC4CmjjdrVWgKX9k
DXpn0j4i2sBhotJb1MoI5t1qboQ/XB2aHkQ1Lz27vT6eoFmVouPVNcOSqLjfJQQGjiYAwBVNR0Sr
HWCVCOUs2qjTjYzps25hUj/qRBaLo+Ehlut+CS1lhDYM/iJulqjnzm9O65Ygp5hZE9K803CZqc6C
F59tlDJH/DZzuW6lglxbq7PD/+PQVp+QiBG02rFXh2woRjL53joL03rTgy7BwDcMNzeuLzTk+Xfv
xuNU0ItqFv/T+X0D3J62Qm5O/6+dKm8nUctT7J2iIkcCuMOKwLgKnLDnB4Kn+uGMRe9QIWB7X8Ce
wuMpAbYSRjhKOdVsJjOBd0YuMScMw2OAsbs9tu3RMswV8Ic0xQX8xYnvWizv3AuAfIFQAjkWOKkt
PaPfwQfRsaC4eSZReWMjZNav2FGLWzBGFztblvJFfZXD1hGjENeOQeT3AQuVZwrquQT02cTfy97p
4ACO08xKOLPkGbXdaCLsC/OygDktf7Qyjk+jgn+UFbpovjVFO+agrxLRauykp/blTG5pvpv3Pwus
Y23VODOUb7QBgFnIACKc3LfqtuzzoBqLM89zjJ5mHQTIsKLjlYVvlunj9mYzoJCG4Pl7xxnio2ra
f8yFul5EKgDA8I79iTMUPPEu/Yn86Xa1vOADN9HPEEWIcL5980qRmqeEaV5egSq6dtHj+vAASHIl
kRXUn/j0VQ4Xjr7KH4jNfI436bphWdDcqtooL3tVDbZL1v6cBSM3aiXjUXhNmcy6DrOFBkasdTKU
Mk1kaoU/Yka9q204BFBzUOH8yIde8hhwNxWTtz5GIsnqUXRn378lLA283o57Y3JYChNpCLfFR2VD
On1h6a4Z400DX0NIl0ZPjdKytTuG+EdI1Y3asHTtsjO3NbB58oId8z0jhOyblhwnYX9d8gOD5tv3
P50vdCxsNoySbOK7LMmTS2yWw1QHP69GVk7vl2iQ4ShumOdFn4pJTLz6DF1FcFR0RzefPd2iTmuE
5tH8RqkD5TUvTsslyyegVXr+GsVAvFE+Zf6tbjWz8aQocuzred8v+DsXVP/WMasXQiAsZ6vxzF8x
cAwe8trRNyUKYtnAkUHv5pqOaoM17/XE+Yp1Omn3CHzTtvUUn0CMuasejdkvpaqRf6oaVZ+qSM1Y
1eztwfW7hLGpvXFp0Lb9eYCJ+afQkUxJSNaWheD8NmQPTulRIlhaxHbDhWQyEMbORl/QSCo8K19N
sZXQx/VjAjYA8L3TEqXOubt3tdXW8oFVnc8jEpHCvj7pxV/YjuMT7AWG/UM3uLShm6ET4ZOb6emd
PfrYFj6FMmsgR5NKxnCZXj5wlEDarWHHyI8FrkQzfw4R42cSKR8Ly9Jr5PXyxjDtuqUM3C7nyHsS
cjmnipfTOL7mJL5oFoZPhDmxgPdgtGbFIC/3ly77NfOcT9LkkU74WSvc4xlz394J5dXLLGMtcyh9
sWKszq7KlmUeqePqZnHTDdfkpS3Y17AFA6ck4t7HJXm87S/l8wkG8UWSo9GwjE3ldDeLW2mcWsD2
89tUGpIGE9XT84HIdS2oJ5lxQZXDukl2/0HHA4mzjdOZiRHJtLkldXZp6mdSp/YneK36WOch140B
LhT9cYhoyFtJKFIxkXn8vH/qerDFm3vGt96yDQ7CSe1r/lMxDaYBFoEF/Xz7UAfGt7zSBcP8l/Nl
tIx5gERONTa5t9JrBYpZmrY5nMMcgszHs8U5zgmPgyXnfc/3+6iGkSeoki/APMb+8V68QO+vvina
xDgEPCH24Jw9RD+JeKKZnk5CNkz6hAk0n3ZyplM1biq2G209GibbDIgMAUUBt2BfOCmFy3d8c8TS
uGoXFmRSSnFzlp97pPWNiSVZp3cx2d530saAhsXQtQkCMucwpu6ObhGN0u8DQlhNuL/9Z4AG6V2K
m8EH+fjGF2gJZ+vlthY0/kqsY7Arx1TGr05iHBang3ONx2ZIN/+xU9g+BSRfHoKCzk36P3rspqVI
QxghdvHlVUJfy6d2AGg5jycsNkp+ORCXrOuKPuJokv2Dd9OJIOUrssI+EQFsO57ew1YK9Q5eUhX7
Z2KPrm0rqqlGrhu60lQleP1PCyrxrq6JJ3t95RqYPKOTUjWcZM0vE9gpnrNVT0oG2/VvYrzVirKW
GIV3lcpxT+W0c4unUehmDg5SFgWvD63i2KoedHIuOv6kbU0mxdIBThIutCYVsbxyvh8UzP5L+jyo
jgZXXsEHf9sg8XMfdMJ8gKpqEb7V2uR/wGhqOqe9T4+eDxX4kK7YH6czfAcVBGwcpN7lRPUuRzGm
NPHcGAT30M+wAo6u983yPA0fYYhwOXL2w4doNy6vscdq/kgn4TmsFPJym0ZBL8ttqd3G058ttQI7
CumqwT0MrZ7QqbPwfMzfZoFbmsjx8AiOfD7A2EKUhsQ4iM5uAR7B7lyEcDVOxSvHHy6GugJqtQx9
uU/CACw0uXt6yMIhXNlDo02IaMVrKvIuonF+9aWZh0U06QjB2sQK0bTD20dCsNZ+gN+/3LIp+OCJ
2fgnE7ogQMESp0n3glHzF+saauJIo9ClaRdUyYvZjNXc+mvYpM1NExsqfTSJw8fAWZmecfg92tVz
bn6kx3uMTSPsHEM9oofrvbD3Ui15tYuqeWl8VJ9KAv9M9tD+qJ9z7Kn1BKQRjpAVHgLPZYZW1rUi
ODM48rNoiiaPaFGM9qncnf79z45TDDKz2WTJEnXPxuvR+aclooIk9QyEttek9J2MlFAH+vU11BH1
mnKBda1tSKLSQLuZxpQyhN2kKu1TL2AqAbjfA2l9cOAIhJs/rnx8jOB7Pp8C9g91cuC+4pZGtDfP
OnPfwgvPV+iAFDBT/pJ9o8zleOXTklz/QF+zsIlEcDXTo/lgQJyunzw/HToKGFsEcD6sdOZerzRY
8jw16kqbd8m3c/uRCSJDet/cXgsaOzoO/n44ZYmohW5N7xTlUcUz7rxBj79PFG5uLEy8kJieInFJ
PpEL9j86MY87yZRBzXUnbdzojckFRhW/YcK6FQlLQzOEw0/JCJdkehw5RJuQyhD5fYTOfKRQjhNv
bs22RTeprz4GU3YM6KJV7UAgTbgBEJCAmnm3aBYxw3gllFWOX+FlvTVp4p7XVCIaKktlu2n8BK2j
dzd68uyn/G99ZB4xsjVgG6fxT7eTjsMhoGv5UG5nAX+wwPj16sWaMTFEaChJZUHGobvX+obh+LXk
7nLiflfVL/gmbhRPOBogSLuTZQUuHfJ+oVGrRA7HcZHh6gSt56sGmGt4B7R3Y+FOREv3Cv6dIkFZ
yPLJ0oLXlsgc8RH39V6hllQjYb8YtYSuBsnSWJTwexMkXSe2hSRtZPVQJKvq+vSehGci6KUwyDnn
OMvl0YWDxpVCLtX1QD5eL/agle4WyXlpCH3mDPrjyH/IOW/EkFc3ROxdfgF2xKSOVXop6n5Kh1/L
GuM90bvpmhSDQJ8tGY09QiPrFH7ULnV9jbDXrLP+qTVXAztAg0nhICdXyf7NA4qpSO7KuDGfay8X
rBNh2TEBo2oefTkLpPps4X82cc1cXhgGUYe12VzT+NkN72nAMQ/UEvS9XntyCzu1lKK7Ek0rWkTQ
rCEqV/6V1EjkzTYr43n2QXPpgQJPVfkjOtMQKyJkfg+cguHBLRLjLc83s5beyUkYM0Kac0xaZ+3T
ZAkJtfThNQmezGaIjyW9m6L3lkE7FlOcpD2knmgzS0UBSdHlWq4YidSlt6m8ZzZrwdTiPNTdDGBC
sEBTLfEDSIAjMJ9aUJs+EovutQaqBcHURXSraVbuzNS9QLb0FDUXPAtPsgCBqK8/f67EUiJu4xUi
6atdpi6TAqqfAEKNUg1fhbIlACdqhFrYXw5k0ROxytj8V+/mXghjhE97THw+swsCDAHUol4KmdNh
ZxnVfA0FCgQRzdpmoQtkKIwnNyQWCgKXVuFnOXXG4Ik6N+DgaMblx/uBQiM2XwK9R4YmySyuYWmg
vKC/T5LrrfJ5MHHBnDECN9Z4n+Mf9WumseqDum6ZHH5uDT4apOXUEo0DzehwaX/fHKSV6aYuSZHP
DTJ3NVbntEaTBqNJkFDiqON2gGKrtqS/WFwAIFgtjifvyrJBNvCDFcIgUQQq3hmaBALwBD/By2Nl
X90BGyd7rO8jj2m72cM+lwIeOKEDLwEcjT4xNrqyPm7mkKdDFPKoEHApAsjIhO8U/7o9YQTQlKkj
wR+8DVI7PZBdCuPZfwr1odVYFjB8DCEDev2FOg8fTvHNDURcz6r09bPUWtXq44f7RaM4+bUhkgJy
X7uytx+X29z3GRdhrBtgMugnAmAVSYUrLCOOrSkFvEwel+JU9zqrpxmfeWqygfbBxhEgloxf7b4J
kG3TsZfTg2WUFCoWa6DtQWKFhwNpsOx14OQaNwGIm+h75YHX3WevadAUEv7ma3cnRsK/iB4oiOEG
op98UZx8VNFbyYRmP7Dis3WN3bVS9Lfaw/5199mrqoeCvwtyTYojJ27MOecIdBNxn/3XHg6bCQAy
at8B/tLh5yJWC2uebIzDGMzifeRW8Nbx1+ahJ84Y+8MMmtW4jew1Mas9JHiEJ0ucEooCde3FgIqU
Bh1YYlk3trBeawlHbIeZUiG5LXGY3LsQFpXINGkhyGow2Kp5oqXmP30kvt+ENtKiu833FwlBZ6zu
ydYjMSJz+QQynktw7E7wDnJTQPUoFD0ns2VhLene4HlaxRV43Fg96zsX+NtJY8Q6FCVxKQP0idfy
ZiCLBQO3plh6uPl/AHFFp64MCdjxCZ/WeZsx1D0iZuJe35RiLQns+ugEL138ZAq+qGKBKepWaQm9
Qc5FYxMhWrwTuPi626WRes5BpovF1r2zijGI7h8a+XKswJkNdD9CqLct25khQqKrcLi0/rBDWcW2
CIH/8b49THhZDQZDkSDo736Pm46hil2D/U2MG2FZQTSBr+8tXSCA3fOmnfk8JVCURegE2Fh91HD8
ZNNpaZNDIh3RlSgKoJD+khe1RUu7ECeptcQtrGrbDznmS0C+KbrnYzHc/FkSPoxf1kAG3+OCECvA
TavUy/m9pU0jyYj4/N2fogzLWmxQerFgn0lrPBYhSU3AGn5D8J1/93r6ElJGQQhyLnoqkFhEkw2J
DTsfu+c8Irr2s8hKjaa9PoELlvh6X9DpuPI2ARdWSM6jSMeK+NqpoKdQ8icPNCwWGWl0OCzfadEe
ou8yEctZklRa6JIxEWc5dR7ds6/h9tQbpRzrIdysgdzXWnregB5ziYEFsnVPM7F/6/NsY3b0K9HU
HdIEAcEQPTV5UAkec1Jj5bLI3kfKEv88AE+sZ4sNQq/n2vsLmkEPtPrHI4aYot6HlPcR57xs6MKc
Wa/rPHumb6fcXiM2hxuMfw0PRUKbftJPLqyFWp4rr+69jXoBMBb9nje5LJmBXLd/yJKkYFxPMbVG
wuNZQHhjl7pkHPTDQHiad7zOCDpqqpZ9WF4O6+oY/aGAdD0pPLp3Ie0Fn5plLrJN/HfrYDBVxUcV
hwZHnXySk1pzGjY58gd/zuAUbUhUpWVWhO+AWOE4NS3clyiGurxl472TTfuOwGoesTjSWzNAw6aL
cxP7+Mvo7QsUPd6bN+L4RdxXYB3s86F6bHj1P/lufRKdEEf1QkhpCREhncJLAV40y8nVWA7yDahx
b/LAwfJxgntbrt5VJjM6H5dOE/X2xHzqSENo/xM+wvHtLka+1P/2BymghVd91tSf6ydVp6RLpS5o
prrg6R/yoP+FWzbembZVdOvobvRGyQiUqO0GF1v8R67UgP0AaXsNhLW0wB0jo2O0r2WKFKhPyu3B
5mK3ayJKX+oGMFSVb3XOpDPOuplCBuOtepF/UXb07k9E/fc3GvK8Ha9DjSRYoMWM1mDtD2/P0884
LSDHneJDIHRWmLAIhbt/BcKMFu0fxb5bDB4PayJKJxcNHh7CFMVUjGfX7n77fax+ecdD9VVj0dej
Uc2gZ06jo6N0aN3y1z5DMc9LppD4TwBf4JAG1L7gUvoq4iwL6YsSU83Et3Bb8CUFCE7Imi+xRZ/c
rsWeEgzh5saIgmpKCXONjRpOjKQIIs7GJqeLbZcccXijqXlneRpIw4Yj/ABOASoFp9yPNCaVT60v
UbBsu8nmaraXB0w7pgcQCO5cUecXA7aJ7kql6xvk2oMGuuTbSxvlDneDUTGW6JsSANDExa4lHPg9
Ldo6RdchA8Lb3hxQLUzAJKnWquVNqzHke7ypCWZVnYLhuhifN01HVWDwG+xLoFCrUGqAyVcSBLTf
FVGCagXnWLHGSU8gr7B6yAjZMRffoo6OI8GE6YhrRFvt+w6uKXkep7lkXo17j7HnXut1JJGNrWDf
peefYgYkxDAy1nmaU63WRLACNX7S+XfvGfJEiloCPszIb6ZpJunPt6/2yz9jIoH67uy0oPsBXgam
mfom4qaad7y4/x16NJgdBYiaMvu+ZtcgCJbhjCwGcj/fEkDltdgPgb0AyTGwkMK4hVJI7yHuL/3O
3ArEWtWiYgOBDLRN8f3v3KNFJqhfmL3VuysWWTix9VuLaC0Hed6Z5O3zOECOBr+Qcx12t0YxC9v2
lB8VRYmEc6/Fz26tX0l83MGiRwXtnzfg1GRhAnnXN5iHemU8NWSE61bafWwMBKz5V6qAqTDFXq0N
PYHFzVwESD/0NjYyobTJR1QGuOkOVF04aUWwTWAVVJA2cbcyC37CwUwlG2S39rsXUgTn4TtZDxnT
5ruVkIm/C0xRat4xq6c43AaDrlox7FFthxIH+J24FT7hrJf+rNqS1EVAirISkOy0n003JWVAyZhA
YWF1WecJInqDbXhV6p39V/FzMAusv2bHKvKDLb3gEFRpZW6zqcIhDr0epTtQa5zWfXTjjcohDdcM
slar3yBjXV2NyzacsBtutnqYiIbrXJ0xNCfOlQjJlyjKtebhqdWSkliARLBoIuURH+fAxqCPQjlx
koK11OJTe/KwPuORqLKp6PEKef/q6Zwq0PqM3Xj8zzCOa3goK3yUMqTW/aeuU23t43EnhkxXV0eH
c8rdMuyu++YpUdHXRiM8Q3xINElfdm4ka0OHZgW5Zhq3tqltZGWpSQJFVGgqgzka8fd0zLT99VFx
DI5joAxllIeoLDNlO0Okb1T/OU7SSLZCORGVIWzDsi2dyHCOR0vjWs+U/eofg8x/4XBMk8qPENyL
fDO9bktj8UDSKLtj75htc2dfQvevCBz4irdE0BfBYByU7Yqawoof8+oJJ49kGbMujDG/RExhsaip
ztblGisXeHPMXyr4FdTJ1sXM+brkIQGEVnxH06T0RYvjD/ZeVv4xSCwfwcvuLAKm7G5Vm7HugND3
zuHPg+x/ftthwYPL3AsTzQEdhegAqRhzN7slvBYsZP9iHC2RtjMQ5n/CYgaqRoW+YfVHg/aWnLe+
q8tveOBCB2Q9OpzZftiF/8PwtzRKpPQUuMC1t9MdHXk/dc/Ehwiqk9zKAHIYxBsS8KY3Nb7Itc6j
qwgkeHGM5+Iymeho/b98fxoOPMPIiH9HooBleLtzxxOhue18c3Kfx36LHCjblSlr0YKZ9hBb/gDb
OjMqQtAqerCEX1xwXBeS+Nb0B9QG4IhSRgdfHPCIE35K1G8xsjF0irRxGtHfxoaDmeUXTU9X8h7p
6e2dIodSW8u+18SK2laA9RV7z0wm/6h2jdhEiV8duiDOG4wNFOjJeIT3pGXWMVS50sbROMPrTU3S
2V7nMsmZQ68L5r1uF5vIUC+S6EGWm8+kRpl2YvgQBC0/hqtGw+vZF5IhkX0FpUwJqfL0AP8NDV//
QlMB6b9axVs4j/NYEaFEFy4n3+ajjm1cnpq8zJZl8MVLa3uh7MI5AAFCvrRWq7LLIj42ls0rZgYF
660Yf0ua3rBdrt6DTnytRtXjxadljII3erv+5wo2lNtjVkJxx6aE5+GUtFqlR92YX1mhOh23BdRi
eZDY++Fj0RsNigzcS2k+2iBxiG9pvCdjPX3L3/aVcg3nTODckDEQehrwJQXcWnyrCT8wHDiYqmK7
WP/1NlMyINhatr5S/SnHKUnC8G3jSs1ZbXASoN+HW1BXUBT5bkTwRsz4QsShrDA0BW7kz7aVrEBb
nAoTaxZ6+Mu/UFb4po7kPzBf6GcoSc8W2EZFbRFuuVRKSfC+RsSffluVLUrKSxI23ztM4ijKtZkV
zucedMs1vLHfxj9n0wg6ub7rYriKUQNSlU8X8WrmQ/k5A+bkZemSQFmjhxuqv+1OqBJc77jNP8IV
BLT6mwDbTIt1dISfYNrNQX5SpQd5dAs/FkJPP/MBvmc/dSjJC5/Q9xKeDgyErwILwO4DnaPJlxbM
jKw3pgli2KT7tbXVmwCOahn7NZiApF0XW1byvckF0KE2DF4QNdZaa4axtHlsu03eSn6PX5flaH1N
xNYQKjw4dts/4YnhYdgYclqD/GA1DsrLRXrd9phy9QqrtVu9fVY/T2UMATkgH3sU/jrWRN9+Wk94
dMdkCryjuLHxZ1YNF0DD9Yntk+RI95uQ27wztVcvsCsA/rcZoyWInIru2s+biK+ELl4XGyB3Yypt
+KnYZ5vEVhU33b5qwFOvM8Diptx+AVnMnVS6eIgduvHEPudmT7fFfLqZj809TTmsBsWiXayXJFfN
RwomrcX448MDyYay/G9plhxs3KeYVWziR2lTEJCAH0Nb57wM+4DuQR+62Tx75dcyavwRMugqsf98
jmw1sPVjuXIm+Lhdy1bQ6KWt1BJ9DJAizcBLF0hEAvRKGtW+M0VFyj3WuVh41gYNK3uq4XBsqy34
CFZALFS15XAcAirD93deV4LTC5grcQpMsffAIoJEUP/Wss+AIolslYryFdka7F1tOBMohLkyHzpT
V+BIcIHBmh7yEKCzsXk7DrZRS/QNEaD7wObnr6HM3CeOQMNDS6mc1MkGkReC15Z8AEeXJxeTzTY/
r7dpBKlb1g7TxfjfOVJCzuy9h4zpULd5JF6xdAm//jxCTfXhG80TsXFgSoags/ESiI4mC0nSDauM
MF5D2ArbRTzS3MLQ7rvePmmWHONAESeBHvansKIFn4NkNF0h+hdwx2OZON3kmuRPAJaJMNKglswi
d8rZvp0Arqq+S/nWV6+IrfT49epzfgfoEOOXtOIcq7CxrMaCafsb6uKWF1Tipcd4Fdk27ya199MF
2VFKf+wjp/M0VOe4ghqwhHApr5SG4ISwfDaCoeddrclVK37TQ2E9Z/5dmpt5+MShoNhEvOHDqJLJ
8Y0Ajthde2OZ0CAt32YY2pH1iwPYHBCUDQjKOs0qS6HRA21B9PK0DDd6hcDHrHP/U+9eo+ad4zuY
eiY+nHp1j2eF7a6RQlaPBYcJE1OGYO9onBT6X13g0i4wtPPGQwrVaWggLmjXtgXhRA7e90Kx5cnJ
pBQmkN60eHSEtpoyhIYUVw41SSS8xMHdaMXNAT4mUYFAaEmkT04ifYO6cIgaXGGqFAAOiQg1Ba56
kpTF1ncp2N8z2twU54aJhkSFKDP+XcTYao8jU+sYFtT6l/Tex0Cp8ycFWR1jmaYSM6DZSW3xm6W5
TPmctDU+wJP6dezGzvNEVRWAycO1qycWokPDGVuHcQBE/tgiMVzLhGsxzks8aLk6ZrNqVC99UVtD
C+e2czGUWFX+P7wsyaD4wihskyky3SizmBW9r+GpwPto2PzmllX9mO3xyNG/eYRd7CFa9kouJ53D
h4DJNWi4eMkoIpC4g6IUj2VK3XZo/4E8WKlZO2pB/dIUUmwTUy1GL9PquMtM0pVKws5pfY7XJLBl
1V2Wk10Lc/hZ86tNX9TW5YDiWiZ9o2nCvqDB9n1taYPEGYT2eylav5XnzmyYXHvCAqhP2b4feuvd
Q44jGBWbgvoqheNpbKCvwPtPVTasetWhQVJsMper4z0LJMoSbpF9C0ucGOdwY13/3D0ysTqcg2xh
GaVpk6oHH6vVYcIT9NK3wK8lXfeibIz7TzJx3fXOz8vlMY23ydQx0dXqPFmLpzIQiLwJrrNjSVfM
oLR4kaoRbnT8VyPw5yFoJsW+ZpZghDh2sLdVkkX2jwIqdU3Jveb/rYyA5/0QASmbcWtvzt31HIFd
RgCKjLnYQYBbbR3RKWPA5uJq0pVYsvLqW7mA+hxiGMuWJeZll8qEfgYJR3pxEb3CnlpYBPwQw+ad
U7jXFvF9/ObURP9w7MqHzeWBcj9eZPtvj/7q++pYzJ74Lh+tnLdT+rwOvd4ucZCqroZGuVMINQNW
8LZIBt8fPsfBp1BSkb8lKxUgjBUyustB+WQj7nyIHTgz9VXkWH5snOXCUdKZys4Vf1bXEedD4gdY
fYl87PzkzbCK+GZM/haZFs+7tQAQzOBpVoBKNlf7VlyDuq7EjibBA0NzFRrNmVtaJmykrhsxNAS0
pfBtQyFQM6TSct7T6be0j1uJ9jrsZh3C+upqDPT/jessGQJmTNo7rWSWboIVY6I+S0FPzvl3dsVF
hYMU5Hv/UI+ibQxnhlwqc0NEJIuGjm5xsBthL4/9PL5REyBe0xmecLChTUNRxvZaHtrEfjtAjoHU
MJ052b5PjuroZ4narXXWJd8fDJwnz7p8kkwEOd85BAP5rhCz6uzAK1HZrOS7ax+cgFKGEs/RmwM5
c2XYJBChkR0/bKZicl7Ka8ODJ2MJYpBgkfJlRVarPMXdCCyDWlKcht+R9ZmO4gV8pwSAtgY+D69t
R0ItHKO65TCqY4IvRKrMeSC/ZERl0LSaxMQ26nKZCOq0k5pfoFiGLko77Okd5y1Rpjn5IYll/SYD
Xij7/B7a5rBzJVoE7Go3a4E3TqCooSd2+85aNiM9/1pNw5bpLSt3XkWZ4wCwNncHyML9E1CtW+wE
AV8j9C72ttpz8p7UxLevfeyRcs8GfP/vgKjf7sB+wPD4jUMZ0Ikp1qPfjMhL0nPmNTHc1RhTCrYy
jwCDvCd8bEfqloIJV5AE2piEtVICxlZFcBn8IVKisXPT1jMflYMa3YiyHqxw4nhD8Jfepv2DpAvK
oPGf3OWH3yo5bv+cAopi+2HqSIx6Hm4+mQaFAfyT+kxpzFrYCHPGDirs+7MKH1fN+hVoKCup1EBX
x0aNfCdimbc+r3JtZXQ8GFqDYEhLLi0YDllHjSaw0bKX933X18t/+ZjgrRuzr4ySYgXJyt+w6N76
yFYSCWJWhswJVpFLndhPw25ZpONJENc+c59wwGXfX4UL/lPU0PHz86rB90CCnU+bY5QgCe9vuA5g
7w3f3H1EH6r80Wg2kdbEeFphlVGWhNy0PPhQ26/Ud/fpO+OGCp8gU0RpdFqpwXVLfmAk5CSiOWEG
JpP48Jh7NeUHd5B92eyTI6hD2QgB90DxdGkB1NiCOcnehP7fQ8R1SBJH3Pyet7usKpEcoXa+7oo4
BaDjZdchQ0JDtI/uVC0OAbbieQkxQ4sPmYXzyV0zUfDiS6Qb+3zll3yqG3bqcWxgELiTCfxY00xB
FJYEyc1cBcW0UeD7H16gas6CWrNBfj8VdDCx3FqoUVikzwVdINWC1nZrjf6+SwV/T9MVBruDjIt6
+uvV751f+niSlMayC+lskst/06KaOqzxiZyNowiWIh6mHvUtuYsVq96a2+A+O48u5LnLJKclxiV8
Z/x7w13TLOKfiO4i4OR5Sa9QLf0poDTqD80C841eZzlOXVHLzj0ekojjg3HjKdGNZkee0Zzx/8H+
qXPWQh2DgGoPB53HQLdTTEzIwtpn61kepZmg27dhmf/V/dHo9ICcEx/MWVdQPgpgXuza7RIbqazv
cAD43tkCddlVzSGonYgqIyNCQUOWNNDiWcrqLXETEWpXw5XcpHI2DolhUOkCt/+Fbv16rMbbxpWC
TNP2AYPHvGqXR1tCQ1PGFmUv59q0I5Houfgz/9lB2PadgG23OST7380Hf6k/kYIsc8PdXnOKg3Jy
eb6Su8W3xJhjFotHe3c9nOLwkUHxY0xn9QyNl3cyMxKjl/RdGStWhNgZ5quGOpArfFlC1JGQirsD
t6ple79c6KG5AX9mdqnqeFQY4MmQQqjMGrYtzwZPuHpnsJqJyN+Nj/hJRLy/oHSflsGzy4uUaSCm
UV8jCuTgoJJ8vIbCyasGacNPL09ZOU9sEhaG+CyL6H/rG7y/eKmLM/uUxgSl/Le94w8kbfHRLvzq
BlHnx4oKIWQzhIRvctOewZt3x/NFXk0xpguGw4SwvJxRoJxcIkxOCpo00GoGXu4+0jPxCC+YKp/Q
JNgAxKEinMRVYujtayoFbtbCI55zUBtFMlM4jsapciauExceYUjCByROjIWcEMsh56PReklHgGqs
amt0Prqm8ywS5iDCmM2Mjfj8OuKLLsO23fDkNba4E80n5sP6cBEuEYBBblDzMP0OIFK3oztGZyLS
txJDAPCOeGh1Renu4skT6JkKnQcc/GT2SycI6+o7MJIb1YYJ0wtAbXml6mmCw4762LO0tZxFX2i7
wRdp6Xixb0UUs6KPYwdGj8AzSY4RdKqIa4Dnu1MiR/gQ8+TW1G7cST+cAq1KDqfa+F70RnD0wZgq
KWUMvD7tHPK7FUgJjHajpCz/4w5yPtgbiqZfzaPBNDYj06+C1+PNjX0xKkhZRJYG+XWBjUH8eRe+
unP4YSi4odgli/dLAvjwj9PlMdvCSN5a7R0t8/YcMskPJtDNXHd27Nae2tZchbSZ+M/BMflvsG09
JBTckgxW9XZlES1Kp66OuLWzW0LOhhN4AvRngpRKzqU5BgHAoHq9S4H+C83t3iOk9VgdaUm+lPhV
4ttgIy3sMJSH807cH0Fj0Ezn2KNDXZFZKCP2RjHZr/cYHeuj+Mh1sIXJT3Jjht+K9Z4ugGyCYshB
/yiUwaH4hym/NDMj57hclQA9eTIJkSH/bGXisbOrlQQzjH12hduZHIvZeGwP1UN7vSDUq5tbS6mp
//J3TMIn4ZogmhJwx3gB/3hCPEQJQqIDj0iregsYeVJHUcgsSGR06Pal9sh6if7O7SrFb7jkHnPC
mSMpW/ksPVjNyVIiU2RJnVTCSuwy9oLPVdPFvIXit2uIc+lp9VrCyFwoV5glu1cJOXFKl7PywgGv
2eSATQJz8ajDLHhsV9/AslT04Z039oFpnxmk43GOuzVBluTN9XGQ/N1VlqdnhywFt8z5lSAS1sHM
lda5Y/kGHM1VwZ8653ZWLhoMT+/+MaC2nHGwB7q23OZT2nXCdE8/0LlNZIHGdg0pQTbQmqnoGTu5
H5f0rCtjwxRt/+ZrKqMZxmGpZDjx+AJgucclJqWgGrD89kkNuzMNKp7ZHju4NSbUACInCk1kU9mp
11zmduMUKCFTdg9NMRFNgkipCqp7Ii/7Z9CC/VdFQ3sCfd8Tu7ln3lt4aNUj5LQrz9iDCIm0hukU
YBnP8kEp1C/LmlDAPuPoigU4Yl/7wVpvLtSzULw2UsRv6Yll2YV44pKA+pl9+tS2IJa61zjwaQyv
B2XMfuR7OQoc/8CAthrkJmRh+w1/aKtye/xcQKwebN/lIv7HQH1eCKPebxoou7oD09cxB8oB3OQm
4QzpTNc9O2ccZTLM2ipZgvd0SfrPkjSbx6Jox3iogRxvrX+1mzl343sLMASbcKKUI4RjRkSgtq4H
U/oO5c4sm/aUmMPsqflKm84uzuNwOemFWqHei9GPs6L8SGm5466sR0CVniOZQ0bM74IYcS8IwXWJ
0jebSg8PF8Hz/BqG/Vr5PJpNaR/mLh9SXdwcPRvcpImT+dKBGe55gTAIcwqQI9igjDK6nYXwkawZ
U9s3rDWbAhLrSXwfkno5v1yY3tGNfISB32v4LN7DBQMHbLUA+0eHMq+idi4BFJpaDKU24qzV42FL
Zk075rRux32lZpotNc4bKt2UOaHRkbrNW70hfjipIUQG2JYCqd+hG7ASut4QMc7NMDhYjvn4erf6
sh07+kAUwgCzCbBu57aq64WkxJdOEnRsABUh1z70+TnclKSDuBwMNJ+I5Ig1wT98ktPzxsfiGJEk
oYZBfeG6jWku/rS1+Vz5YFasPxkuV5zQwjJS0t093q9YoEECqzflMd1vYrUd77jeK5RN2Ldpnd/Y
D7+f/+JUeIzUtaA9JXCvwXbzgPh7O7VvR2fu1Fg+YfyiXL83h55ZJOkdcyAmeHfAXl/oDNBGXKP1
bR9v+S4jQ34y2N2+r9Igc4jA2IUMQSJaD4Q3uS5Kc1+54RcU0eYJvKlSWyKUl78YptRtMMoxQF0Z
qwJ4gyItTA8TPVHpmXaD4qzqa0ce6Hb5ep3Hn6e/mzhdPt9ii7S9RcNJScNUh9gQKPWtbh4xrsji
Tk+bZRi3pY2rmBFAoQYBN6cmPpmX/CUXBQofYZq7sGkIY0vr8MR2npzx9KaU1T2TVQOi7hUuucFA
4I5HDfCOOkuigT1RcK3VMLrxQxyrb24fAtnWgC1M6eQm8w9glnbd+wIfL0Fba13fA1u9EgVJJPR9
0pR0tIqWRH5CBkXeG8IqV2bRVDxIun2UE4ulttT17LVkGjj5PK2ZJkxIAmBlqjBZq7L4xQrYJTwA
OzNO45nCi9hOPNSeM+QvarYnAs0jIuMZkL3vHDqpZazZKkiFbt0Lk/vsmkNDJsAGgpWtjnZrKy9K
7XgegmMXyZKeRPG3PBi+G5unvOTK0V+PeG2y0NS/vX0CWjXs2Pg4xCwv3zcxyeXtZmWoFKJ/h2v3
bdvPvi1NXOv7ozJMdTyCYhDxC2ulmcETGO3SUUqFQ20XE5Rb9lmBm+upUxOCHJzYxh5kP0dFAJFL
+Wsr2DywKG+Krn/+IfSnif+A1iKu8gRNr0vU2U4bEuNRqI/ikKdJ2GR4V8zns3tj11i+Xqd6+50A
nyY7Ilrpb5dQOcy+F3QxWJolEil3+WrEYFh2V4lKwqmlZuv7tfJFk3/cCuL+rt8i09E6+QfLMQTP
dxVqIQN75n40OCE9xjUSwuAwHc1bHGHiU2hOWI9UXRgf0m4RUaAmWh+deNC/lfZK6LIiePeBvW7/
HHCQsD+43Wsmzf6Ctzt/VXQ/ZzZ7KHfuuLpSZiJY3FOMUKDB6/dwKIQunh4JzIcgu5BGWw97CTfe
IToToa2OZl/ylB50MQTVnydnIMb1+mNbccR2gOnGKctFsGlJETLUiZPp9+kf+zgmSkpb6cEWYd2m
TqGUyjxSisJ3GzVV+OXztC6EKU3fbH1szCVTKNasEPz6tYgSSgnpcW9/RNjNogD7m2XXHJI2B2Jn
1jQjBRgh9ugrGC/aYyfzyocuW4zW70NRt5vgp0LaOXXIf8RNFvX6NTIJIxxxPcQYCopWed9s+wpM
f8mZ7yBc6GKRLm3P1v0ntM2iKRb56pyf98Hp63dsNMIg+bWW4TnrRPe2Iel1r8b+FXWbYAF3WH0n
K0dk3HQQGAEz90tAv/iP7FP8L0xVaZSZP37aZ1+XyW2zcmnyBre18OzpBM9aplzGRq+oWbA26wIL
uMmcKnfr6F0Tug9xLlprcoiMIVTRHTPNZufUeXKDXu2fBil2RqeC+sTxLHC0LcoKoFJixE2fRTS4
1Rxp5W4Ul5l1C9tzpXtXjM15kGXzvXF5cDD5cTTk/qABLST4bbQfYQn2rxX/dSBexlzIGZk1d7HN
9OPwDA2vQ/+cCb8X2WV3gWgeL2+vfd5J/CWlouaybIIIGo6JiJTy2s5hd3SP4VkHj3wJylzl5K+F
iHiDDt2oShhi/NBizVNaf8v8d7j72WrFB3GWDvYLZe1zhBUkTiHXI9nP8PpScJoQlR6twzVAH5OO
/29WKxr1HR7grr0XyavvKpOwAjVQ4bV3awVSUxJhx63REK/5umofIe6rY2RFx6VQtKzxo0BZ0S+W
DsW0cgwZcKuDU466LZZPVMOKOV+VruQ1xIOexjunHYlGMCbc5r2H0VvF3seOqx+goZIp1ZpOHhTO
R97nbzZvyyCNN5sq8k5Tp6rk+CrSy0dZdAbR6f2sXIvB2GUx/ntXmKR1ihsQnk3oAlgqO+sIC/GP
fKhpHgEpd2FGxIAaPhxh1ToEFjbEl8Q1nUOedg7YxYcJYZWfz2X7smoPMOoRculDYsnL/X0duAxD
rCb26zNwa/h2/OmmXSFhr/ptuzt6ScowmvC/TYt9YH2VEu5vk5lxwsiePqQmdQD0Jr2SNC5HYQlm
Pl5uFCibikTlOMemrifOIcFDzikJMHcF5pAS+IfYaDxBfh5f8IUW8kMWrHpmt8ZdWHPm7gb8oFVl
i8UGHb6av/QhiRe1jckCfIbZX8x/zPYrwklVuZdq1pniI9uAyUL+Fk3T8gvFbA5Mw/EaJXq0G8zm
TIHT3I711qTXG/wDMwKSD7BMGGVZtg2MPYhhzCR9VxK7jvZt4JzbPsAy/+H3k/QukPqp+LWXYIo3
RFI8txzrGCZzT4t+E9nAmtD3iX8jjw/mtExZNDS7fdN5nd3gUN1tO+Q34vE3D+Vd5YJa9AmJT0Hn
JMl6tuWaCMkg4m1mnQsJ6MX+O7SgBGYa/ym7dym4XJoSYy3LJcBQXpIaI1j3vaYkJ9Vi9NxUh2ID
o5q6F13QYk95JtfgC3XA14tjdyhH8SUCyFkJYqhIUK4trXkoINt/bGvxE1JxVEl7Rf3KNtifesvB
ktI3kWSJs9Spzb2zq623TPYfeBBljj3D24cZFzUxone9PifVYvSpccU2AEF7Ugwny+yUNxLGbk6+
AW9AutarBri/m0RtT4szNsBPDF8u5JYTF+w5wDxwoU83OYe8y7JfE6EgFH+OsTODurRSRJQq8j4B
ucHE9CKpJwNe0cYX6YnJ+SQeAuHzJFnLAaG/QSBcUuq2T/VIFtE/817ssFikjzBo0BXaG3CaNtto
kkpn/or8UwgkbdvSepdRg+UYsLg0TXaLOzUyRDfDZu0IOonq7eJYifZrJ3waOPadxqTJlPAuEVx+
v+QGO9fcoYanjHHD9BMP0sqlVVDgGVAZDzCgHdsB5tsWlLY8M/7k7JIhPbfk9vqIepgnJcJXkLC2
hRAla2c/cZraGQh6YgjPldl886y5FtwNtP8DAXhN6Sj5BSUDNXp1BEAPQ5aLeQQb1V6DaqSknBuU
zWGhGA3MUl6QC+NowequBYOXH506X0tA5soQBzhAOXibmTHUHIRXKzhkAwbQPQLO8r7IfO8a8H8J
LPA5y8FM3dp7Cy8T94e5ShsyH8UFIjzN1SYJm4UDNImZ3JJidy+sqg4uVbTFVjT9VYeXnxh9jPLv
XcAK8zme6B8yhCn0OB9GB0cnOSruTfy1PXHBliRNLBKtUVL/HdYANb1JWZGd//bhtw3/7bcjgTqd
hLvryi03Y3/d32z3mh9zJ6LMGlGX66Q8NjrGvTzckKGcFnbluE5BsZFsMa7RaDnKA/N5Ox/g6qVo
WPpL92vk0kjhlH6h3y8vj5jwbfzIlNp/EiDZDwU7bAqXv+ntze3zpfPd7fEwEdNfkGxwtjh1jMHF
r6AwjAJ8bsMCA0YDX8PGoUF64GuC+jzzak0INpMJj2QhI3gkS0Q85PJsReW/cIE+WYFrNBSAQiLM
42cxlQ96KYbqetki0O1UcAwwB338rf7mmggkxOj56xKIVY6rP+2UpGezTLs4R3IGMr+/qkQ50nNy
8xvOYs6AgqTTEcYU/eFbidIS5ejyGTAyYneJgBeyVdCQT4YS+rjsSmyovYGj92cYYaHkugiygRvw
jOW2kUOmaum1vreEEq1Vx/3vvbcYMivQkXIn8Y2O/rfePBzhIGPjpAL59W3FToqI6bYGvdZdziHV
qR4P0A7LJsOciiMhSg3XyflGdfl6elRsaw3Owe4KZF9icUGIGppzbR9z0uZOIpi3Fh8b5BuTagTp
XwCxMwFCI4q9EVZyIf00uVdCTKx+XEX2r3/HiDSe7YywBeocU3XJ5n3L+p/SyOIIWtJScaS4nYUI
m1xUMSfwqtXuxisR80Bbju2pt/RuGwWEaWY31usCxpn/ns5FEaH/c4NIGK7IxUB1FFSMrFP3+LqE
KoswHUPF3er1jQsKMeJEMLg6s0G0CvA13rF6MoI1N7SrmBhkKvlwcxfyQb+r+Rz34TIoPMQYJCaR
QT5g9vNWHWLlIgunv44idjIFlUPKOLT7wCNH9qahEkCKTeZvlirywuMHR/fmLfDTime3gqhoJXSe
ftyLAA0ihycUjr+f9d/js/A351R0Ya9TZdkp7hUUzMMZexyZBlc6uyacLyhdFAumJme98iXIJXQh
vc44G3DyET1UJqekbHYL8SZnU1C8MCF++beGN51xUBOszcrfLkjJLM8jiOG9YDw3CZvNnzud3QFJ
rKC86g/bv6gNKYMgPADsmQgDe5TXDAR7leogtO2Hon27m8gyidX8Filwxtzwsh/YzTZqVLQ7EHY1
9yjIaWTz6/BPooo463kb28xCLcnC0WqutV4ufgaOAsfHL0aC2DYCe14ZdpxWNlUbmUHQrdYWVKO4
zMAbLImDwE+E+qfwf25tLcxiCGa5rjDD6iEjJBs4y9DrBCTPQEsDgB3bXpYDHbzEL4T2SmjBl0nR
Z7I+QeNA96mcJtt5UOTl/z687oFnIGkp5AwsVh+O+pNIJyybQOrqsFrZBXhuf12dKYJw976nyyHC
nJ7K644nSd1uwTghEgw1R8oHONFYQkaIMHylWPW8ZNFNdF1JugLusr1yspmc0clcQPLLrPpD/ZYR
k3FZCXX26D2OxiaEqAt0dQbyo75GpF1dRz9M34hnpEDvGGAlZT292K3Y45e3lY2uuvPCpdGn/qLh
Rwb6cZmzbjGB1wqE+P+si3ir0gcP1uE9uUr2YbtZSEh/hdZzvlw5tJRgc5WvNPP/U9Je5WKh8As/
+EggFaQemuIxhxClWZ2MvAP7phDMoafuOdrVK10iQOPV+7UNDw9DzYUbRT94q5t49fsyLlpbm23Q
gZiN+uO16HpKwGwj0m+BAehW32AXSnQHws1mRXOoD0B1wrgdTD8+oeKy5YZEoppSxEYyI5SIDsiE
sXGzhRoQtD6y+/Pj0abcU0z0Dxj2m82LoPxdgbIHm5IZbirO4x1t9l69mPYPGRtfaihq+unJp9BS
vh2YPKxd/qqelDbpuu1f5SqUh2duE5jJe+L16nFzmPRcoF+JLCwx9+MWU9IVioPG3AuqpjrNEMqh
mhpw5ZgPq+7HIoP2egi/qOGo0MFxEeHw+m8x3epXTFixfzpTn7Fow+6ZW+oSBphtEU2iuASuncZL
C8QN1KouXLeNzQpfNsezAcf1Xy58PCZwVM44GMDhICEj45lgDAQaDWJLERu2aMHON47hcKzPx6S1
CFy1Xmk2s8qoNfqfYvFJq3scjb5PV5Swu2SJhWaRu5GOmeKZPQE8/CCw27rD7N/CBuPFS8msdpsX
uHuqkR8XtXB13oQqp+xmO4c9wDU/OgSMrVNUVYlNLUBHnDihTpIPDfIyiT8C4DsTu226Q2V9fpD+
KWywa+H3+vBRSP9BppNa1yrLhwk6Sp9Yc657xJmhkbKRVmn27/3WFiZuL7GgMwDcU17qJZU/RqfD
YcLetCr9EPRDphDrWzkvdVO8heXVMEtPMLsAHg8TlzhfLu+XhNFiROk9s0qdcMmdYHpg6kQyRQdQ
L/dIRXW/3Q7lDbp3kU0ucLPZt+Vd/ewECwPU/q2Km7u6reSD3XrWClJx4FUvXt+5yytvkiwfykPu
cPCjIybfXPuCsZgRcyKqZbuivQ0qnQ5fPaqaeZJ2hWm0xtcN4mbq2p41Je8d/s6vLPu0cVVvMIN2
7HTo5FcEMpiTb95EzyR8VdLMV6nyAAOTpk4fQcPKE0HX3+oGr1qfg8FEak2mYTeZqFlRmyJrz37h
Af4sizxwy4jcj/9ybkJUHfdGA1bLI0qKUAaqlaEVaZIOHLLJeCCGAkCcrg1bBN/FXOaWi94ULkvN
nRPqneHjaGdK/fizDNTCSDwSxK7xFrW5ZQEgwotBEdh3GblpKejRyTfVLMGNh1WmDT4rugTY1aKb
dG79EiU8WwRJs64Fw70ptDb/QyGcjCnyoxFcgZ3MIpfVi/c/q0NCFRAXA6rFqf/d0Yld+6TUHEZt
PvCZLfc/CgsyoFsQ3Cfq+jJw+RW4JNssqCemwfOzVPj2gPleOlZwCv80IVYLTI0R9MuBgW49Y5gJ
DDj1NCT4nXxstdrkvIMlmcAB0PTNnOSEjl0faADP3hbeQ7qDPh43ngjadmt80KzQX0QCYUbx5ool
EMeBXUnJnggn6fPH2sVOPUKtUmAgED40Mfzhimas7n9bThatfh/ihTXm7nGWYdvb+lCboVHzBL+c
C1rNDKX0Vm7K0LoIE0GzqCd6RT05HDQrBePWJeycxwSE54tmjqXhZUEa1DrRV9kswb2rEX1fjebZ
WlhzIDFY0Hg0BWJRlJYMyHL6AJeHz5iAB2JsadB+j4FOBoHAiEMwIZg7yLOnt8j4grEfZObs/Jlt
8HN8RuSWF3FDoYle3dX5Y2zvs/RSBvEW+KWd3u65TnpndGa+gSMFxHbriKsKRH8fEEVJnupaaVJn
9nFzchxm0eqDsw1jsrmwD7sFQJfDz6qJPCo0OvWCCPCWamijRIa6wVnEgy0sTb+vydiP5IqfGluw
GQnUaYbmFt3SdsOb2K+S3U4vFSNxL30Ms2VqNQ8WOo6/nZvfKqpGm6NsNKDv6rmR/t2si2vCnbBc
11IktV8xdXT0JPKb0/7t1E3YBJD43IrKTPBRRrtwGG6wA9QKLh77wH0dsGr/QScfuIUgVXTz0lPb
8bDXz7DGdhw7mOXyWWI2JCStgtmEl51SVPzE8WEWbvH9uq90jxYPHGXm41DpMqd41Emj57joNq1K
7YfLsGHF2X+We1QQMbSYhZuDPktFht7Hbu2jYiSoT5zwkc+zZuB5l7nzzGtPS7q9aDsp6ZsZLd2C
6oaFVIoQmck8qZiBDzXY26CVinbEFHyzw9xjv9OH4BiOQ6d+RJuxysHGFEll85cKaciB77sFVGUF
HYOlR/TTmLQ7hPwexfqWfuyzOVEQYak+0GDSfbZ7wLeu4BXLxR3Fee5UKIGTdOfLe22JIRqtflbO
4HV5FNLNCCstv8jnm1S2BMmQ/xSpfahbVCcQljTppbJyJfOGqKdhp71Wg6VsXGi1IaS6zwcCgCQf
7UrZP+dZSp0taot3j+zY/0rRDgNXMlZ6L6AkrEmIc9f7SuuouM6WXuD3UpABtiXipXxRmEBFi400
Xb/wTzjUitedgPxwaQnZujXKVfKMCcPTLtHCjJn7u7ffOZyah30NYyRqArYWglG6oyPrp2WI17u4
HEviHECSZpmxy25yQim8XwrwfGyQBX7CkBWQ0myMF7x1Hd5gmUT+fakcsFfijVRct59Zc/lmwNEG
SuH5Egzw597oTKZfRfvrgYbxLdcM6qrXlBqg8VjAraz5IlJ7gXVvSaLF72h4xFzLsmRmjqVT4L8O
ljrdZzrkd3AhFmTtQx7OWuUOPTPHwmEi1fkZascXEEKHo6S6Xrmfrk/Ox2dqLv6gA06Z8mMTIeWM
tJuLcqdc/DI9uV4bOd55Rslax00PiZGNiIUc0ZqB+9zslb7/2VNKFvMs5R1csHgkOQB4YRTuCuXE
xXG/+V1CCsqn07Rns+LAKmI2218XK9pTXYPT1Cq1bTARSDIfbSr7Tq316gGiMul19mCqEcnxtLJC
iM0Fae+9MaagUSoKQC9j5yvIcAAiYB5T4VOX9LrrUxecs5tIRSVPAJEEv2LD8xn1RvpeRE6Qm6w0
nu9n6OLX/0gPA1p1VNQ7mO68XhZy70UfDId8IewzEwJwkkgtWUGpVt6L7/oml1TQHttP1qbExTyl
qrYqQlGGDCGw+sBdUFi4y7EZ6YGtIYhX1AnZfUAgGnxKlLE0VHYgaM3RuBoltnlQH107Mp0rTQPR
nFE9/5JpdpLgmuLFwbDkA0OebcHl758FzmydoKXOUmskuh3rCdniu4kM6VJdvbYJb5+w7tt4+kPo
kZIiXl6urzMi8WrxDaNKNNbJfQVEHmm69E9YVSFlXBR0RnGSWYnxG+4EmVBJtFOgPqXSjP+MLIhZ
g5xDLsQ3geDdVbapG6l/dl212WAS6lszMdzrq0ju8mkBQ0GrZz+Nxeq1LTJt/kjBoUXR0drgOIoy
uay+6s72kh2scTAfL6Cve8ZZF8TOFjRJn42J6jKZOSVufLTJlC1Z5NAT0leQ6qGyD+YDJsV/CCfy
WSxfQ+SrZLoLegSuvbsIQQYPiMxjKjZGbMfZDc2JJ+Fg/48DlbekXaOxI5oPMv2XlX5pVe86cVEU
VD8j2Zq+9SiMLVO2/yD/FHKPWvlXVO+M/YfTgVyVrId7Ds54n/f7pIP55qtBFrHaFXlIbFP+ky84
6IOmPBmctLbwAZVyuDeJ2y9vY5C9CegvE3u/00bNlCtu3RYuhglPrDhMlV+LC8dsQ4WUFchvMvfX
pWJ5AFCbGAQpQD+FmBHseS6KwVPJp8K/rSTkAdNnSiXfRW283FEf4WJpAxn/1c2V8NWkdxR5BGCZ
jv7fHUof5MPJdLwoHDQvUaTcaaT5cd+GsDvoTAjTtuLG5tIwtz48N2mK2GBpOV71gHigGC9M/EaF
EF6PaqfbsmCanJBLQIIOBOhGJx95tNxpd7Qp53g/Er/bpKJGIdjYjP9003pTX1wDc/nkz52Q05po
JA4mc/yaRvUpbak2J0VgAT8druvi22BsAL8DSGU2QQ/+Bp2qMbe0lMe/4j1dNuF92buYTJZyCMMp
AIMRE8v1jxnoK1WeBBbq+MFtFFZwhkoa0GRVvsxJafoJRkIaFeHT6WPdNvLir/7B04+B8cN09yVN
pPbHtNdNucg5akwf3HGHguovCu79L6KpILBZFChbtLzMF/GedYLFPqRAWruRxUGgFpofLSb1nt8m
UZTwcxfwGht53x+i1Me/fc33jywuLF7COWBathTQw0u5KZCTNz8iTPB8NFL6YakQ8SECDljKdBkl
xEA/C/0WFyZF3ffxTujM+/IgFn6iHTFjHdLSp9hN86zYYWywSU6yzA27cMpjfY1wXaxnJxs6Sj7S
oeOriRJn7MaiErOFM64EDxUiu/KMe1AacH+hBFJGK1rXSSzzyE/4c3pCJvDaHeHUNxf7LKWOAUB2
8npb5eEbbBRV6T9sAwqFx/e6Q/yhK0KuFwT+XQVdhDD1Da81NSHMBgYKDjaMH4Wvk7PYJ3ZU23ms
uN7DBo9mPeOLByz/zOMbpMQVIMxIhlRf9q1Gvf5VULrGiupHdB9N3xnVQt3my/086PgI1MFoZ65y
O4ygNp5rGYtNx5+Unbe8XHdDNsyRudmZcD/UHJESQSzjjL0xfuNfTltvQwCB5kEbesuRmngQ8ZQX
looEGk2veNkxyt7sonxnIjgOH3miYg1fs0rBA1+/XUkm80PhObLqjpDYzGjqyf0zQZCCy0bk51Ed
9b6NOPq7GuSRBHXJxvW0+zuAGx5TPZnqHP/k/AJjsaz+3c6ELxYVA4ZV8E8dTmoqciOhFjh3JnCE
kwwSielTpp/NzgV562+zPDAhr9G5cpQNJKA56XNIazndJZd3vYTS6XVSGF3b5WMMMkqzTaEhiYos
iqfocLBbCtu5qdSETuFSNOSMn6qxW0IoVYHsy7WeHVuMI0U7o/1DQmRol0h2DjZz92wLfdTDCiwE
8fgE6aca3vOcvvxWPYQKYzvDAgsN347U/ZxZIRdJiAayrcgz5gyevMmdOP7+p7BFt5lr0y5SrJSl
HcVHYAv3SD5o1YaO8jSsWCglZe0Hp/aulf94i0wa41MsVeXAx4o66UM00GW30MKRmVWGuqJduecq
IPd+C6Wwb7UkWAYIh549PaHwHkzorKTCrc3dytGD7u+AInuX40jb2c99TqUETGGMyt3EA811CF5G
rCBPwWHNE1gY7quwda8Ef4XxofUkmKj+tlnSfbV42jgIm/clLz8DKUo5b0o9wm9AOlOcAnZZospy
x8XLpfTibmpGEWDyAduMej07l8IshOvLRHW6+IDtJwya26B6rJsmOb92pku4Lr/t2djWxC4dbjre
318xE7spga5Gh0n+BPcTXlrjguB3lQkKxeN8TAjTQLDf5Hkt/yFLLbXzwv1BHYa/5rrgiKTP98Tf
pH4V/rmwcIj6MaLDLT12rTyT7gyAGApndYHvDS/joD0myrSMARy1coRX8jjLA2bIu7vPWxp4u2wH
UggybhBiMYM2SMEpyPp1c4OVHzD4ma8JiA59BXPunIA1pRiPswPt/w3X78RkicoiKAfbJOQDAyme
zu/UH6FqFjdDCk/hctDfAKQMVhCkXQmtvOS+cYB0517vpW+C4cwgBSz20Dhfzg6f7cfEXUj/avpV
LZWMMNqx+Xjv+zM/ETOw+g40jGyYMgJRCeqwde2Y3u11aPaHqRcKo0x2AxEAkPVToU1S5KBbhBZx
l5KMz1S12Hd+pKAy6bBKZYqlpPiRBipwZmAlrkQPDI3XGTLs19nACsHqNIK0sJLlpkrKSWarTk7b
G3qliisJ9Oge2MA58Sf9RoEdHbgTd0w7y+JJt3YsA7CfuWkYGavNa0LvotLIVsHg8FeApgGf7jA4
TebJ1HQ+2hno9Qw/ZiUfda4V4yvS6bt+ZtnzpL2urnVnxKUnbNR8m65rsqCMldq4zd7qR3ICW27y
VmSpr0cKyvbPoYf82ZlcI3ANX8GTPi7p+DVAJTM/4MczsJBLsq81EsIZ8dOz1iA3FaALBcUlPtnL
q36UmlPV4BQQR5JCWHGo/4G60fIYRni3FUwEjonp7Y9NICk+y2MxXTc8MGdQ3Zp/xMwVxaCG48+s
9pQohR5qo7TQPvNpg/dIgZw2TKyRKCXDzAp3PyNMgKb1prifYnOhXT89uf5kn7w8mYlEm2cu1Wft
fI5ecokvl7VkQFT1FHVmcdWsjMzVT/aoIyZ5ezwx77kDC8DbqUz4YFXkUeNz0f28RBXWAl3xfHze
zlGog6l6oR1FTTgU7yb7Bt5IVPI0mMzKWaNiwTFuGn5CCXxbQ3haeY1TiSV5Kv6ztdY0KUrLS/T6
mSpU0bwjjyV4zej98S15UtUUCWG4CJgUzQ43jpcS97XR35SAUVcb665X+fJkqHz4DnFie5puV+54
CJNx5BZRsa1C/6zDppJeB5MB2Rqoe5ip2OkL7rdx2EYPf9C1g8Ha5EF67rRSwsbsvk5AJm2mTwAf
ZdbbX8QM1UJ0TZCO+2W9j6wesH7Z2DIrOX9RdNedI7PeVAUZp1HpTYi9eDh1inbH/Qc5ydojym6V
oZ2FkohbWU7G3en+ApaFh9hgMMZEKKt/IIyU1CNwJGeg0EmvyGkakU8NYntWo2z55/XHswk8jdw1
J+521nq7sHHMD7aqcKMddyjDvYyH8JhkAUHc/MIQI1y7BcbVf39nCe+LZaV4VcLLvBvYoNG7za5p
Lf9SoT4TcEKLuwAhfDpeaTV8YFpx32L/MqMcy6AAjm92GLQUhXibP4tU5fcDS8ippWWCzaleUplh
g3+d8DoPIsusf7SASx01MUC1h+hQSDRYnBPvF7FDMpa5GvaPQZfxx07GPBIMoxw7QCh1eZbNOC7h
6z51zwTW1imk3gIsHattwjRlB2Ehtpar+P+HFO0zLHIwESWxORAL2vf/huNvVercvhocAcuuF4kQ
/y/qKdi8jpuoO23jepU6/D/SOVxmlWkK4wbg043SYObE6syTlzKJsLC2FUiCc8a4VCydaASEWlag
X/+xFvLVbi+ATBDfvv04P4Zm1jfE28jzodfkjDlNGUjEVzEsOyIPcnJBpqJCnXwPWWIB1rIKU6h9
tuyuAAOSQWzr3Kg1CIotrAqwVhVXPqapisxQf801xLJKlWsVj04iXGwicI8WeK5dWFNKQKk+Tuyk
IeAcyN3+fblFbr7XjcoqM+EcdHj8DqMGr9LS/VikOpq5sHTH6o7uTC38hnMp93JNKGulMsSCof/8
8ioL+wNC3wTjER15ekF0cmxy85Lmf/zE5BWak6PT6iXLHdCK6EE+NFCJ1UUNmsIeTbJH+u7dAqOJ
lznyioZyHupSdihrrpz8Gz1Uq09Z2NBbvXk2F0tcXi19yC4SN+oPUCase1G9AHpgoUL8XCw96LD0
IRhqj9xyw2nH2RmyA41fhvKILvLJXrqx3JTCBrH4dsYBKu+ZdORxSl1j5YGOgdsM+o9E20lhVOpV
eVnurTHalhhKOlmNycTt7D88iMcEPE/eNCKWSwDfPkZb5pRJcRInyCM96FmwMrHtltluGbuJ1A/t
o2UUHBWzi5hzMu0WCyUjaZNL6AdsmRAaJYmoUQcvef5NGHImF4PYMWs5EbDI7LZhrxxP8Z4F2Ubs
UEOgYR1g+N9SybMkNCG2gzBTu9QxyG4ThvGaFYIhuKrUHTCfyGTqKxBitR9ejkrJ1eYvJXHxyukH
e3xT8fF0JF8cHtpRFt19ZTG8qi/uKMYIirqBhIRoQC+Cu31Z1LGVyqNIumm1lArSpVziLqaVNmf6
AFrPKMtM8ARW4MVGQsHX9FCyBkBbHYaEQpFOEySaGRT4J0idm4hNBh6udquP1Fsx+Ry+912TrMuF
1WzCyUBxvAPgLKXV1+xy1NhneKMkqhZys1sGnfARts7O0vmHCX9D1SLeyETzF85zP/9GLMCKIgY9
tc9YOKq/YJ5X3UTtMKUua2nASj0frcy6XUiGms1OXpQWYsm0MUU1CJiTvhflIapvmyGFG+PLVnKu
Xo1Ih8FxZWikSpsno7m6WOG6Ay6XZpRfVaXmFgS9BXkLHEjC0qQSuQjuRAUGpvdcIYeRx+8zhIrm
rbe4E5iH+xWWVuOgEH44iWsCNrT6CiqdjDSyJxuXIQfeFXABwcKc8pTu89T09eYdtr/zISHVNdZ9
kT3GsC45pii/H6wXqB93QQ8xUoR6IZGzgd8/iVBnoedOCXmMXcJHK02cLCWg92XXhp461ikQcL0O
tucpAQNzzNVak+GbYKYDXXkdwbeBBJqK8v6mHX8qtfjQdKkHJ9UGAT9EdSTNmZgclE3xJfX9hAct
nam3M2FHT6xf2jhX92iOBiURIvGyB5yVyRQvbMkiSqmPhO0TQdvbp2r5BBOXflGsN+HFrYO24zNN
WX7UPgBryIfH26dutWipGmOUCQmALL6A467D9i1QDeL1VL33rt8wSVduwOx0qg+ywqawbYjNH9EV
u+OkycSMoGtnMFzEhgjTigWDffxQLTXVV8Ca9BuNDunmezuctm3n7LMe7b62IokvxNaT9LdO83R8
2ZhMFbdxqEjMWtuvH//GcOmZBf9QLmK82qB/pBSp/dT/XFwjzbxAkgrCQu3RrfkXm8GgKPQQvTLt
ZTmm3w+zNK3exKBQKKuFS9fXJ7IDIoMJZQIyvUhTzCnIpCRTrjczlZninbz83+YzwTeSEEkWFpdN
fJLGrrbT0AoumEM7XEVdp+xe06+t+KN/kTuLxciHpAYwoF8WCB/rUgGWAvvHgD71jIYhcsJm80GL
CGf60gc3ZI69vZKtT/EdqcMYf7JcfLq0txWbb3KP5uxZsv4kfYCCZoYZrFC5ecARE1GGINAGHbBp
gVvWkoHpGpQouo2RVwY/lKK0JDddogxGbAriYyEE7nqxQIs344qlJxWalmP/FJhejfWfDpPfW7ff
oQ9iMwZRPe+MzgaeN6A4Xw/A0gw96lM0+LWnXCwyi0tWH3iMmtTDyhRVMbHJjDIKZrrZCqW/Bndn
zrrfF9vqaQkCB9Loe21dwhMR8JBavbz6pHmWEPzZFL5YsjkvjHPkX8Sd+70elbocY+SM1lZ+hxjy
4w2opB7aQtmNc7GStAO2wwkwKl6Nfcw75lc9AyWDj1QwOSx3oQwFISFonlp4wYeHAo/Aj24zKe1g
dCW3NOZMKrUIaGwZuf12hT0TJ9TUdJ01Znx+AH71OQPgAn6t2Vfy9YH3qd35C0+2fRzdKSJ8tm2H
vFGnhxeLEV9DSQO0HlCGTdAxBPJAvdYUSDRjMpDHuGz2MJXedpWZhkIJH836eUGbPV2KfZ5npE2b
UfrcmBKrPaowYZCzQ11ZW9MMJfAAhCkdwtDzxeXY198fF9GOymTSOzrLufgJl5A9T7JEXAp7n0qr
eSbN2LP4D5XDGhx3JgRN5DwM9bOGlQZMzgSPytLJnCuETgBJZ/mmAT7S26iY8rVseEDgc+TvzWum
5VON8vAvqaCsksXAbMna3WbiM19CXI6AdLCtdqdB2DHXI1z8AJ/vP4lPUGORBYAw+9pthohFDyZO
iE7cY7UDf/xA/Rrc0zppbGjNC9fyXQZkFn4s2I6z3b04tvrmIUK/yZSs9S6ZMZL1xdAvfo1Apfz3
X+8z/JmrG/zKVhtoUp1F2hYdH8tjBhFi1mnnihq/hCjtUg8wXJJtV0IGqtxLrcVMwuk3kKb9cOkj
5doA4skAa/YjJc40QA9yP/C7R3VlEzQRu7i0z6agJONdY7Wg9Uwxb0yxGMQtUPVKYJOwC/lrwT2L
ZxpgzqMtyEIxiGkFOquC8gs4BcXthv+ElwlM0XDg5XCewxeJolfGHHFacqRW5sDRzbcfu9IJzySL
Y6FF3ORCpw/MJ6PuWUyJqLWxSIimFTWuFB1fhPlny2n6sH0W2WKnmUk/SiB+9lT4Hy+93Knnrr1C
iBEoli5tBMnScWq8tA7k8WhxaY1Wy57s0crP6+an9OHLh+Tq1Dci6RYe2lv58BOXa5iWosvChscb
JAnj+cOVHSG49au8S++y14uP/r5w3jiZnD1xglSAHSBLHFQ2XJAhYwrjhfqB8fAbC5cTIeO3mdHU
yfCZfmnZI1cR31sTUZj6YiO3WjnTOUt3synzjr7fT08BsC3msMTn0f8Iil1YJ5efi4vOfOhQkCNx
MwUlymNiW7+l5r4oIA/swoBVdW8iTKaZHn/m2Jt7k30sqYAQUMuzEeKqqZPu/KwaaJhvolzuXGwm
Cdxw6xcjVdv9SPReYt16EJOKoQr1NWVXVwqpkJUlc5e4DD5gbwSN0QWhkplsn5srqHHnpw/1+70h
L+qrXA9jUti2N4cAXc7183UfOGKPEVWrVx2PfGOWCSMR0duuYbABuuEAg2XVI4DhE+XJtAiPFKv0
g+LOovqj0QFM1dRuvOrxifcfiHgVYUJ7mrXY8auv5U2jod84L4NfL0K4jaB/in/I24MqOC54gz2H
Pprc+v84npUsvWHxZYF8vttnjFfGdaiEnAuBHm3OeLiFj5rBvCJ2y5NGP/qkaA5DldqNvR/cDYgN
bfEXoNo8oeCXjuDp3biLd5S3vPOsp09hvqKzsyCTfLzfmwsM2LwWuuJQvNHbACjV9nK4hp0pNQCj
qlvMdwkrebKvQRqgmiIgFFjwhMLhfHphATbvmK/hkAjRQpn+ZGmoVtXFy2E8weKvdP6Ua+Au/a7R
S5ClqufiGs5dRB14DpwYXJ9hZpzfPhqvmM511R7M2a2C5fKuVXUEr4hTg7FgeIHB0dHhw363kuq1
jOdy9HpJr9dgnP69EIqX+ycUGuJ9hGCPB2dMgwoE0u4YUSHJDlVVQHfkuv0Shbra7zU8X45c2ADd
/uA5ayqz3SYI2i7nXf2SBMjVxSt0gUCxqmgghcYa05/EtWXjNu9Z9/wSZiCHahiXHmQTU7zTL3Cs
uzVlD+wVfsj3JgsZy7av2DTSrTguhO5ktpQN0Aw13rJKYu8RDm3jox6ORiosgxCkV9r9tDaAWmnZ
oSNNAxamgE/5aYYukYszUjet5FEkYdAaowXdlPJfBQk3TrDLkq7AqcrDcPhtGA8KKHMf8NQxDk5q
nLCh/p7654Coh/cd8h0atWwpZgdRZeS1Cr7/fODArc/yA4nrCJxO9xNXefZMRzFy1S9iFcQA1EXi
pc7kvdBNAYo1Oq3D4bUriheubaJ7D12jqJOIGKdshBlOsLbYqE2Y16EJc/NJADhyQQuREes6oLaC
/D0GdWrdz9YIxF7dmkxaZqO+dEXrZNaOMuLcSq2uhqdKeFnPddPenvBDYlrRhZXQ+IKcKTlghyZQ
chGjYb6WyiCZGrO2XGFmaZ0PobMA2ENkPEiI+eQYgKKIgcg7rG3rGJyJVL6fZgrZK11bhmeR8mWe
YcZDiDGOI4MHRdraFIPHBk2DA6P/194OFgOye9U7eRjHeovYYcINYI5xa7Xuw86xvR3k9zLANDey
lDHEDaaNxIy0U/mVPMR9eeIEWNGeR+SSwcfA9D59Y/4i/+t0K/GNwdduXhHJEqWBj58mOJSLtpZY
I/mHr5BBWvfe8MWhWMEHq/DfZWmYtwIwWhMaKVznNS8FRloAYg/Ep2aQEfkvv1WjW2H5kR/fAC3b
r8Oz9SbzEgY9VPLceGBb2vZ5uZq1KoJQhkFABsG0Yc87gS2N/PhJITzguX+/gQ5K9u7ScPDbIfAf
L3HDoY4yYrZ0XId7vbhgMP6gNREDgBbKppJuSXhdLcppuyowZ9a37akZ3NHwqD29xobGzZ0Ugt9s
yjtp/LaHvxX6FgOMIbcA4a/4CGsAay+k4Io6yQKTFjLoy2x8ynfa5jJBR5eSBDf5R87oJfo3hSW4
vbJVUB/xNlJBwZqAT/d95uJ8YB1519teD1bVlAKkQoEWCjSBLidVE20IBhKwvGaS317210uIaiQh
SOC5Byv25mtKqzk6xs9AG1gUNtYojn9YxeNI5/RhFMDd1YSPRkYNdtCAF8Rcx6+SWv0su1fXupyh
zDUCeggrDatTGrFpw6/gu4+tdoIMX3T0jH+5R1oEuijRTcsuO5lOHBqD94iDUDDerB9oUCaIWQxt
slve8RmQqtf6n1sySFH00PPWWdm/v26v0WPnp/ru0hC7jld0+16RwSJAIjS0Dijp7U8emqi6BBxo
uxGcOpWBkIBTt+DdZuQIqF6yJx7N8KYHAJS1kX7qwGAJwT7wfmF935pTNKW5dUELfmZfgoUNFQRz
bz7B7FN4AhHC1ALTfwa8GHDaVU40QSXIoqFJl10YjY2YeSNWUNAqLCzR3Kym/ZhSTEfrqHJ3e5iW
jEosnT6oHr5j8IQHBVkBTgNmqevVm1U1tu1g5RPeijvFiB6gG9Wm2XbFdHtkXw5hzM1ROtkmwhdO
/xXL9CLjceWoC8ETAFLE1H2JdjY/NcWHmEtiCzYIByKH9vS3w2sT7Va47rBlmwg3ycoMVbCy6LxU
T5mkw90KSssAXe02IcdWHWhxb511dKgktruQrM5neNzMqgW2wz0OwmoLyUBgIo7ELioxWOr4hFtL
o2WmvD+vh2ZjA4WHW2UtPT/oJB9UqHbziJr/SFFjGd1jm9LCCEpgedx2zz3CihWhRHAk8PZPBzNj
KYMpRYRutdBzJMOnKSj2WUq5dNVgwRPAru7jzgBCvxB+C0rx4CSKmYdV1yNzg5cQUhCoylsHpdAD
6NAoKnUu9rJJszP2SRjIvaIykkHR9suz83EmSrLGuIb0jDfowTNxFer0NC2pSl4J9/UuXWmwEJYq
DMqrLIN87Up2NbRdcSw1mImptbYXaH/XjvUSpOY7XnM8uVeM4RAUCiiZ5oYApsAbac3plGnVa7Gr
yLBK8Y5Bj5Nd8Yukso+y8GJcnGSTlEfGML3kcacZUvgk2EonI6Ck4R1ssY/3Dc7ikUC7ZFOrOZnt
BGwpQDUTnDu/dyKEn5JCZ1ttYkGRWYcBcSgOmODXxfSshLLGSHpFQMxRhPHDv2H6ijRBD5DCKB9S
LtCagJ6Sj8nLMXGSh+CRbaFi8h6UYxsCTf4aVKUVzuT6YZKpiW1ueeGV5Bzyd2oNmfromFEy2qFq
J+dOa+QFCzKpf9RFufA1lB4IwdMsTtXIr9ShIQNoO+wDwANZbnG0hhq0FvnRIIO+aTn8l4pAG8c7
7sKDOwdaPBPjv7YQX7kc67ItmZ/9z5H68KEkxxk7EEv39x/eVde9dilLkHh5b44aMTjemIA7bwOk
jq5HpkYaESguYxglZDKcNCBUO3vysqQFt8gVwp6H9nrMti+d9DJcDNCbyk2vgzGDba6D927KMDK+
uUpQNuo14OYvdAxX6HU2EhogXfelxlnSE9/jovvMs3hkIEzvblf27hMDZSqv+8i93EoyjA1gIvZ0
tWEkudXxhTGazxd0GowktUZWx4HXzgbJzbePb+wuO1wvpLe1OfktuGXej16TzZLvt2micKZmOmc7
AoKmJyNozgYggmVfO0aZcI6Wc0WcyNl3+MtvjZstL10x1tDuVGi2LdMGSoErvNKGZgGfD1o3xjxy
r4mknMXJGK1Rw7k2IRKv4B83tioIztLY/4PVs40bpdecwiRS4NeJhmk6qFi1w7DIqDWqN64if+YQ
yX98WLImJH7QTMJ/gpgH91WeTwRtFlLSO/l2fLsoXTrOWojAfOFsLffUWhomK+8skNZMZ4t0W3mh
qJt5aheDb8yn8DV4JQmRirbFoQphZKa23nFrVULSR8K1ykuy/j40SaRNic7css7htrL56Nu9RzST
mHdEE2kPvXT9kHeX94Lr8g3CNDJJkF3BF7ZG6OaU3KHc+SVTto23+O6tIApat2hvy1HQeNWtmsXQ
OD0Bn1QE45ZKEvKt73Qj1xrWZBdoqqdyiN1hk3BOJ16AkkD/wOlLdR99q4vAguTo/fLHgBIcvZSI
oR53+C6rjcIBELx3aLMz7F57PuzF8XGhuDKA5bOrApX/wVHVDRZn1rrKhTxNXs1VAFEaG4OvRLgQ
vXeh1v5NYE5pV+94cgJqhl61LYWGLerAwZrQTMYJ/t3mJuQL9DBunUcBpXu8QxgKn6cU2QL92LkT
63jDvx7s+7siRvniOHAHZ1v4PSsqRJWnBbpApsGxEv9nj1eDgb62rKLM0CV8X0O+Za8MIDHxIFWa
JRSiU7QKgAWH/7eKh2VXZroPPsOkfh8nR/nDINH9o3PJ96ClNuaHRCvHEuG4PJR44mF7ay8v5ZQQ
Ca6Dt0zdg/I2ZKcp5p/PijhWZqOUbVhvr0yL/VM9LYJeIxVz5SI6xMWpABlh73fOLjVR17ksJTG8
8gSvJf5ystLJ+JwpbQg7T85a1Kpxp14Z9JG1UMseaivoqIt5wucdfxn9fC/HBDALUMCS7o/34xXY
ngSdQ2BB85DWXgSZ/AHti0eaDHD6Y80guOKLYrVVUcWUwxVcQ3FclS4XzWvvT3SmXehh+4Ddd2Kk
PSZZucYdPWc4SbU9W6M/+R5grf3BCip90zcqQUdd0VSas1BPZuoixOJviLlUdJ2jTNaSISfZb0tn
qqkeQ3EOgC6jd+kNtsLkvGQBo/RWQ0kw+yWaf/+XsPOZLDhP2/2QD+aeq3czDU30y5nAvkTy/tNm
XvC6gmTFrxjUkKn83FvTz/R9O0kleql/0gJqJoNAMw0IC49LKZg+sRIskdiOxsQtd1ciGDxmphbR
8aJCXNFnKoNlNYNQ9dtmQ8UfmVLy6Hiz2KR+QiX25tv0HgdlBDBNjyIOZrzWip6f8O3dRrtLRn+q
uj73sfYW1Y/zuTJZlwbfMNHMOyV5M8TvUFC8haSexiec271oH2i/9zl5+Xl14mqgDxRvHVIENpXg
N/TSxfg3QyGmbNMZIUFwPayDG9CnrBPM82dvktl0ESauTGbLU+vEtFO3kNKUYd0add9eLHdmICY9
W+uHGWxJ8AmTtKMUzSsH2iNVDScq8hTJWBj1mewRgFjP9gMaQnancmOBJHAw+hsXr1KJZAaTt4Sj
1QOFl9k2iAaHdLfJTiOfkF/dtqubm23Bbngl8Puh2dkhAqwKUd1hk+qgGD3Zd/g8sFH56nS7keL2
eMzWrJHBfKqTN1eAqP/QPPEd4G2dwEFREV43hlVcwd6wqWeNVP4yXPggK3W+fTCYEH1reChmT94v
g4ezgJ0V6WGmPcbKns7H3G4GyYTr6eVHSsq4/ZoZ705rBcMgim5bpktrsBDI0G2LisGzudjhJ+o2
vhoWycTkZ/lw1SpgUc5fXl82KgsPlnv5RBBFVjwAUiMq8sn0n2RKBVCVcStn+Kwmf4QAlMqEOmX0
uFTtl6ju1qhrMEdIEUvf1BURaMTc/54b+lpz/9d1Rckqyz8vW1sBDIwvSqhgfaPBWweGKzvwfyUm
9gUtrkxMowABhbTtSX3uN7JTSt64vL7QqNCpZnHbuKoe0ZB1dWMGNuXg6tP9KEG8Ezh/rAL/e73i
D4gODOXouauGslwwH9mXu0QHaKYx/TOdAdbyierWmSmDihxkvHeneI2d5LLFWgaisTcld9sKNi8f
pCBqR8JPkmm+FVNW+PxOWyZjxekXd5q3LzYWT1uV7+9+yufZmw3pG33+712meRyX09k05jC5gxLa
NRHOa0T2mT1a1+yOZmkcEQ1072s2R/geW1vqJJ2lD2PIl4BAAaREANGZwSRgl18j6yKFdPkKQCaH
8OUdlBoJ1TKHfW29dftqeP9N9FkM0geQzMtNt9vvb1kF4zUK3BjLppFZR8I33KSAbe9fTihWpAv2
ns742zkJ9oCF6kZe8sQohLjZXYrOghrTEIzJv+WyLfssjZB6ovNVQHjRE0kTJD0WReptQjBL+r+z
i1/hJfRKcikw14ewe1Num7v/03bbntIutXhYH/6+PY0D94vb178tCuGHPnnfjTwUSunsGhTcYOKC
X4rz9ZXV8N0ocapltem4gJRvY46NkXObD99fy0g4g4yyLrhtwKUGGITR/l//oPJfNcgdhaILmRBa
qlzDUkO6NJuu6HUpX2419r6b2X/UWQSkqQJDV5KsJMCWU/jU594NP0fY0bRWLyVmcUStXRRHgzPa
tC9Wd1Ae0Z80+N/MchNs49RJH5jhjTpNk6WtdEGMS2bDT4geUcgR431SEadaSgBN3QoO6/eHRD6Z
HS6qzaQm8RgcsG3OwzjsV53fKsCecTHVQlIYhhohIHQ8Uvg5dR6heXcTagxPsnEBFsnUNXAv7iMX
frp9MiSD8UVfNaGK0oIwaWe9GeZo7m5bmx0acnWgUExOy8TD1Ez/A2Zh6SogQmxJWmVU6Tuy6kql
8NuGomJjo+meO4TpuXJl4zyxxKzrfPZrSAbnh25ehtL8w7EDwW5pNCRk6GqvZ321OhjOnuAhROS+
8OZ21T2Pz7heuB7f2tpUHfT0wIKNmSPQZKShYNV/GkDLCQs1DixxQHy/BHXtK2hGr9h979dDAieC
gJ4msEwjCrMc0LwL4haEBKxb/f8B5F0MSRHtg2j8rGAqaa5vJ0di1A38LIfjBmRCbxXW4BKLPanm
crTM1YaZfVQiihrM+Gzyqg8pdMsjkw0pAW9GHvHrvsn9tv3GSwsETnDpeB6wntxXUkxWxS5oVbPB
V1loDppmQRlvm9UWO+8BwGlVSZBpNL/QTQ2T20d4AY9leDusuB9sQ6mnnk5Xig1tA6icXgQsHX48
GjBSJiSD74ZUaD0TY4nH7JbQVciYkwnVoo0/8wxKDF2zPgFYe6zOjI3ojI7K+LIVAiu7IW35lCdc
vLWJ+6hZnqZt0V6qM6XbMezcGehKrFnQ1p5NYRvZQwYOtYOXd5m6htpVocwhnzr/E5DupcPmUtI6
KSZA1taXZFHdQYu+IMdW6kPmEz5o+DlO8n3c60rmHBcLxgwKgsFplvYCE7nUejzHvh6uZDAO2kAB
+dt/+Udlv82wsRvTg9miljooCO/eazbLWi4lTr3E2pJkEse984drXKLYAma/PXc7kdRnjFWbMp/z
tBfXhviou4Cj3qfZJxvzhirnK/ziEAg+BOJ3da/+lX35Uo08giU3icQHDgjqaCjDjozckze80nhe
URTue+3er/z0HP2cLgqY3KuHD8U/FT2FIKk5pu3Bn4PT8qMb8CDYqDhTnJRSRVSRwpLdbm26V0hw
lFuWN2jMws1TTyDhRHkxPT/cwh5zcFWEIjQ4McEorDMG6IG0VZ9umZdsMWAArUEKgCW3GQH8U31p
pSUC6QczFC5Z0kSbf4n7KM8kqTz9cO3x0c6mfhQqDDWJ3nT2vgKI1OdH5ZYY+ib8Aj+WbVVJHg+E
iMTRou3ZTqSbxzsQH4Tj5bj4ybOHBRQKj1BalPjjOe14Ercif1rNfet/dI1kX+6rUogDP5j8ZkC0
lkVs/j9D4W/DtFO6R5ypCIUSTTfu4Kqaldp7BI0EYtCCCHwyPvzrXHilpR4Uq6o7oSAlo8W2/Zpx
GkoCSjiLS2br9N3J+tKAAZlaBy0xqsfyJVyFhnJNoSXR33ynrvEoMmCvwCo7jlwiSL+cvgUBbzbp
JT/DwB5ApmV3gmu6s6rCsUtAAQ+SrdLzKXblrWlcM0ptdrQJUxl82aR2H/FwaKEObMfLPSMxUEMW
hJXc+nAeRgQNhB7QJpzJ4+QfiNcfvQnNvMMJoB8l286y+27dvVNx0Tj64m3GZB7E9yxF+g==
`protect end_protected
