`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
GhoA+/icbT0Ipp1bgfbThTLjt2I2k6V892hq70m+0koChAh17VFgHCtwKFaBlrgb4ja9gRHntw6Q
TJW4qKuhWA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZNvGNxdfqWAbVYNln/3iD5E8MA46pUpubTf4/wcfjvusiO5io725OqavcDDxVEm4FDdpLJD6cDWq
K6q7CdoEP1htzw7kaJoztgODlp/FQKwVwFtDht6psmvhoJQM4vm1qI3Rzh6nOaMxeY8krE9V0fUQ
qcPNdfwuFW8kvR3wLFE=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Eg/+bCPqrNn1FpQ/idY63ixAbvltPNqOcwbiLnQKTdVtFeKc9Mp6THHzJFYeIMwQnoLLnwD8boZM
bLNF6yfgunAGECNC+NrrTTFh5b+37nhWMDaoaaRyzcbn2zjFMljb3IaRvtvUKcL384fqXX1rsKM8
aVSoq5MoZ/rabnB1u7UIf+dwb3SZ76q2laOybyoEKOZytaohnxJWXDs4mmn8U/Sj+LvcNPaeU0VO
w2hUqUcYdBqHrWHPDi5OI6d5zRtjlK+i9RgcZr9r1NfJ81Q7yM9xjWO1nArR/ZO81qIiHnYq5Yfq
9Uffzaimni3W07vbEW8Dna7idH/FApfMBEnWFA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EGH1DZdxFr2lEbqtw3qS/IMoOFKsFmRhrTzrxKYfOYXrjIq7/vAwZoCAmQWpp8a9xvhKR+DnGf0g
4X5CSkH8NIUBrSnfZAWQZHDXlNVhR92lxfsu3qMauLIZZzPQfogE2th0B39lbU8vk+Y5yRbFmywj
ZfAPKuB+DyPP6zbc8HE=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rwDgPcXSPMkww7qDPfm0SUJDvmV2Y1Mf9xKOPBS2f/ZqROQ30YnTgCtCePhqBy8qkMT0SPyAW+GC
eVKxJtWVu9TdBObhIxTYga5sLxazigFksGLQPrK6O/53ABhyjGmg+6F7E40pKqOwtZzbXSy6W5Ha
QAvj3KLASvT7kkoBe5Uq/NKMuS0mCJqoAcnq20FJsDzd7JqkqAu1V38p9YdHEY3Ws7dXqILFKhL4
KJxauMaAi+zHIvslEnQ18XdH7LGVmGfQjFKE9UlGfXYqCwOI4ptaB0dUKUOUSjZmdbTQUSQyD0sY
BPWErql0iqkEt2hE6FVByB+lDGxTTRtBGAuCSw==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SvzBe4uqBf1Op2K0cnCIMKZHuDYvseQZlDoUAZm3B0vqnXskFzPjZc8z/K35LkgyMyP6rHDB6aHz
oAe5CuPT6e90oh+KkrPSoGv3oWDtFHqQ2vzgXzWSwzHvA9JdLY0WECkURxJ/WvvcQ2FEof/8mtpe
RHeHlScdIwS9N1BWSNsbkdGFiex8P7qCU3hbjN/Qj1sRx+x3OJDxGjtRsO2wpJ80f6w961nEO0hz
LVbajdAYx19shShiX5Ku09QgFbr/V4O2uZHn+iM6ufLM/dlPDW3J0ktz/l1ElcJFlzOV8vb0msX6
4oC5ZUphBy4apJrwbL1tIQdDVOD9juS/8NQ9Iw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 119648)
`protect data_block
lIJx2V4eCqBNB4utX9Tb//1kEv9BtS0AU5WsFuA8Pfb3q4QuXGimIzVWPAyJ5/KF1zq4Cu2IhNmj
65MBW5u1vgTd/4xV106ZIxB8NE9vvv8Vfi4SPIV0SxlzKXSfdewD5ymDJvrkHsf+vnvjcR2QrRNM
0bf8j2XJli8q+UKA7qb/OHEW0dSCww1H83AhVfOH7pA3mKRTXlxcjpExgq/4NuEk4HKpfLrAZ9mV
wimQLM5CUUMEcnINurBT1t9pEtue3FB/gS+o3aCIG80NXInN0/Cy/sR22IyooFC2dMIUS+ikIH+g
iLNB4kBHROdCkj1H8wCxh6Wgy9Cu8sG71hZIzkCtqLx9zrZD9rS+ZNJ+It7hq8/aAh4A/LvVmoi+
vlR94xxz54ksraJVzpG3O7k+52p2psyU6OktLotxnDN9zez9OKl6BPAFKXftXsojbvTuUVASrADS
Cbe7tU7DGDnI3LH1GrOnUiefnR75gNbcG4LWcMaflYjXs3Sjh5DkJ6uLRjukVsG4d/214r/aTQCW
gA63ZkZ4bYkBCfDbvKFhC4/y1hRhjQlhumjt0ggkd6sVP3hGGIDld5Wtfam14twPCun+ylxbnUGQ
N85ScSPzqYtcKwHNsg0zw63yWN7gKp6TdZvOUNqLpZ2qPJypDKpQ69BJyENO6hfyVfScyy5L20ab
3PA1Y95BW1YzB6Kai7b5wL1M+B+br4ThLv8dkhKGdBKOEhjhzHVT2BK83eDSb2IGCUk/RkLBmIhm
gzOxKNwEAyAeOZDfDAVErO2XgVCSL5alfbm0S8Q1fweFPbjVDa2uXOdBLyOpn0EGnJp9xhIkbnL+
kAQWu/UaSO0/PKZzfAqErw5apz5gbXwWWRYxPz0ZQXsTfrFOZIKhQc5g9+a/1BSoShJ5RCNisFas
kubVTH3pt6KmnC26JpD20BuwOa9LFqr4uw2a/4C1xocEgkxnCOYPhKJcXrc6npB22yrXe2XgmA4v
VvSTpXGm72lM+mlSXawDubbSQnd2AS20AXpdLYWfD5CPgS7uxUaVVamDhvuNpJZWvNcW95hSTO/d
/ZmcSwLj6xanMRT8bJ+OG1Gu9c0RN2U7CoYtXm5RkgH1RrfTUrjOw3P1HwYT6jQYj+sAioKasJET
i+xvjbsuGt0S5JSKzAt5Z3dP+F3d+874r/VABpzxDO9YtP3G8nsQW0Dsa6Wb58Nxf1G84pfMqyPa
/+RiF15cAb2gSThMO24OgiFlzppeHJhbS6edAZS/irZsdyfQWXeaZBpuZJ7X0h9GUobfpqGLMvIP
6gBLOyZ79ZhhzgaIurr3TX2fo9O9GxFdhtqsxaepZ91HscJ2bxKN7lBZtrbsh4jyuskqly+Hm1tK
GGt1yuJUOVs/T58oUIRdKwv1pMVXkCm+mgGe8989XXxrVNyqSjfEpooz49txg2e8O7jZmdNIAV+g
NcOVaMNnpBr+3KVEC+lp2pi8HNLJ0Q23AEvM/HrorVL7Dq0Qq0Lamuiz1PnxJ8OcIqCkhHsI9eaf
SXMvfps/vepYLiLYISCPtF87UPzCNRXZUL5DrutNoUpgb49Fhl1i4yjE5/xYh96j4olcR3rtDOU7
8+x31OhOsKpylx1kMAr0Amg6T0fiM/1jOMa614Eu/ZJaOiZt85i2T/zovRdeNjLlIh2lm7aaQ2hG
3iIOZYaQxgZGCXlLxErcWh/XRRe85+G+Xl15foc3nPZ9EOAIbh0LRJhK2QZ95p7Q5uI8SQlgtMg/
cbtIr4sjI28DtYnfPdWY7z29CXMRYq7YkmrlWSaKSE+FkARrgtFU42CP6YLd/376rBHQKPmoXAVy
dzxa5Txk7yV/2QZxiNeBDJgbt519RAgAvT9s/lhzfsyjMPOd0jyI6KunKLol18cj6CE4ykVoWIq4
us5FKGmgnPbKTzey5F88jbKqNs0CKrcUvttsdOPzOQkUaLj2DGQifZEIR3j0jrxtwVtR7NPtdhGA
s6nuxALAYh/mFb+ilzYSrLoe3aJvnoPlwf9wCltrF29vm9Xbcq5H8nxkbXowmFcywCVPRuR2fqfH
7UcAS9OP0z0nbl8TVRoMsKgnswH8OEch9evDCIhvs8SNyPNJ/QZ4mipYXPYUflT3+hyNddTF4u9/
RMLV32hdsLFnLpyisuauObZG+FbSXaycU5FbDQzJxOMwHAoRdoYHtyXd8+r9uQDJtTKaUwEqe4ZZ
33SZfy4lFSMgpKRUC5hw6zF3LAaPenG3Z9+ntSBrovSreSdETwiUTT0B569fuNh89EyFSJda0TJ4
OUsbD7gCy14UZ3NVLwD0t1ZM6q2Fo+RtQ1zAuncV8fKb59w4MkZRjzVp2cqVVG/Fo1jRBFvYkNeq
44sGJkXKb8FtvMc4+0noO48Jd9hKGKtJiqUI18xj2QXnIHarsX/QnvrusTN6gEwcIzs5I81pfDYD
zGbOrERx1AcIOMOKgjsJlBEsQoJlc5qpVz6KZprwgJi9ghA0ix48oKkpSCxBnT1bo/q0vhnIInhX
kS3baunjkhULTKSwqGfuysqdPrUKnsxeli26He0Tb4pDHuHH6DyCA1xcjJRY3iDyaQ4Dcsm0kVMg
JKVwLia2gHl2FZexfu+lZWrGz5vJIn2h1U19/wjy1qyR5lnO1rx5DasHf3+PP09Zw5+91NFoknuk
olarkbDSYHR5wbqJIBmzMkTU4/6oZh7knfW7ebXG5sJHziDwh5y2ba0uzRpJ2xYc2Kw/bIpr4VwE
5M1SMnpSR1mJy6Iq4Ki7v0Aohtk4QWpbErwaHHBlAuzySLkKHmfXtpf+TeJZ7pl6L92pWFJUZLBY
jTc7C4kG8mMaimRjmWqtctzy5VuZeCsBu3gf407UQmKiKmejCL7QFQEvPPbLvI8zn6O6OT5tTHXM
Wn8x5qg2e7/qYAwV9tKAlVSbNGhixccWWqVJ2Pljdopw5FNjJu1Ok8PXI/6l/VmzBRuaT84hDUnT
IWGhUu2akqYqwOsssjNlAOag5cB6yor+tWWyYryMcF9UHdfSR+R0AK7TrwNqoTrXx5mB1L6XTVc8
EvGPDWilXGnDB8ZuYOHJkd02A5ngJtq94c/k49hThHAlUfom1vZj6Q9LQtobTh0hcd+tAwgUHqPn
u8VBS5XNMF3dbwxvjh7ctdX8IoJUkSE+O82aVTtnJoa6wBhYKLhdaax3UCxdVbGg/m8mYDnkgUAt
ypg2SmxE2eoLXRJKugH98Djq/cfnEtKuzHPN0EiwPCL4J+tFIDQw+1V/WIWtA8H6bglL1Ep+5JKT
7gFz4B25f0xqN0HA2qrqo2eQQCLtXYQ0/NdjHotVCg8N2YA9NaAWFgWgS/opgSSAxgOQ7Ng7roc1
Wum1mIndhYn3QiRnW3CMSn/UwS07Xo0xWhze7mrx+Umr2EqSbRsOqN+xDqDDA2iEnwYq0SwV0XAk
oxwT31bbHGNkHPay7CrdIluHVaxbSsTkth8yIetmxz3yD28oOCGI9YyjpD3SQkB0GUtpzQ0lONvs
OpcfxbVsFpUI6vjU0gDEmJUwroULCeCacAiY813PZk6/mfJ60PK7MijefLFqbxaw516FT2WSi3fC
CvYmc+G03AFAxs8sInDS3+8fFjqe/1tEuRCj3gSOo/obJCscwsCirebVGw/qeuAKGz/Fyc83RMXr
xR9VM8UUrpIJr/x+zfzPVrKlkKDysM3sFvlqjZO27Y163rz7vGykwGvmWCWOKin8YQorrHJR8tMM
4GL6zXhdJpZKjqD6STXM3VEFQrSaqaPnrNv7lCk1e4K4ZyxpWwiALyJ3RjZsljJRQWpZKeEO/uJ8
HhhxxClS9Z0cKNrPgDqTmxBXmiDwLMiGDXDHj0aAsucu8Lk5NJLdmNSqMLuUA/V3FvXJwnQzAjku
WX1aRRaXMDlea+JlDzDWF90E2lfViJUBYNjHbZkSoE7qMfYrI5nA/f6RALP36zzzpMh4qoOvF8NW
OjzQnWfaE1NA+6gDgn0ybCIUNofhWvByZa1lV5P3i6m4X4yCJM22e5S33FC5KKkyLKrtfyBpyFF1
Bvb2ukVUE2hTIMf4ZdzfcZxve8ctU621YeEXphFWdGamXvANKlmjuPhYSN/f5fiYvfWcpxXlX2jf
Qof526oKaAteKBodIuduO2kPJiFw+lwV9SfGBpUuisbFfjz+EpovPBQOgrAKVYwSWceXWLuq5sBt
U0HRv/DxYp47mY67Ho0xthF2Plu7J4C2AYFN0Fyhcf14xKZbVFQwLHREARDOSVS1Pol92nV9Jzi1
T7a1mozeY4F3MoVNN+lONCzPFoCBufYaNTdxKCq42/qH6bY9b7d1zOUmo2pG/HeLxM5BfIzfZIZc
+sbzoF8V91wt1pjBBlnPlD9REdgXfISCsvDLsXUlGujLfvuwczn3gZu+QGN6Vj2dEpaEoptRVJrH
dX0LU8Qnzxgza4oA53oKTMpNz1QeJjXPlFAP6Kf/0CONh5/kekUWomQpB6+p8BUK+YYbsBeHRp6D
o/FAIysCYUTZS0EVtMVF4nT+wDsBPEICvJYHibw36IuCZERVxTU8DeDzyzvBIUkJOguSpfplwARd
+eHwsqCJw7k2P3F5gxRwdcy/ipBoq/ig24CnPShzqiEBIvVxLIktNo5ADicywjrAzuba6bN4C4jV
/q+P+i09fHaWQTZRWGFqIQ+TF8ZPRDoFvOqOmDQv5P+lw7GDjkiA0eC9a7wongp8QU/n8Ygi5WJR
eJFkLqAvbJfHXEYfd0TkbJez+peu7j3wXOBk9HsRvYEpzgqd4epOm8oWtGDfQGOCAtkcEj3VzDdb
kCBxxCLEviVLHUi/5LstqBfWkcXIiH5bak5KYK+EZBmSdFjmpSMgdwtW0pDTSqBqgJAjQOWk2wOn
cr3Hdp4GY/xJi0xPdMqC0LrcBZ1wxOGIpT9Gk7dYRfwBwPXn6xzB6WpdKIarKdqcbCiLjYgHhy3B
xfllnboF371tZJrIhajBtIHTaVoM7a0zfWc9KXoJysbaeOdFjUZ7Kg+RFOnYqVm1TtQmhUt0wM5W
fR9+mlvob8b3CGFbNJKFonRfzEf5ninweCnQIYLpNWNDhP3zbor6J3eYmF/wXz5eTFL/6v8TaWtq
yrPsEGQUg1Twij0Hm2sLzIjBJwyaV29zDSyC5CUAd/oosiSKDk2FyzaPyeG1tpnqNJY5yr/ZkYVh
VuA6ttNdYOcL4v3N3oRZukv734GoAk89TUBHXYKjbTdkYjAcFcIsRTLv5Go+2jH2u6Di6aCLZIG6
p7odbFYwqfzgCxKFerwaVnKcSh9zKVGQfZSCiIQxEH1IvsiL0O7/eIgLMwXPm1DaIjac2UsK6GY0
LVx8RW+C7q7C+NRjhv9rarUVqk1mRK5HNuSM668E0ekiaLMOccTPGtRRUA1LiPuKqm/4APnVi+Jz
8Fq/8T8gFtvT3hjvc+diBKmqW4Y3Kqdy8Ya20Wm9FrWP6UD4LUsvqngWvU1nrXaNxv7TjEIUUXjB
EDES5rpPUymOCCnD2H/T9ZD0xs6oAhVQR0k2gbEkgeJ7A4AH3KyTbUO+5LH2uJqnF2NloLDWPcHT
8fTiRprwCq3+W3TWULzmj8CtXqhzHst5WNT77w9QVwE7FLqM06PgjDuM8swKgPzVEUH7zRRGsq2f
YTdJ3Kc4QgDBrIenN66JCNu0sQ5se7ZI+R38xNBAm6985RrZgCS6yHqdStqZlx9IlV5BKNnejfko
nrhD0cfu8R8DyanpHEyffTvLqosoBu7zdh0mWGvc09TK6n2f8PPpAfQ8WFPVi/sCMzX+O1umc65E
VhjEdN8f8uCBa11C4Em1xG4Chy0HuVRUsJNv3xJZobkmDDPPao2G5/D6JGt84djfYETvlOY3v9eV
LCuzTG561AhotCAOA8O1t8tiWBCP8N8Sc5VJ1NcZwRh7FyJjr/GBgitXuKDhe9shaQ2YKHqb3N0j
jPrdXPcGuPful0V0HTbP/O8qhc9PsC8l06FSxjtPWDyazWMx7qPOurwtCCN6D22q9qHjmyASk+SQ
8JIPvoC4bJJMkNk2pw/Rsq+56yliUSBQqAu5uJFSb0Ndsc6y1RXvqdzkqesgHmFFl8V/febCSti2
KOgkTDDUx50Fx6Nq3xwvDmIyUI8E/EeEjd9lDtVy7FNV1nwVP9+dSxofryYUAWnP+wwGpqyAYJK/
SccgPaD/m41BVLSv/mtGRD7luwCarNhWfX/INc+jbpu5fytTTeb+SsZsLvdteGxgJQcOSff1aAUX
MG0vCM2S/RDBtKkDyd2eyD6N1ogzmUo4Y7s54mGG7zVXvkciTP4bvojq3jzxvvkKrSBOLsr386Ed
MjDh2QoLL1TPj4WVuafpdf/P88dUhxYcNgpPtTt4ny1mHL1ohoZ59eaixlX2wHtwr2b0LSV67M3O
V6YglATkknZs90TFeeL1QtCC5PuHcEi5WBUuNaNXTUy+Lo5lUxQ6A1hfoEfImscEOJ5f7nG8kgtq
vzdAruI/bHwgl5WhD1WAXIjhGvV634qWNLy+YfYAWvJiTlTBLDCezSxT4rN7K4JwMQotnHvtyOO5
h2X9ccLVj9+ggycr2faCtq/tloNUWbBqrTxh0tLM+7L7NZ3mQ8HpRpX9JFUi4QZKpFnEmoANGyrR
oLMoRq9ueO1WbFT6d7nEHUBa5Wb2/F0n0O3w2/EQKko1ZwdSZcfHPBgiwK7sg+DfUaR8vbpNboYS
dH8PDsPUE3VmkjlECzbL99kgQMz3L7YBJ5QQQuOeBw9ZmjVCrC8fqPCew84ELKpMQIpxuAeRsbxM
y7Th5XhONrCe8OTZ9wz0+ic7JAA+ACvTHf0WfVJmAc2F9KpHcFLFxdvO4/wlJ5BF6NWcwEXp3Vtw
TZUkc1iRn4Hs52NsSbAZJ5Wf+El9kSK0gvPnQex5LLFXtdgbOhaX7I0DpEaMCTfITOz4nBfHikbz
yXyuT0mJH1tu0g2e18TNe8NyXspg7swV+5ujr1IhuLPMOlowMcXwySrBF5cmuwIJqUu5OlyKa5t+
Jq+QLVZ+CEe49gzRbQHHZOyVEKBrOZs0/1PZINMM72XHEUixR5ORZS2JuzYMJEGlkKFnOo4xpbYp
Ldh204HwugxlYUZ4X5YgBtenTP7o9UJF8KEygTPcXqgZTBmmBqgzBbDnxH1ItQhFnnfaNPyLQzqg
HgfMjE0FBLBdKulzTkmJD+Vt2yrWdHdFtcbe9fjeZ9RpjfXjG2Y4BnnArq7zlgcYdsbIuh7O9CvA
Hd0LoBSaI5ApHzR3+eeZcRHowx8idg3dnNJjMs/eP5LB1jAMf10zigz1H4NnNbm+0+tV3Pcub5/+
y1KzumSEmp02rS4Kk6U542Ut8jcVXERAEpe8N3tQy0ezD3tIJKBs7q5iGNBQGQEmCaQZP2IgHGtw
0r6Z/rYNRKZZI8D4eIpJSMNzMaWuQcIBjiYuqzlB0ITbttLtS2k/ScX14pMaW8WRXjDxWxe4dYFx
jgnP6kJV9UhyJb5LhFDr4CHfkvo0209O7snSuiT7Urv7ZXUSMJeLqdN38prOohoB/OKcrsxVncTV
g++yFTQYm8o14BcFJwAz2/K6X1hiUSIGYd6VDD1148sU2UnXybaX5ZLiLczBA+FtkrKNXyKg/iQ2
DF2eiWS6kTCOrmrZg6LIA8lZPrBRGJO8g+QqmZHf8QCsaWvt0k/O5zhT86UnX+H4uR8oEWxFH9jv
AxCQ4D/TIafYmyx5WI8tGB82eqCfaX3fX9M60V+vrFX7t2wXIGDdRWn0pyUtHHdgS1J2Btt9dmJY
xOkk+5IYSZDZ0LaZLQ5nUbmNrsBHSpYtZOCNQbxjnYt8y6whJmxEo2qY1E5HP4ul58TpbejL5/F3
MIiVi/WLq9FB9nijDt+yUBrAkpTnOtI4J2tfJGALIDxAhDX8vEhXUwPVnokOxpWgj5LG7EbLyDcD
8zlbNGfvKX6XH8KUmXVRmvGlwsz7Ir4cBg7IoTQmRXREzDL9I837RGMl3QVCHMxSFJ5AOuv42Bn6
d16ZhZ7TFSu49I06T242oxJoUeu7OCywBUl5BHS9phcMbhpu4cI/iEy58Cdo1mLK9MdUySx5ozLi
QaPoG48rsPWRNnD4rF2j3l3Vqg/Q0rqyjX4SmnqCMF+6cNhcSz0awdlkQB4RxlGJXOQ6Oqcerde7
9fFajgLvXevYx8vfhF3H60wiPYnX79zg0j6yufjty2JUDz040fKvWOKmlcdoJX0NwlEWEdaXfzBC
9Ve6xI1iLpC4ZAYCzZi8yIG/rWLVRm0J38JRRE1OtIIJt9TdQMK2Qwp9J3MPG8OsClEwf9lJPcFE
KKrO7JseoXP2jR9BQtNL6Q5BL8H6LyTAa6KsNRngT0b9TwG8s6cb7blnmV3QCsj9pLlVlC8LFpDf
VQaIKQyQrAG2AE9jqgZskMJtKDotazC9GBXaBQCPmkx3qsN9ApITbrrPoiaO7gqTImDGTS25wxzl
2F/4VOG448UUbyeL7VXcnp0U4ifKwuNudPJ2HuvqXm3d6a7nA4X5i7dVVZRnNTKsl/nIMlZta+Dl
CebSW2CZDGz2Rk8NVdQXf+R0Qr1J4Qw34+gFrKxRY3Nl/V9SZv0MvqPkWE1HPgke/xYtDodOdfBL
pWLMP15Z+3Qgnhr0AvlWaUnLdUxX7fFOOC7v3RgFzQrlG5rPcEAX7TANBRcK4VHZk4VXcMwzBDgJ
EQAXFpg4FQr6RCg3M53PAMRu+DU1D9tf1gw1p4zI4Gc04vH8POmFen4tWNCUz7TEkf9iEZGu5cFk
36y2riTEr9isAIGML+yVcSlE3nJZcPZunXA3SD8Yd8oBQyrwk/Zhz4OBTROliF2oCDHk/uEk7Dqq
rTkzOO1XzvPm/5RuoTNSqp5Lv2EoQxr/NiRDABhdqYVEebSyzmaboQ5blVMpaY5JaZmPvBF6gih8
pUSp943i66E9vHsAsuXbiHQ29koJiKJ1bDao5Y2qFH2konOmtm6qxvBg+6f8GG6mNgWa+Xyl0Ndb
y6TBKaBBTheCL/INaCLMHWK7SHek1Zf82phK8yq0jzUIq6EHu1R7MG0Vu1wx4/DhMCsvvsTeb6SX
GLxrsxQ4+JDWt3sSSbJqiwrk0ixfJWqML2cNBut9gQn0o4+2FIDghXcVD7sGWJyfsirty62aljMZ
ZWaDLu03nr0cVOdXyw4hbS6EouXiPS28F8QLSUSEEgPYWBxZYebBy86Fo3fW0BINn/HLzu4W2biR
Qtcu0lJLGqmMeCDeLdh+s/mG8eQTEqcEoC9c806gwEyi6qJw63njMErGqhYSvbyhwexz5yVzwDix
pBMtxN9H6HQkYfQx+rTDbiV5jLzUFEtu5H4+rckSR91ImIjFPx03aDzVdUuHStKNq8PkZbQ9xfFO
wAKa8P5rRslLEDr6iygzsete5uihlOVU53QOPhqWOaRDdsvvXXJ1srcpuHXHIPAFQ2F7bbA9SS6k
n3PMpTufmoM4h8ox4GQx1sWswf7HYbWzoXdLKiPy3ygVw4W01IMiibk2NiPd4g7WiLmBlAPfuWpd
NUHJdT170P6ZR7lgh5RbXagSMfGbs5570w7HR8QwcSJ6Sk4b1NPqJeAhvhboITIdmeKO4Z7+5/oT
FvYurMuQbC/De7oNxnOUNYETmfyBz+FxffbWALBHcxGZRC6edISjTkXo510yr1HjkSQGceQBthCm
6MPN8nfHgzwdUb9nsEkUQT+CIZhdpv7FFWSu3IwhW799X1e1Kws2WXGy/PuyfBIO+ctp2KMP9Nmt
K7GKphHQOAqbqKRpraZsYELc7b8aH8tdt/RFgWw7rc6Lxe/hXg9o8kVARvccrh+T1qNfGzYmJlmt
T8tFcHP0XcVfVRU/MAUl5LeG50IV7G/gurj5TB6g8U+s1hwiegzYc3Of+xVUEcYjyPE5xAIvtrrc
bL2xvb8AsCX85q0muteRwPct8JEu3K5rH6uhb/HBjcxUYWLAhcfHPMscGeX4Kle8HUMbfQ6vOWLL
FupmDj0g3hXTyfl76TfL1LlOW2hACsDRV87dmufOnRdZEotwACRxqOhgBRJXYkZdDCT96osi3TyV
s808x8Xil65Vb0PlAFcjpNs3QgFv1kgSh/Zw3wVKQ+hx7XfX+aBR4pUN3/4GnVv+EGibsbPnstr/
ceSQ3OUgx4q+01jvpcV4S1VN+4BCw66sG/YMq9Oxqq6qvlxli7PpPI4OEMpR3DgPwrGAIeXTtjrb
iqhQEcIOtPbMKjUPc1Ida6l8rHVB7TEtV20IODSrq2Iv0ECAMf7rI0Heu9ZCbO5EkMdWyJIMc0Mi
qbAVtWg+yOsa22CjMFRV9v4V8H4jSZCRxsDQKazcVX72/EyiKGCI4kq8q0uVlje0QQqOnIJSLuoo
T392q6vQTjkHms+O1K94ewRc6nMBfW+/fZSSv4U/62mOv4cEiLHnazUz4fKsz1hFnbOoFfo2uS+0
mrKTXztg51IxXMQbItEwAItgB5kUfk0P+LH9MrPhmTwcBPNvXr9xXo/gtDAwnxjgoP8CF3MDqI5L
mw4eH3tqqbj+qhE9OmHNZMwDDmmaywSoESXVyLy62yyFcRA7B16ou+JPZQaE8OqBFgCLW8EckFO+
DHq7kbJpsu19WEZmwmxW9dy6Lly4eS8SiRVAHWtskWM/LApbynWmKztOiJwsv1yN1PnSEIl/kz68
b2UltxHDuQyUYd2dY0tHKk2S0lRGGeR0DneZJwD1WGdiOgHMGbdQ0juNI3eRtj6jGgNWNBHqEX+D
YPL3O/bhHe4a5C9m0t7yafS5OIEbLSxu80biYtIK59jIAJ3MY2ZRbvDUyTdhlytWFtuuFd8wCjI9
7NCZse++r8+lgnXlBZloAN6nyCFBrGsCQ0wMFc8+fGqpiAO61PiCoxR7EJ2BDJ1IpUkdYPgQVHpe
Jji8mUVbVfexS3IOZ3RhiTwUzxrlO3Jyx5vb1bsGqMxkoQG1g5uunawS5GPBu5eIGUPsHAGhN9pl
qFTHd3JpTqJ3XWKt9Nar0JchkM+xBu6TfFJX5483WT9kLWQm7pptaOnszL2UJufQaboNkf91DwyZ
9zOf5hr93QtLmJjUv5H2I6quFHx3WjsoVPUt0kLgVxXDzQxx7kM0uOnYLbn/pexDXTck5PyfcbsR
c3+wLqlZJWecL8rEgzSxxB9YZg/furiYb+UzpPBiFsQEaaB6XRiwGWKWhUHrlwlAA2piAISFzkNw
DxupKMB5yc5dL47PXk9WM9pq/4EFuB0fRhQuwuKZ9LCSVrAvdUUNyuOk1sQkXrmRXlNLxtdTaMqn
3WMjo33PzrQjRB7+1xCVrYHyCDKp4C8oXMMACMHMVkGY5rizoixlkVl7xA8VxHuqCZkSUKj/8XAF
kzulf13wiQnPhFRAJjcElNcMGqZwVlWNjCkGDEr7OpTvEyk7lcA8SPoxTfvGj0/985g4T+bmsZkp
5h8o9/j+fRY6CErfk1QOiP09r/lyXdO3s1LNeNpVcxGlcq1p/FoTNiFJJyaKKK86szlIZhvcR9di
P57cdtneiLaFuv8GoZXePeEQEvnV+Mw8Ipra8lcEkvfnXGMI95BlBzuOnJeUohAbugQVXivnXEMJ
+5uus0yxEyob6eDZ9lM+9H+F0jgA7o9f77y1PS54oTgjOKzH3upHbQ6SNE4cW7Lv9lMTvzg4WsoR
MKX2d032BdXP1QAXOy6kD7GoRRE3KHP6fqfBi4I66woIN+ZPdumT/l8AWOf02Yj12zDNSWv9/DrE
Ht1H6sc/9UQx5hNmQtA7grMaxAPABcGG6lNxY+Z9f9vMMGXNVv8zYP09UZRc6RJLgLE//ha46Ym/
CFn1xopqTK6u9GrV4N4Oets0VEClhdSsWM8vzCD4A7CNvyPzl8aMlxDLGpp4zwh32+Wj35QNdFzE
+mHozoCipwzFT6mVIVsqTwVTqLV06yP3TYyyqlIISh5jegKxsA8I04P7RfHxDwRD8ZIrBlVec4Jd
FdLfSoNeTbaY6/+b97FjUXVMJCrB1gfee3XvmI6+kkmIIqxOfpTSdiTdaTDZ2dzh3jhilQPpQeWV
rd0szoGcxlbezqLheAO45b/khiCPsPABGGrHom5y9KFn+M5tE78sWqukP5FJotbKDORlr7nv1Vk5
UUFDuHf14aufJqIw7NjlKGfXVMu3mutrIdwlk49XoXUw2llVFsFnTz5kN7fmWirJah+mza7UTJ9o
Lagu5hVUMojL73g/nsVQGSkC7MBh7OBeiq1ShiQn7cqfcF1t6p128cEbSoMU55G6dG+oMDHbJhNm
iL5ecGd51vQY3QTPS3gHVN4eaDJbw3x/yj549UmBV9GuMKf5CfWPDPAYyuiruPwP4ZWeu1Lc4Hmp
kVI2Jk0dckhnnI75C/44Pn0gGBM2sbJzb8jQ9rVWRyejItML+n1gSaP5i+kW2lZJ+Yq+gWu8/6kq
L8laBdq7jnzPnVNg8t0UhIz9iHIzU+hYrkyy6VkO5ZRfCiwrWLijpd7G0DL5bJEP2T3EhfhhgJC6
zQrZQgWi0Ri9sJlt/cSD1c5l8r990Npa8oWmzjSO2b3bR4X8LoB1DvaCSIaoaSXs6Gd3BYju4x28
4ujYq6wbAU8gLvgfaDKEpPkgoVLtIeGrBRorZEAu/b6UgHgwZ8EwyndySXx6yHg7tDhKsjSWo41U
LRaZywRxX85pl7r+P16t/B2x8omgvRBoT2KQ4ve7szZclCImsGztOF4hpZ9I492jRtl7iffPh0bB
2L5kMTKLG78CqgI64vthA1/KwTA0BytaYhHf5JbXDIYDCfAXm3vSezOQIIDr2gxCewsCk0hXAccT
Ckx2AmO0vCK2bUz7xf0ZS9/3uiUsuRbKGVv74x2L0qtiGK0eEXQcgTMWlgF05J77dkp8tOgPRP1K
bvmQucD3ozvMvxkIZEogkWU3HCrNZRvwdl0KbHNfsGLB0gMAXAWom9fovwx54/39GUt5T8AHqz46
exWUX6t213wBDHLp6cdWxNHEI9/UdgmpsCEfoPZ2cEZfdVf1dH8mjrsWEDNVQm6PZKIYhFx+NCBb
sx/HbRecnG06cDxUO7N35aJazcmvcM+u8j2fk2P/FV6xtz1ldFBeZZeW7Opr3wNfwRSdMFbBOCVX
D4rgmoim9EMAc4ZpYt9yM8f73PjNAJD7T+YdYv0qw8fZUSNcEuTo4IZrC36e8C6DUy3LKeWTzuaJ
oQRiIpliabwxCBcIDEz5uWqmPbHp5uC9pSpnc0Pz5kXajQmod0n1ZGyQ8E0wKReVdX+EypwchScK
KvVBZ+dSGbEf2ZdXuc15ifmcjmfGl18ZqvA0czyS6bAmxgTC+otlMDlxuq/4cI6T2YRcXb4k58DF
aZamASpAbqfAFzDdscc6jZloJZSLvp80pPpY2fC/41lHxO+Q7DdnhJiNtzWWMGAmKPuOsHG3wN8G
RB3yH6X96nbPCGPY2cR4TaAzINi6eEITM7+Wrvhplzf2t2sBnwM+bJ6Na8ZVEnMjH2sA7YhlO+2O
iXLLR2leWhrpc4cu++UF/moLVoAWqCQkOGFKaC8+6UpjjbtNGpJfmGGynBq55YjS2MgfE3a2ybSQ
g6QyrPkCubwUkXLdLDdqsYyMbly3aH7R7CeaOFir20VoDa8lX0QLyfVFr5Bh3CGon3jo/ma4QyWK
SCoBJyyHAQWDEKDk+FuJhbrPrVHMW8OStqRDYV7SFo1Ie4URAvsyppOsSI/NdE7sx3EFjnNlXKmf
j9FvsH4PIlWXAfdJQ7pilJvrQ//VWgxygkJpP7GFJiTJkBcbwIuIZ6y1EF8kIulFgr5XlyKN4v57
X2XY0B0EzRCWIP8iioiJDmANJDJ6PQP2mxTYj43+gia60cOswBIcCdwrCGWQfnN+1XBB2Rb/Ec84
xQiyjmf/VxEJMRxe+gwYmTboFSp2K+rGtTpQOc17Q6c4Dc4su1HPXbFWFpz325X5g7Pw58tdorrc
c4IOBe9RLW3/N1Ub6loASQyjmzMOrjsiZLLvhBp6sWfq5yn/ktV6QKv+RxdaZGf5NxyPaHG7EQ4Z
EqXa0OYEK72ZqcOZtWnrLclBCneMzkDuQcF5Q+i0kzGYhnsndHx/pOvDGVLY9v9ZM/E2XaqBKiVk
W+MSYAa4bc+DpmMXgnif2qN8prfL6q4w2YCxbfL3GaKuNk5dmgPMRow8jErDoLBSXkOOqZGLxv+x
5cbnJ+kgwqbDZgy2g3wcQjLLV+XhRyQmQgZLZsa6zQ3agyTmQuaQE/FtboAjeAFjK9V4PSXe14cx
L7wBnBqz8DhJrcFsrSYYy7NgDUtXBXZBwd4Pi35BkfiMg9+qXdw0rhzBoQ9baddT+j2vv+nbSk5D
d9LksuRQakZt17by+cVh1/SlqM3M29vrY0fT9NXYAbfCc+PTLE94nYheL4YyBfrpGSbIckHJpLuz
vjB87VlRE0LtKBb5C3Om6N+bMmZej6cZpQP90oSl2dHAVFwEco+yyewUbKv3jR6WC85w9yFNKhxB
p79imnmk1fyyr4DnXQsdIMsx4SArbzdoYxpY4JynbWtVvjxJ/TfMZ6mAQ4RvpgrlYnT6HzVD1aGO
NRM+48lqqHquLz+mUhARqRHJlt18hLCba+s3GRsK33xCfZj5A8K/PcmKHGvAJt03TqH5Olkbndz/
EM/pUKr72uk8a35fZ+J/XIivwDL2RPcO2Mn0X9wqkvm6YRvl8ZnZyeDdPreXefIQnqIGWNr4ruMY
8uAZDRSaqlBQ7VfnMwCCoSCBk98AOgqtjh1GI5dRKXnFRNfup+dB4Z4Sq3pMf7ipxkQvhprxTOL6
WBP+qmHcMo9/0qWFSRFS/2WcSTKeqxGjstq0EOJkgZoPlOwdbYWVCN3VhgoPVf9f388zWNbhPuRe
iJMQFyzyQtyXr5FhS7oleJfa/Ha66ceTn8QJ2U2U2ANQ+30zCqKiAWtRWV+6nYAXknKQ90m7vq01
UD8s241Q0hTezQD/4m1vMjpIFiYKr8JHALnCJdM6gXOR1qXCki20QlsAvEVWttsWuea01wD96dif
xwqmLf+aXuMQqFSJM69iYakHjE+sWcLGzHvWpQBAD4sB7JGIPXQ0IlHoc7TIAR0IXT+j9kjtfivH
069suibK4FUVGvF3E65ED9ZWyZ6vtEaebjoJvssn113FLy7/A3M7MWHNjgRE27tuw9YZ5KcgQQ+k
ZIex8vT/HZ9I8CZFIi2vonLqRgazuC9FN5bJbP0e9fHeKgO5SM2ZnujYjk+i8OIm3fiI3P+9TXrx
pp5Bq1Cf8x0yGhbyEDqAJqYW1Uun/Qa1Az4cLaDPsEnX5cwgFLmntAuVz/6VmLSW4Qi/+6M/KFxg
A5QkqlKFp/+MWsmWJPIWIaE0mZdpvFNbr6JPMTqVJGUPZcnQliDwzfmCKOlEt6rYRd+uCxvzKFXi
Xx9GQSsCDumRYZBbwDGmkCGcG3UMMMQcHBXkG80JJE6d9cPjeCej7ki6ZRWL42HT6/oLnH3aKILX
crsNncn1DXzZjC8CAzR4EFRrhe0qYOWnQVzGOunH2WR2k/kRsZ6lbutti7Ow+S3TPayjLxQlTLw0
F6cETGAFzo2puq6KdFN+miDwiJqLqchPuyItdC2n8jZoi+8+wOCp/srVfzQ2JXklc5sbIwbBCE4t
/sAiN3Q9IDzYPS9fET3puSZRJ/fnV3sGjprasB3WhV7G020M8H/buiEAQkeRZMuNTJD3R7tJLFdz
dBbXWcQgzWZCuuDtwkcz7uwdaTjJCk/rzna/XtE4HSsXoMhdbL9f+mpl1wlchPw5Cr68lL3YGx7X
lUSQe6VjpTVHpQeI20xl57r02ubH+Gc8uMqsJh6NFqGDyxM0EPpJoWBFxixsBvHWyPzFY+aV6gX1
eDFMWt+TU/gF2zeRQygb4OMhPzMYxV6AVB9NV94XQ/TzxJdGparBf2gy6YgyeL+PWEi9QL047fDn
af6jLwWUX4aVtKPFg7pdiUGdsjwqh5F+qP8V4r6CyDp+LTV1zKIJ7HUKSy2H/xJ0bIYKMp3LhABb
YXgJF1DcZqVZLnVtgXtqiIjbq8xY+HKyha1+vyJYJY3LDDM5aXbGgMexevZ9JqGp3y6SWCv9we6Q
hutnHUaH2NHatoFWhvPU13G4YrGVbO7sU22/lS16bBBRkE668lRzVAd8VL5o43OLRUCqEkBGFMvJ
24+oAcFYGHCrjJ4pcvGOxberPg3+JvcXPLHMrUVi++OP/oT0Thmt1nPbuhipR0KzBNvCwUI5Zu7P
JzGc/hjeoMD1KxfSciEbbCcOOuPUBbSmKnUzzaMn76h39/6hC29BwASjbLkANZkz5nCeio9El8TM
FTmnwJQF4+QoHi+DTc50E3LjJLrl1xamX7exxUQJC/QhURaoKyVyHTto4zIjJ0GJzp/hGlF6wcp8
+MsTBAm7d8CSgzUelDyhu9Zd990OLRc+zFGO9qn++xFEmcgSr2JT3LzgXx6cGiSE9wz5URI/w56u
isTc3fi+uV0SVNtuOmaMz9FWthbpjaAn7BqCNPEa3FAKnLMZYY/dsBNDx5nYe+IfaBHHCfTLc0us
3RbP77EBHpZjHYyXVVG5K/w8v8zH5ZFOLfzDAHjaQBtFMwtz09z13l1zyR5GETEJ3cK29GwGt2UJ
mw3+lTVmgOWoPBUi/VSSHMy6qH/HpPQR8BBtOTL4tyibIsUSHCtE3yWoNnuElzBVYAxPFhP+niow
tigeR+zapsB5VDkGsmQnfOqAph49VuQyymkimq+XxsW0/65P5i9PR9GZNVMwC8gLhOfy0TkefTKn
z/nbIQQveFWigzmcg04s1O4mLc9MBvqYEOpKAwiMK03A2MX2HfRBP1NlcA+CseBMqbJjBalfUazl
wmFB9T+m1WNNqXzA1TublArp2rbKl/7GSd8xB2byRJoKyxXXPS8Yir8iLipFBRl8q9/lnUpUJPMd
ARFmL9O5xDayQutta2eyH+xrwCRr72HJ20FWKBCDYMAoxv40bKB3zeWNMD1f30EwIWNfSEV8yu3v
HWeuA3ZdfJRH5MiXkSsxKIabOcHfS5yFIcP4mhikTnLrM+dEtG0qHbWsoLl2lmFEcbFtHO5nNqsz
HHLCyOy4fv3mQ+Mc9FwyaII47EdKuiqq6avlF+pjziqBW31lSWwx9dJKtC3BwTy8FS85Bs6qDdMf
oAUjYPy+9m2fQ21l5tKMUxdb2hfaqC9+QMT/7K6spvMlXsvRJLH3zTwQ4T6/zrTEPuWyUQQR8rXN
aOlpY+HutgEvYrEtf7sEMkEQCfOYFKJrhx9GoGAeL1LmmSu5yAy52Al3tqBlO/tunYm23W+Z4qjc
J1iitQX1C/R/Em7LpU6TkLXKVqX27iCafmy8cwtZy6lMm8yCadJJg0zB5nwTEiizLhMQjTAxM7J+
Lx0dEemcoZis8Mwulmus6D0fY8G+08ArFl3QYk3bsVf8nKUiJ2jixQdc4ZBrJQq8AHn+CIyrVEsH
+Bg4cW22NNWjAZSklY1m6WQ4yokg2sJf19QfJNcCpKeIvfp1SQWICmaB4a0ZqYxGu1+blxquvwOG
TChSs7gVb/HnDEihgEPTdWECwPewHJuZ+c7zgVedNL8RQ+8n6Qet1Gt1EewNXceLqvI0F3WtKT0j
RJW+nOYOU/r4r64seLjRooZhbNqQNd8hF7jWWc+PHQggDJGESEQ5ulgj7XPHvqDP5gwwgo9AfOgv
MjCV0zPJXYOFIYoGvLG+BnuPZNMJ6bCAcwZglv1bhUS5IhC23eGTjEbVc8V0Jf0qRkizGIYvoW0A
gRCUKZri1f94/nCmG3S5mam4fAcQjyq9UIqYwocwr+f2TrjWO6r9TdEq6tVIlBBftr5KKWe9XAnf
quQXGJDaGN4VI78Z71bDd3zApM/PzAhy3LYyLkuSRymMh/MGV8z7GRfRicj7SydHM2gLxRQS04kM
q/mbc5cesH96tcsR6UoCXZjSP6CPqi6c5NP39HunfrPagbr93oLTCh0uQ4Zzuxi1/a12fDGmyTfq
5Ox8AcEX2PVapqm33TNBCTWpfqS66e9ULFGLusa8tYDPTjFKWF9YnDO1okMlwQRWTs88ltFkX91t
nmfe8OyY4d296cckyABXcjXb/U/ZT2Uze0Jitp42AUThSW+ShBKVm6qocc81oAGKMSm1RBDC1RTr
vsvAQca3SzPYME4lOE011ivVLLJZKljFG3bGWV0vok0ush+BNTM5NdvkAq1Bi0vuGX0mbHl9tWuh
GJCSRl/BnY4teXwE+Q8L5TUrV4DLVHItzXHjP0kKyhk9YBCLoPi9KWREsn+5z/l4KVNbhlkkwOiJ
PA8iGsbMYI9T3FJcNSLl1+z5m02GSrIlL48lhsou7EVT12lS4Pm/Hh8YWloPCMLScaCdy/H2rwf8
YMldLuRWn7e7K4XQY0YiSFRuuAEAdG5Yzj9QT/RNH9bZF8k5fcB2MMXVxDUFc4u+zMloCSv69Qbb
/f+43HUjBxxl+yIm3HbvFqQaZNglfbbOWZYb4g0XGsIweTOCyouKJ+ZJA33CkeiEg0kICtQHF7z/
pi1Dr6ktd+lL5t8Jg9AzW5oBsYSDjUM2Gl2QTaQpro17WuWfG/c4JDXUN7yzzPoYxf1M/BW8jH2M
mss+PM3uIv12yMWULCiX34at3+SZZYYkxSlNLR6UuOQFcxRXmuk4cGh6bENcgG5xx0fb+8+Q4K6W
MFzYhdMQQzfWOjq7wQFzhPfHr5dQUIl7+Yb7yoH8a8FChbO6rA8m0Qn00ODMPpxB20C0C69NGCtf
oLv7uI3yM7iZLBHjBUzEmCbyKo1aC87BO2LQQr7+eQX74nWdUPu3WtE+dH84bmv6HMm4ttX4+53B
C+giPW8Ytbt+IUTRX9Q67+yJUe6oPkPnXgs1uoqJU896uvB5MWqmvcILRnLGR4JJVX1YQRxZFoaO
A60k3h45UMV7oHMhyDy7NDLwi9Fb6gi9Tw8UzE+cHW5PS7vptZecA8mldmwnSAYvJ1zbRb3cs77I
5bc10OoTUOrcbRd49U/f3KAcMTafbdm2H/cHkexMPEikSiKsxvOvSLcbWw2wqoT4B+X4oQVg+464
E1I64gYCVm6a2E//4J/5iHW44VaMdiOWZYmeX9sIxvwl2BzeoMipb01UNuYvo++OY5tWBAIc28aI
X8CWNJV8zEESY+Cgtb21bSjdDavHmG+xoZGOff2SNMutyclk3f63wuutvYpCewuvaaqjv9uLpHGi
xegPlS0TWCUe/CphYgu0474/QMZKx8RpEGJ6F2dn1pJImZ31xzcYoVs5FkDv+n1jBdmlAdb6OFTi
jhSEhrz4ABnFfwYtAXIwtB95CpTKtDPEUtDGj5yrhNZQCmc1okOz3dYnINP5wV0w9JqW7tU3lLki
1G03R8SgL12nvV+gWKkBE/5hl8qilWybkWHZBtfUQPLVu/C+842czxOT4547Ww3goVdrq28iuTpr
QczPBvhHgOq0taMhUVKPzKPZrNxjJ4uGU6fQwO2t1dcCByxrkG8CRW+hqGLs9IAJ7VwW0wGGNlg7
4zk0ltSbD9E86dtfYeCzjtDCXdsynLyFgjIuzeHAi1UdIEao8whR895YbQFsz/gpIiXCn+9IaAOn
lvOVQ4kF8//FzcGplzZWAyRoEbwQayT+OLoCpC6vhXbJnYzghhFKqc0TnVK4jLb6PeCt3x4sfgy7
Gn/AXTh5heYZ5n2OLRmoj+RlNgU7x5rQ/Cu6YTtO0bq7VApNjSpLZryDjDFfhjVoRGT6q/7VKDDp
xzTXCYbBu5DrSLlfimzqUxVIGWfTXqCQl8BWYAhnuGZCy5o/lQKxkDv62sFkY5F+fmKWt7XJo7v2
6hTzuLNgv7qVEDrLHZB7fmXOdsRbxLoe6IiOBByFGmHbgr154r0HjDXSlIpy8+JQPyBM872EwtVB
cehLQtD4tZd0UIgfqFWeidGyJDyZQ09otO5BxKQroPz5wQzhzHD/LL2Kea/RO16Uzfxqxuwe4IgW
EZvMopCBXJ7R8WzE4kT9kNkPNp/PV2DYGV1+8+IafTTFvoUcqb5XXJl8buFQZB1d/mCABaZxvFPr
QgcxbG8I4r3yoF/0EHf4iYglV+CCAuVqtjC/Pd4RYjczGFLN6PZLPg9I0/363ueF60e9yFQSHF1q
CV5xoBNE5e6EEovwpn+v3oH4UAb+n5UfzDA+D82v4u/Z1Hx1CzhkWw8p6kyHExgWRELIpjU6Ywxf
lfgaS8bIOvzJcXS6mh+KeqCmcNJLXhozo/e9/MkKAjzWZwL/APyUd2vBJ+47CCDHpPuMu7Hvj+hB
ungo/NtwH6Xr/+jHikaBylrfw0JNr/PymiFkIhuu+PBXrOlB//WKnRDP/t3+qdIKgpLr/pBnzVVc
D+By/s4xHwGvG9tHefbYo0p6Hky+4F1huaylnwoxK+m3bqlV4qSUzOCg8qFe3qjzz6kE0XV0is/F
A8qXFRdr0oaWWchNO4zTGfu+wveUbzrL27Pk8Lk9OQ0o8MGf/tTjI1ySF/OxHVnfoF4FglYs1DzC
hTmCrrKluwBDYgq9RaPyzTwU87WnxlokHepTpaZta0LeUqDdJfoBHH8tk/NgMXM3qBrHrdr5Yc2l
Xk9p6lXI5vkqugnt1nyttKN2/4NZ5VHidP+aOSgsIE0u12JQR1hWDA+uGnyXoSd7AiBe1S3moaWJ
oSbH/VoIs9SamZhtSavN7VPbsxp9sTF+2+wHgo6LMHpFMDNV9PrxVlW966qoKVXi6DyRNCjbgCjE
XT9KQP7jbiobblryg1B6jeqF2sD4adSEXNoAXAjeYsNd9LB2TPse1buA34Sn4+0f6kZEfuFvde5m
jowIVwTCWSbtg5cKmgMFNVCZYEk+J2RT2KXHddFwKcV7zf0DRzEhmuKlfDk71ztpmoYW8DWQ+pmB
s3yD5a9Vv1dQlrfflz8rFiCJxCaeudB5o4SQs51q1Z/HI0F5lVKHcvJ0c1JKhnDaQY9okyl+LJwq
H8U87sCDgxBXEHb0THcsXQamq2H0VlVJljWVChrboNL3T5iNLIu5FSXf3iR/P3TaxsywGcW5UxMx
GAC9w/kV87luAUmhgTKAfR2fUaWQSPlCFoNE86vMcx30KtaGAHHicBoqmKBu/haN6f/Ym6xwwYzK
UxM7A2HCPBjXj9zQfkYhZQRHJwjhP49vvhiTSK5CU/hsQ2PI6cUQvagqO2ruJ9arC1i+iH+HKms4
o91FhSxQ68EQUyRTL2E/cku5ZUlI+6Dl01U4NxB4KUa6+o4/VC9SeQtdL1E4IobyoptvI8kgvoTC
DGcj7mBDYcB1QNm+iNpPp3GjDkvfsXvj4VMU4O5N1wPdqowBB9wimGq+Ij8o7OPe/YnY9jCCtysX
4ubewcE2ZDjwUO55AV6EJ6zNa9Uy5ml2J63T5ipjZ49bVSgMCuRJK3Ex2GefK+kjil1PQBVIvq37
DmPHCP0knx+EZSPyO2W4SC7ui/poB+IqtlI1xMUdZmAmykQwA1mBx3F5aWHfU1v4vd54LAT9WBEu
G3gHnn9wOPAXi1JrKD2fkHXNubEgdsSEiMNSV4jpHrZ0L+iz/5MIgAUaaZ4w0XsNUvIPP8zW+pBo
eaRRATKr/tZtW5f9yjhIhwwn9REk9uKuCbF8QT/YxkXX4G4a0JT9DzVMLvepQ8vDNM1u+33KH6Cw
jenQ6+hBNn21ONUiTk3ERlrXs+DasJX2NC+QTbHhyze3DhLo07ISwsHzwHRtYFOmLFkSRUVK6atW
JNIX2/Ea+Gc+KOd17zykkXB7cQwY8kMXoKobZRjhyLHxyUz7+sdFxdO8VUVMU0l9d1HOmsHPfDmp
ckl/+XWYjHYhpaZv9WFSmnw+62IQ5mRbBiZBSPlTqkWW21dKWyCcTZA3cIwE6NxKNcqiqyev4qpg
o3n9Fewwd8ZDJ5dzFtNzx+FCKSVwPuo6qY7ocJR7i19smAqr7TfLsGw+Iyl6rdZt3t6S0xixp5lw
LCS6rRkUl9RjcSFGDob9yfBsWIQLtGSpEukdSR6+CY1nt5oa2W829Pc4VYAydRz7jXqOxPznRdlV
SX9qSURdlUDhVkZ9tEsAHVK76hTapTxhgZqw5BDPfn5xLKrXfO2d70kwTlE051eGvd72bcxOTbDD
xJPxx1krayo5OtovdW0dHc0Jrj9x9HwM6pCfJmDcrjSUvOtKUHYuqknwJ3JG1JddiqzASm92s5bw
Ptc3k8cLGa04ExQb8SH5C+KqUanKr9VaN3MAFN9BkxM5P9mADNP5IC7hcDIoi2TVA1nXYSM3jFN9
isLREVj5EjZzQCUgCCpZKYhzs7cWMNRk35b9qgksHXaD/1/yYXIlv6GKbst4dUvNcikcQ0AjSEU/
EOzYx2To/NrJ7YinDA2egdQpbgMI1JJ7qhEjFYrov1qFSCLS/yOfuk5i51+zW0AY9iOjASCGhpQj
jS9vAQFcz/bEgVycffam6h5G3Reno+rJOM438wmKPKlx6pgH10eXA8xLBwwpnZ+T0u1sv2BX2oLb
8R5QkJeHDSigVwgkExDLZhszPRigZYkJHg3ZrPCzEwQxBwRcS6/1/OX81jnN251CyY7nVn860LGe
FOHMC6yc9xWY8OP0M84lL9WQckiLxtL78gxd4Gnt89jnhTM7lgGixcIwKFl0MFfsAnVycyb2vlRW
kEhH+ug+8pYeq26TozpAoL8zlKqgOSqP+/PfxdzuNiUKw5cL5jS+NLOjiBimcFooaQAIT1B33ZRE
CchkwXAmkkbe8O9bOLOP4QggaygVKKBP+PbaVV5bEhMKeQ36odlFY1MaEcml2WwFvexbHanDXB4h
xqOzAP/DXWbwV/gqY/vBuo1bsTmYSvjprYMSjp4ro7sMdWXes/ppZ5GnnQZUoQyLiaiNVjo299Hu
rf35WSX74kgkqOVDf/OcUbVShN+vh+u5u5Y0fxs/oZKqcJbmjO7Hf1ZIEQAfBEZN3indyUANVezj
IiHChwdvpmtt2jKgT3RhF7LrtONqeOpo5akZhKWdheoyiyV0l/YtibJKniZkPxjoP7c3pMUp26V4
zT2irG8WRYayOkgtnHDk2Y6OU9XFOWjXOvIRvHONPvoK94aQaigNwX/9SWx/CXfjPioCKudap4sR
5wBmD4KaAHSpRUtNgEkk/XVU6z7ox2hPjVnThqaap4DYUqy0mY1JpMqV7RDKeBbmiFZWuxjM259Z
F+oOgE5HUGqTpN8dJ2Mccwjkhu4rIamIMYc4oI/6R2CbETto7soYRruLRtzk28rBymvxelQfhpwB
8WcQ0zvTF/Xl/diAq38kEBgTJYtb+s5akCovcEEiueGq0L2ukHCZBdipEslXAJhw5AtNfJCMXuT3
4jpqPXCgbcYIkVkBEva36IwAmOugTXNP3zWzAlvORpl6Os5Nk6Rkphocplnbcke4dqQJEbQFwSuR
WOllSW0/jBFRMhTRMSUJ3h/Z0utBCNpzEFGC9DTS0Vj496oAuEE+zGHUB5aCozcAywFlvsxyBjC7
6RvhCNZcXP2BK1x9wpaZzmIqS7VuQcQ6NmRg+eb/+J9QPSPpaoouXc1ELpe6gbZLEuqxiQc8wA0R
LhfpOCQ17oam17FNXsipsjg2VtHJL9cLYWvYeon/mECbl9Wf87uFQBbAx57iPg+cO5j0CjBTuArx
FuM9ggbBiLdoUu6mNYFDEwP6z+NszFLKT+n2cE5LzDffzuvQ18MJM+tW43E39aufktlE87M9BcAR
vrPOmmK6tyz1ngVsNcU3xhqcCrG8d8bBHfKl+id9xThH0v4HPhi7hadqBK857yf0XLIl+7o/71YI
ilkrL1+B3x+AQfhTb3lRb2l6wokqD1/j0aAycbik3YEvryx3MjY1r1UUEZQzCwIXegtdc8Rd+VY9
/y7be1C10RXtPC6dBl94JtmjByJIxdqQcWl2ATQLERXBSRfqCJy99r9aQRrtPemr+l7EKAsDlpuw
9+92i9SY/7eUvCTa0GG6ESfEn0cctSufglXPPIWT7UCNB/CrjCBJpL61Cc2ZykOylOSskhLJrBFW
ByglpVBoi4nPg5fnGumw66WWa2kWSfvg/YCMBe1pxCtSz7jWeZIINTjfml+5CndCRNMsNk9BHZ0i
JaQtm+W+cYVo+xA3EvV+Wc+aw8MiHO0WhqkiPqPreU454O3EAwnPzxpKkj8ulsWXH6iXQysgAVLt
OFf69VM4ltQXNuuDlVXxmxQdnZ5fLeGl9aKuGB7dWS3mKY0tisAvr8Es+z+CmCvmxshlTKg/RPDB
pOk1hRZwkjfUFgssN3bnjIm725EruWE1GXSyqIGsYXJkKl+HVHxxUh54aWOju9m7e+8KcqX06T+o
AERxECuk1Evs7sXgkRysGPfsW1oIuilNPZB5SGbpRBGkYNGdQPSkVAOxfPjgvAL4jyoiUehCwZQm
U55J99rG9/VoxjyWh4vJyKnjuQEE0SJpidQqj2JxPCKmNxD+XRLiVuN7MKIS2FY+WVOKKefZYXwR
difMhNEbgwhFyMvp+AXEZGQPDXxyucrXOt9nHuer7o5tYdmxdUsVGjHR3Y34EDlPE12FJzZoEza1
ttPozEnWM5IsyX8LLdnhSxsoOuF7ASiBTzfEuuZNgxzwgaKUCLerJMrI68rRFM6OrxHo0galIBsq
6q0AsuEma46ZW4fRcdUYzr41r14VuRnlALIp/XWCXOBSdtFh0bt+AVHH26rzBrpbN48Ig7Jq/tQj
+NBa3ocCRgRT5FdHc8+ny1FmbkYVo9/CZOHcxezqdXxb/L+ABciRXysrFoKStd3KWie08kQe9lIs
6V0r1W6EJ563BOpRKVWszJzmV0UZfJTQeprfeYHWOPUoWv/5/R/7p4UrmxdSkUsAMiuFrQtKdkDb
Q8fXw4x3rabjRqaLF3bKbzrgwc9DPCDtDZjyC+VQGVGT5YyDpFfz8D0ZDR+djju4Nf9btA/YFwdt
jmL8tOu0MKmdLfuj+egTFuNKjCHD1FHnGvsQIGWwsEd1RmJYoAuVGNQj41jX4x6wnQ63lEyh1f8v
7N9VNc8KetpKfWbIDtBXGiYQzYk25inIFwpcBtyzGo5v+uCklf30oHG01LHvePR9bMZX/dKpKc28
r1+lhP17ruUdHrX7zbFFK38c2BpUcOSxG7gwpJ90To8PR9hzwJe2U1zPuNg7YUvvepb1RdpAa4Re
t6mqBPFmPRUz/zGbBI6v5UDbfzlF1j6yoHND+jTfbaWDHD2IrAO+fgi3Un+By5vM2IYTyqI/+imI
gkiqFrLV4uk2ywFB46DmWAuajbIKENOGdyNPO+9cjwPvD2MX73PE+v7F6LtfwHIxioXWph7Vwevn
IFCJKypXhJFeMRtrjWDbdkpBcQomPBMPEI0h8EVZr/5oTZ6mdViIAcyYOGVniBKzgRufpiWN49os
Mhepz7RzP6GwlxQBrZ51fmz+ywkU61OH+7UCdtni2E1k5L5WNCrb4djVj8E0Ii/Gd4r1sbMr+RTg
OfBHGPAbwytHCic2UnMTEHyEbapcdQ7WcFhS/6b42T5D2kskAKZ2F6ovfPexpqsu0Js1jbECu9PV
dzCpmxsvTE/THraDeRDX+FrUem4YLGhf2Ch0QUI55BGfl83xcXCjNVCZMDD2gO+Ebjt9OPmBe28F
No8qny3zqxPDmEl16c3vue3UeXqbvO2e1iQx0za6TUWv2zAfwOxr1uVe1kU71njVCU10r/W+ayiL
Uo0KyQNkLGXOM1U6j79bbV3gaQdGTKWWNbGVZTq+Lx0NzOBXD983Zse3KeEXjl3s6SRbOBmiIIl5
wCqi9tkIMS6mCHlEQD2uf33rib2johJzqR187bm4/q+DhjsquaWdkAIEk8zGftCULWmMqKr3MaAH
mSABWXcxXlx7o5yCf0FYIzQDJIPOiqcBIABPTg6ODosgAOFCT75FL90QpP2XxTfoeX0pjQBb1Jb0
JdIIsNeMe24BwYfDc9pEf883qgFiqVsgYeDn5pHksFQe4TCfIlvhRjtG+hoFtbtfOvgJjqwQ6XdM
ZTdt/PgQS/vUKW5AisrXnzTKflq5bOjsW1xLNtz6VRAzi4BzPPkoz9ImN/5osFq2q4ZpnZLl26u3
pKvA4kth5tYEEwQ3LJsgwSzcMywOnR/aY9qiRMJVlNbA+AD7ylcPS5HVDOmH6gcTPRZqPh3sFZ41
xLDAqk7jN7Qv8Sl8bBXB+ds9wOZkht22jnXUl5wdfdMxLLMvBhe7ZpiY9yfybQg5K005oZ7TN98z
/WXwIRYLGh5Sc/1hLEBn+2vZI/M3NsHK2lror2YgGlRooOGyW8PbjXyaxx/QcbwP7Ju11m7v6Jd5
rO53rPYB75qvBVZbJF6xxl9d5afUrbjnPvaBKUEcL4719cMliuX2GVyenISqFtDE+C7YA7cXSijV
QG8F3dWZfEKbZWE9HXef+SC6PRpt0C162x544LxjGkeUW5BEy2dUtlc0eODkTPF2QRSdm4JdVAO6
ddRZjN4o1Y3zFmuYTC6AOt018eI2tiaWlEGLnC/95i6zeg78GOd2NOqtt1jEkk+InKBY2PsIBsXG
DpwwQZHyMQU5blF0DUN0yDL2dqNQPF7ckJ9ajIxzU7qp6qGbdV40F8qEmDyzeCMqRo4BxaK0vyK8
KVZtCN8GqvhKVSrFugIQIX7qYHLXa+WXlir9/ygWoPmDGwkbGN3g31Cn+0me2en65RRXzXMjlHBh
2vcHj6dSrqL1RC5Yodj0m2rIgSct5MmwAB6v8NPHnfy8UlUFwhhd6dCkj4kLfHsgWhFC55gD1ZQw
PTKqOcXOLzWIi3O4EFRIptmkiX3fno4UwoKV3AcW1QwiHaCyxEcMJhnLbIIOqNmo3umkFH7PBAj5
u4ZxWpMMpZfVxkhRtTU96hk6ULOY3LP2yj8tnF0yEtzM3Jw5rA2aUqR/gY2cb5dbyeqoz/BaHzTa
TVk21RySja6LCBwCv/TDe7TlhI8N8uChh5WgEnfwFQMPCpa+cavFfEoW7qWqyHOWKKeWmyVGDg7h
tPb1i1Hf2fI0LwsDrksGVgldT+orK9anYst9wvaJeqxBfZbXIeO5QN1qRf4vq9NAE2ancUdVbg8h
2YyffDCqq0mjwLzIr2+R0gSxe9uTW70O/O1nInrGbOvJ0SUi+HyBTiG50kigz+Kd9ZjZq0lR1XsK
QsqYlsj83js7IpStwd5LiG/PtLBV55aGziwjU+RqrweqOP0GRFmQi6GSzWxFEy57zG1Uj59y4CXJ
3afjFEri+oCkoatNwRfmlF/TY+QK0QNiQwApmpcDLS3N6vJhIa5d+J0ZHoOCJjq5VXs/hwidwnof
s4bL7EV6Lz9mCMFxSlhCszZ0fL5qjjSnesYKxXUGWcCM/rOb0Xd6AyuNAcRCejVfFtw19UlvEoCf
TsRZ7rENdeHi/njj8J/bxS4hC5XHOoECtcxHryvogh2lnDKift9eqhGDxe8uS34ItuSzON3WKdtC
jVzgbC25d9JwVry6R90SQDvv07ATjmKo/uxNqw7lP8fLEOwJ0yhcE50msonRULvhsR3Z/ltd4xFF
DTjY9+x+NoMTTMn7cONO8Fg4WRovPmHxzWx8zN6ERo2mC/XrJ04OAdQK8o0IYm8I+b2BkD0sOuXB
5yPSjLbLxgRBnIXzKNz980HF5spcZ6sE42yAYt3ZAC1kAIVF/8Xd5qDfMSYV1DM3yrk8n5VvnUSL
2UYTtVo32LAyZx8s2BgaSDHPRkZE1+Ft9RZXdga66OLwJtkM75vV8LQVK/b93WmevD29pqq0DyaC
zMBvCMciw8Cr41rhu8qx8lqVuF9pFIL8+l4SA80+R7ZhCEzqC/q6VuiOfu1s8bj/oolNfDaIDJCz
XIgpNstYjC3QmS9nMIKfaTfCq+6aMDRx+QjO61hvx0XuawODZ/sxN2WLvu74RNN+O08LCh3zC3Xw
KxTz321jq6TqW/d4beON2H2UdhY3a7tdQxubiZns57wikBXlTFFki5ywlSipO0F5PEzp4UXRH12h
dAnFRf37mX4oZT3KmqoN0iMHeET7IoarCaYxbrDzq1WVFpwaEcLdFEo4aG9eRyPOZOHLp8DMOp71
roRk+F9XKfVYMZp+A/opcFzLEtIft6x+A64tCXbmWzOJZZQ11zLDFga2t1UZDjge5EelMsiUDqdy
VnvYpswrWQXvAk+2Yesi7OWW32DZqZtg1hP8U8aTLerRYDwjmM76iDwLxSZQKCmo2FPZdNslu25d
VZ7F7duZ30wcJAXEyGRF5OrtmgRypxnqv3A7nsP7bdhWkZB+B4NX1zNlBr0H6k6lMLkM6Gw+43Id
xrBKP3+bvofXZXcTGDT+UhYvjuPmBi5J9x7+3KoGLkUjToBAl3ikfOaRhOVL0F7V4fh4JkC0e1pR
Ioze5eU0URjwSRk6IVkLkooRGb+V6iTLtXe1I4iuFyvAkcvyShaC+Orvxy1spswKcxABpEkXWM4o
XYLiqLCscfFwVXD15C2R/q+fYfkQhFX844PDtcksqzq/WHe4/5+nBd8lKvhbipXO6NYaIq1d2EAH
rZq3S4Pky+LpibZYW7PPQCg0hyA7pDYfC2UmsQnQYLk/VNMunlY++S0kQMvubPrxwk41e2k7JrYp
HWXAH2zm4iOvGb1s6xDUwWfqogh7jm1l1QGsT+XOZsP+YM8FPQxppzquOoX90JZyrPu05+pl+Gnj
2DtxRtApESBSW67B4T52RBSSR64yx5XSQOzBrFL6dcZgPxscuF3JfXDgfli275Nh9l0ENwJ5NDuA
BqhEeKypXR4/eqL4axkc/oH6b0z1oDn1e98C8UnhTTPcu/as+dLYaPufz30bT+erP27hsYrvnvE6
qd+hw6kUJ1UpnCMhINx9mEw/rBQa7mWEkJ+RzUvc4DHg8XLLlrZYeNlGAgLg0RjoU7krKwr0bf5h
Byv41ETrMBK7AZ6m2WRW7mUNPUSO1tJ/b+yXeD6Kzo7fFovecW9y3BWlfsZTImOKc0p66Krc/maK
dWsss6q6odt1/BpKmYWwBLuS2DukQ8qZv4UmEE0A1cX1u/Cc5iuTyq4z9LyJyY+nPaspn5wZpJyk
4bSU6FrxJE77RQRK7nFl2AYshI5vbb3n/cVB52iNN57xkdGu1LIM9uIHXK/CPWmhL6hfkUsN2zGq
LEF1YLNJ70NiW4Ee8kHrov/HTjOHZOY+/xjj4y0wbEt1D1HINd9LAAKR9i9holujjO1urQFROaH4
Hlat5qd3lk6Row8HcT6b33MNSWQyDAAo3P0uO8FUeC2GEuFM3dmQcdA9oF2uvWeW4/nNmpOkoAVt
9XrQXGzYC3xEyyHpu2/nZG1lYTibSBychb7EYqmsp8E0VwudozJ2sT4toLkPXrlzK8IDMAUqiF0Y
QkA4md4e/qSkQKJoAwOZaXn6mRymrIj2ouy02DZH0DDgljCQryEWg+HmHWvQahIBCFvl/R7BauEs
2791npwZXfV7y2EkJxwertB/ImzL/bq4vxg22ZuDhznG16hmRGghRd2nCyk+Q1S2WZZQObA4JQcI
y4WNmDFDgLjl0jxLOOueJaWM86OTrVXcWCImPjD/82810+vz9iQwMdY9PhMY6dI2Xx87MF+8BTb0
hhf30r9qenaFeQYG/b+SvKaHmt9VlQOuvVF5K9UTw5o6YhZC5wGUCQbwNFJZoIxjHkCRQXNJB2hK
t9nzE8M0nBQjRFHI/KzLc2jDTsAC7QkVarTI8+WASVJMxWo732LLbk7BkPMSghnJv4q2Pfxh37cp
1bI/3nnuRw4ojN7O+JX+ux4HIhYvFHvS6NuaywJUt+658KZqGSAzp2n1G5P+jKESETV0jbiRmbGg
l+xL0kO7rcc5L7L9OZZcSJC0ed7b9+guKtImFCj2+Omo9uw4e0qXWh8fweBVMc7ESdHjhpx332UX
mbwkjh18kPYVlsdDDIln59q5+BJAdhzHJMsK85d7CqoSIHJbdALBxY/ZmawXiBnHD/MKO3nuwZU3
ULqb2DLuDtCn2I/NtfBrpMqdyOdnz0U5aczpumSbAH2wOnkLD55f0jnzuSQDSKNlUxIJiEe3nXeg
IIsQ75wNYSwtaOgUZM3dGrZnC+RgEDcdkeAUoP2DVHfnQ5CzF4u+Bl2UPT7xxHEcVVaB5BZINAHK
dE+dsD303jLS6pbe2ykWmGji0d43szZTPX3RxgCdm3iYaeiQcz34lXan8QnYRwJJt58QWqTqCpIt
w+Kmz+CI9zsSZ+/GXvIZur/9FLBp7fi5MNuo1pSMDHBp0xEaFrJzdG5RGYEMry43MkOJtcGgN9D/
p7MY7/Ykidocj9vYHLfNNvSC+FCtA5hkbIFCotvqrSgFfWuub0Nw9cV4LkWlcOWNumvI7iQHx0jp
C2FsxcWVlwkdP0VGf5o85x5A6pzc4/D9O2cwwZbIVSvzGD3yk60rcBS9s0CLxvW+jeEBepM7jZrY
CW3JaPJfz1AgNi09j7XxNqZt/qtYF/Ng7LUhWcEk1k1iQPxwlHSoYtVqqfTfjsET+wHXu5cnBwSe
wqiHPFZ6i34s3/PdKq8AbfBc1Kj2U15cxqBflMrujexKO0E/F266S1SaSe4KS/+ecZ0MihBKgXlY
HeW6BfiPwBgUyi4W6I4M0Ld57C44Qd/djBXyU8z9kfsf8RTgwD0j/HHFOwGaueuk4QJsGxcAJyCK
ZcvOMq1l5OEmdofnt+KorxILRduPfhuWJrBN43CIXgWZSEWQ0OUvvPS57TesJ0TXturT5cIur50U
PB4Yq+Tq8atueVe9tC6qGGAQYNvbrT3tyfzeSa3ahrymmcRGVstIdqm1w85eDXKVBAXVYnetCc2o
I9sFFXtqzl3i27TMSTIDux98Y3yeOxvzK5thut+poVW2c8mwTb4ibViHL/rWz0OZeXqo3v2/duBG
2P+3hcLhWwf/d31onYtbm9UqXOT6XBxaOltaJDQRT+W/xrTX+Ty5q3cwtMyCmyKnXSxeJxJ1W01N
Ba+oRXI5mOXr7nNTGA+aUwOzsUFgaL82kkfX0U0IpuxppS8jqo2ZXGLeEjGvqt78+5IVjFgbK2gk
0bq8Y/g7jiGrydzS8QQoehDnWwrYyrUFSBLnrkmADewF42HoTXP2e+RC64qU248BKTekW+YnzbSk
HH9r08f351nGDoi0IQvF5n7ckPTUu36WoaPzBXuUIVxqLEurZC7W5zjQ27CHPaTXUmJ7wnyUv5a4
TRRrE/djLgu6vHmihMcJRSaGLNaQnxdQR+wZ1um81rFKS8vqkpIt52epB9SC/NozEYlwoWdkXGvw
XOxmw2QlLmSMwynt+lbsOFMcJhD5cVzCc+OBMHjkNkf3HZRNAHtWLAQ8PLFEr0B1G574aQ+LXCYG
AQIQVYlnBaEV1mtcQGi+IGMiGKnoLZsHKai3ex3PDEwEyIYjz1wT8i9gL4A4Jn3U9QDmoec9M1j4
cH/4tqnnpeUzB/32HFLawy47gRejCtPzAAVdCnMefRr+yaBlAhAmcR7TLCyacs1FlSmOmJSWMM+8
dkPQGGH7jVUoHN24egmUuatjPhNf4EYtvsWUHi20UkiKrnhKWlNzNGJ6JXbNFTZKFpfV8Fzozlb5
Zu4V85I6a4B5dSpnxTAwQEWb3wdl7vWoFV2a/GlikiMUkJ0al9P+JV2gzy9Kk0/TF5kV8ltokLfx
PKnLh0/16m33cmzZmVvwnN1XtI/ad2vO3Eppv0Adcwlk0TyFFNZ7+bobg4C5wr8tJylPygBEPICq
JNI5Ee2G4tSWXMZRCZ2QMCKiIqUE/TWw944EQRncaUKoCtb1P4A81Z31tYqg7RIzGqx/gj7Tb3Lt
D/gJgPR5qjNqTWyTIpqJv5Q7vA8TuKuzVaGZp5nxedycMRuLcTfjjPtLytv84LRkE3FvndWApqij
vp7IPnk/8iRM9HYFEzwn64ctfUdJ1rc4qRW5mwpv7j83jjhsC6kZONHNqzgLUrtvDp2VovoAAI2h
3H60tfhgKsSHS5HcXBjcRZoERt5/swYojPZucK++uOU1mpDYRIHTxXxlhmGaebgZus3AOYXwl1I8
1YAvnrrTAIDFDc5lMsP8RMUaKGzaZpnbEls+mgURuxZqxfMTNVkq8eq9V03VRI10wyMyDJC+aVEu
SsOl9SJGHE2YdxWlVPNTsSp0T2xZW4HXo/ccL6YeB05/Q5uabS/F0e1dSjbRtUXRvJPSV86gDumq
jU9HwXkKfFhU9RVdoXkNFDqhovJdCAcfl8BC65CAUHX8Vjd77Jm8z28Uy7Gq6Af0FybWpd4RCfPD
Ck0NT7dEJd7NDj96A6HLyMEx/m6uegXGfziQ35geVA7KCJzx1jyAl9KgM7IVgJvaTdopuSNWA5hW
ADjpo04N0JlzOWvVD/fGJgj4ULtV9gMPYCXzEWWGfMbp3KdIZvXA2n86HiHGRCE6mUD7xUVJEEsU
uY2ZBF9tuc07dG1xBgGPs+wNJ2D31yLloDzBzVdmXPShSOU3cecrub4FWhzeo/2Tjq+L1swo9ohd
2ANb2DU5HzbjA9VCBGk9KYKIKo/WVMKLnVmvoGOWU9Hzfx8dvTMloAXFqg8ruk9a/kap+rv9dwmJ
90Vg647N/pYn4PIKCIjsQtdlHxOimmBvrC9VNHAbX+oU9mL27Dck+3KXPU+7Z+5+yeZP9BS08w7P
A4c73ZSNd94vynOfpmtktTvPq5pVz/oYBhe0WmScql7lbTHZ0eXww7qdBPzOD22rIVGWFGftMT9J
Y6VPxIrnSJgnmgHRmZKI93BFnJ3cuk8MVZ2vqVYa74ZQXki9w+b3pLLJTx8A3CDwZkZ3eBhHa1Js
M5UhS9XN9D895Yv+oS/SqR15AJEDtj7R8YzBZZusY4BeifzXpP/smLYSgJ2VyWuJGcPSHIqobLQ2
FeGEt+6fzWwZntGYRPFyZTqQ7+7ke9dtn8y5oUQoE5NH6BX7ByAAhBBUNtuUG5Y7qRtlJsmmLov1
5Tqv/9bCHr8CMrk65uVl1KHImQQ3FGy3Zv2o6M9IzFcIZ47B7czOTOgr/7RA5W2lhHbOlt0/CzhN
2s8t1cYdIKHjGDlm5SLcVysmwexndYaClzkopNiGAA2+8gVD10jxUak/DwFJct1lycvqrSpxapix
pcjqZ9oQq2j1r6k4wlDto1YnYASlwW4K8uAV5cltGJQcYvCnVgP3caagfaWGh8aErTesG6W7Z3sf
t9hFbCpYa3XDeu6850SRuqRdN5miKvoJ4yWTsf4EV3cElDp4JVMnL31rIQE3Urmq48K4UeRGrwqo
gCVOK43t9iNsZvylKQ5cn+vr8WbPzYNRkegAOoBNeZJwN6vLgIXWuglbmGT6/3rl/deC6s2XCQql
FOHOren+iq39YdUEqbEn2aIlQ4nPimRs0Z3R6L4c2438ajZVMBGuy73nZRqf67nT/RnD4YEHTcLm
bVe+WVNJ7HhSpCtMEuqEhl6KaxEcYexSBkkvlQo2EFSpIh2IUVZVaiipZWQQixps7QsXqxZqa4Up
dCJ7x2MLbjIMLTj9eja0J4OLgO8C/EN7Vql2560UtbAv4dD/QBslJS2OpAmAuWLsLY7iQ2A3zfrm
rxlHYDppg3zIfZ2yL5NrADR0q6YCQZ+iF66sgaUGzpR0nASmbC0rddCUujBy2ITh6clSK2L17W6t
zIVQa3t/bTvZ8Gz+mHgdI+zLQtcf/gl6yR/7MAndMQwJ2imiaz3I6U9nYsK2KiLquOsKvHGFUZne
EilPs9dH7QOid+pa6oyfHUUhb5Cs9vxcS0JZpkOLATQxIGh145v1GPwdPXEJlI8UDkT+o3LD3oZg
Z4WMWIFv36Z9oc/nyakhQC8e60xwxjfS75hJaVVHmflzMcLjUXEUW7wsHII4MW/6xv29Mb/FiDsL
0I5tnJRsqZVB5Uh461dqXTGS7ywoaTHKlktNgd3UPJh6kHc8J9bnsrYkYkZiwcgj7hXQeKMGZIN+
N0NfGkxbDk4O+C/NtQEHTNVUbxHGqsThcKyUEhOdJERSA+drwwko3vvs4NBfV+iOtwYagMikFqiU
5V90yAdkxD/B+QrcleHCjpHthK7PLXLmVgiRdCU8vTl7y7uoopmIX7iSu1lUgBGUm/PBkYBQRsiF
cqeRzlFwoLa80TCIBAm1AwZCVqMU2GdNMM96A75k8YwwQ38QFdGk75tCvomRG18GMleIjlTQdDkV
oltaFGVEBFJpBlZ3DOt3gEPnx5bJW5FOS60KHzvWkBl0TuqkdHjs1Sd2A+jJOmzWOCPst7YoTJgZ
k4kUbYaWUROwDJxGPgX/BkdG1cmTb1oBYa6i9ND+JCyYwYyKTqr1DBYxLirMT/vWO7IuqU25KZQv
OLL8UTSjWBCUm7llhHTCpGcdvESJufmJYw1cZRAim/JD+jPhexQSO9fgi8k10Qsinu1mbErdpK1I
E0nBkxX4ZX82OzYVMkuPsPauG9DlgN36Nsc2NGutNxp/M+VdR00qEZ5d1zyU377ZMn4dugLY3e+v
OuQ+A0g0quxyxxvUWw7kNWl0uwVEEw5THqJecRizpJsgyXXHLmXBVCXDsOxiwQ8keHUKYII/slYO
gBGPdpXPcuJPdcfnPOPuo64rDlhWkugWwUCYiHrzutpA+2s43FMpgLJYazhjpvsFlNgLUcWZnpf9
WpoS+qcr7NTQ73xoOaJUsS1n3qbHS49SsVucH0guosTnB9h0WyHvQaaEXpYOYYrDXBjAk8zb1h00
JJRjZ1Bp48Wc1Iz22XlJHDLhWLlqJ4DuBY1RlcA4K8HWb7FeSyzaD4juF8boV8OQzGcEzG8TU9iN
W1hiaTWdNbXfPIArJy3npfubCVchzJPrsgZ+J4ikE3oZGbvDhBfHyAEyTL+J3A+WFCH3D53u5wrS
x0IbTROerbkkgCFH1L5018boh3Jex8cRsVzWvi5wLKqFgFOEyQpPFw0PRiGJFEB21cMtVIeMsvtX
3R0vb08xPWgxZF00zlGl2Q5Nwyqy/2iwU8eQxof1q/8bTJ1nUG0YGOBx3EO0/2o3BIWRm+ymj48Q
RK2J6tEjj9YWC9FCCzBNVdP3sliIeP1u9KO6uLeSsWSygdHrSmUh2UWglwVDMBipDAepNQLIP7Xk
tB/6YAj39ugRnLZBm5UwtUCZgpUVDMDEmsAygRne046qB6KpWJu4K6TKWkxeefchvX2pbHsIrAmD
5mLk14m4W6ZOau0xUezJc7uS4EzWccQFLTyeuWaK3ZtA7I7c+mrKRV7jIsEpEgxpYteIlwZziF8e
ZbizeYpH9bMwZbP6W8rKh+UuUSAuzkv4m1HzTjhTQvFx+67iaoztdSowiWLeQzc+VjDSmurW/iun
ywNfE9qpiixPAnu+ilQCP9c3QgfPS0dkpD0cOKKhG5KBQS+s2vDxBqgGevXwBbubr7pzWsZhRlBs
2FlgRKJXCpiqkGsmk+68+ROegIhqKExS9KT+/7DMQsm1XNX9NF8xB0/Q9gyCzYdHdh3XPCWiia8P
ntxAOZdaR/392X32fvJ/UO9Tuj0dzbVCPKsbyP153fmAqrHpdiKpcZZVUjMYfdlDoJrQdZZGAnCp
hC1YHWeLtXJgPNwSjQcks/8AeONiQ1R3KXq4fEbux6z7TUTLBRZXjccqV1gqqedBs9+O5XvbrDR7
hhhABrwQJy7T+xHcAWlShtJkVpKUfo3aTm8zKO+8NeY25hspCK7SH2/To+qYLa7dIJ3vWx2mNzdx
X5WO3Le7KX03RzMfTdiPx5kWj4lzxvZntFU5SdpsEukVNDCvZ6ATuBDLUlfyebVrULk1pKgCdrGt
pYyObFjYeKBm0NVvIT8N4SNqNO9YJl0ghhqBEomf/E3DQBwYQehXf9J2F4c7IsrN+maWgDPO3CXk
xaaHNSVuds4maghJdq4vzkhWmi1OgMSIos8xnYYD4D973sq1C/+DneiZwxFAnFLfo3TU4rK27gIb
kx8YEjNPh5IPyZAKF81eDLDIfPFuPWFggmx4ablE87biXe0ax7qqP4AocZGKzoikv7d6Xj4q/DlV
1CI5h3opGILcaC7CwTUChkkiU0lFsbxQVHg+SqhlYSwnCS4eFZ/aQYhUdV8Z4ln8wwn+qsz6Ps6e
PK20RfuPcAejH27ALWFp6ssUcPQuIWf5UiMmF1u5K2bulut2eqCaoN3NQ6Mu7BFbWwCNrs09yIb7
X/6aQgcUsYAqDUiWOqjNlbqnItYWggQR1yB4EGdzNb3z8i0oFge9Ym21Bbx52xmmCzaQWqWgTkDA
EfhgCCTD9P+3j867843uGSS+HPDxz02NsjSyEYDLVpyuzrhlj1SuNu6ZSUirI7G2O1Z4ESB1B/ta
lIrN+68FIpRdqutU5qZUKR+JVpXp90Dmk1V6lthNHiUnK9WBHstrMpwukhM+xcPZ77Sm957k7Qmb
puaOIzDpgJJ6r6lEFvfkMwbiPq/M8gvMMwFz67xUFFSN8fJMtTcrk4JK8cl2UMK1nf5oJXHj2TMW
HYZRgfzCMq5hbe+7lkd3I5NlXIuf2WGWgReeFLin2DUGfTWqlx9dxFQ0GedcmJYM4IHjG0qKx9+A
2YLHPcLInEmw+ATimvU9OUOXf+G0LAINJmoI8zyr8YCOQAuFFRelhSVLP243kzTwwfjrWJnRjVZv
ewJ+LP+rAJ49n+SXUQi1J6ZEMhOiVKuhK0g/OU2Hx0V5yST4wnGMoRhiaTsLkoCpNtP1mjOYJnUf
F4CnCwSwx8y9KOV20ZcVSAZ+T6Gop4p2C9lEQsj2WY76kF0a1iVSAMxHBlE6S6h54MA6YdcJ6dSp
UdNeSv+UUr8mQCW5FYU5M/uxrVTCm9/fCUY4bKwlgKoO4hSgHic0Pas2ywTQ+wIXRFAhbDZZlGOG
jaIAvcpDwBAH5EJDsYVeLozLVcXs9V/msAmly91TwevJk1ognXTUJUfMJHIuS1fXi4rslJtHO1Mv
7vqlHiroZeulYNY4E9kFY8EmiMy2jc+lA+rK+xSUcW0DPAuNTAWKLXx0e4WyAayCwJJX9mTjMPYC
020kCDh/GiWogO7nTZKCXzg9qibVfqpTChxmvkyis7zVlYnBIMBgKM4dQMhbYNqFqXl4MqNgeDvw
NV70ki60ewYrJ4OqAp0tHEB9r2Yal5VvknBsVHjxAD0PAfeZ5k9xsMeewhwPINnLDiJ6a9OCFDvi
+CLDYlVkc2wM4PRvKcDtnwg3+K9YnO6as87zbUgQwGSqYC4aClrMOzdosFQiHN9+YFALDa8CcdGw
HbiW5OnFq5RxRng0CEywjCUCRiK6NuZp4dENaKHvM5BxQKjo0e4zrR4J6rU+4dX8ZPWIwUCkM8no
w0dTUen/9K2QeYwhggcvPoiIf7FUnifFYB/CZDpblR+3NBjdcyXIRcJM272gUz3duLjuJlNJnhCl
JgQ4VgkM8iAAT1AK/mR6lL5gDqzFhm99jNtnBBLA/5JJ2xWcH0jEetVpQxzFfaxRybKzl2iSErZV
sXW04ntH8wCnnHE0AsErbrjbChLDTtjsqBfFlPV9dHJL3OGU8rhz17rx0Kbmq5tzt182BEvgRnhQ
2oCluPAnMy+14xGmUYnSnAG7UyacmqR/1Bzf80NsITSzTgfnL2zz6rhttINTh53xXrxw/Y1WZb1B
p66sxgQjAeD6HTELkeex6eeuBstQgfn7ngspNtFJugZfeerzYtYvkxqo7T7Nxq+B9MrAgAos8HUG
HNJSTUo1xAZz/t8+t5AhWHneVSBEfxxlgqPf3ChVBBfPJAINcRbDVPW1hMnqbbAJvrGdCS7iFU2a
ZEijWyT9B/yhNIJj7VoO+YwYA4+8FS5GxNCS0Ty4m8dDQiUe86E4JBVEzTWnslKnD5uFd7G1Jo8O
C/gEUx+HwyESKf34uBXN8S/YzCbYq1XjEdSsnKZajumTRxnbazKc02U+iRNFA7t0CsOdxfYgSjvh
ehg4Tb7/jBtYSjcmmWqHgF1tTifh195cMTC6dj7vHF3JZ8ZK5jmS1l+Bo81+ruphErp8fFd2KIAX
MNEAYFoM9CJNhmfmsiN39KLM5SJKjIjn/NOO5qXeiQG+D89qkZaBCejk5KnMegvLYBLlmlJp9pv4
qgNlar4dbF4M4STDxyuohLf1dGaXdd1SD9WFggpSHcUKhr9i6g7MVNDnwLmk7ZIGGSOw0v+LfVTo
RVBP28g91qhYH7NDjJWVzxLfvOViyGEgHTErNey6MlwmAXtwtkw0AsNAspIS80HpYnRi9Qdm0KNm
CkedrMcqkDoKUSV4AmLRUAziU5Fako+CybsnvoqqJH8bF1ixUFpb3tEWjmwWmE4bb1BTO6CduD1A
bOcu1G27oZRKMa1Z2051VBK4XqsyqpIWtaIlvbCgeDOPBQOR7p4RZ6cDHw65FeGaWPE+TLjdxBu5
J+KY7uKFxRcwkALcWNc5W1W0yLOjbc2sB/Ym88OY+J3PIajqKBbiOLsDY398E6GP2bqrln6bGc8U
6TICoYWcEDK37za4GvQnCtoDzTgLvCzux9xrR6EiR3RDSn8NKH5OeFuoLILhk++Obz31BdqhnvE5
cwP1ByN2c0BwrUQxd8MBPph1JreTDy1gkXR2h9X+U2OS746/fT/z1N5vL0NpMAhHlfNI5GTfxH0z
7wGh3H9OElZC+TzIryelCBR0/ib53fTsC95PR2dduMrgv/9CUNERUpmlU8z45377jy4lnHro+stS
FZOfYJDn2FeNOmcm6IvkNxN9l4mabhCq1NaNFj/56nvfZCS7dbOFA3cUpWGLN/DJLeVdr88kQrI5
vMHuamR+v3rEB3hljyKSMPsQsRv4meaWidQw3t+py8Z0K1DUIzhqs5W15ynXTylrzH5KSTwR/lVx
dcmwFSXia3fml2P42dU7bQUlGzjbVHDZ82SVlZE0F0SzHLVVSshyZuT0HEbYksgjSzUw2H3a9gud
a33Qm8dA0Rp45hRDNt3meUTRzGz6thiHy7aPtBO4bpxhvnnsv6qncNVlRFd3YaaHeDdqLG+oqz3T
fggPbKzJswHvsGi+twOIygToyH4vDUbnUGDxa2uLA7XewmyvOQfI+SbCM3fwVyVZP8b/D8j3tFvD
Px7MlSFBc3QIehIEp+AwbUovRYIQ5JFXK2xAzh9lgb1GFbCAbuI0CGXHJobCVUVBKvKzqMln1Ee7
WlgbEbSvzGa1CVLrmZpp1Cj/JSQpa+f4LI4pWoXhflJt5p2l0WzhLLBh3FNA9Q/nbpf176nqtgJi
qcMgwtqmwXW0uAXaBfdfa34SFpgBt3jOZ7POkaqeSGOD03ZHjoJIzC/ztkSJGU8UqLLT6SRnwaBA
o26Xzo7GtGEUz24/+9EJ6CS9t/gI9B1V3CHXYITvXip+ff+j2s2oFTQo5VNc3bJlFFpsBWHjN7cd
AwXpVY7wvmB2jADywRRmoYahYngfLo+nyuP1Zi8825SkCXtKcPkboZweJ/hRKWGhYIfemT3UesOm
TzsAq4FtS8t+N5EVF/HR3fZ7H6b6Mtu5WKH4gFvJ3VI5HAa3cBpmrILCSb4eiJXjzKAHUOFxEY+b
t9poXiGNnyXvkR+al7WN3UPL/Cmq6Ja0DFICkkJZsFOTDFi2z4ZY7Yj2okzqHz/G200qpFjS+P6u
8tIssMuFEFA2GeFzIqGGe5531bajLXU7d23QdsFBlAVCaoU9XC3NTISUwVd69Nd8oRnGEMzT8ZIe
BCfXLiBtq7qpU2iXhxLeZ0LbX1x3NMz/P/EUarQyNLCEAtcHS3Vd8KHWr5vkepZmaBwhX0mNvbx+
gVTzyLTJZ2Q0fAQSPWWFnAwlX9oCaLoLP3Zs8kJvFLWY5XALqEm8DFBGuiAB6A2SqJHAka8OQXjU
8PT/BfM59BHoNq6dxPvJ2TeKfgeuUT+8rTcBF6r9UnkbowuMMVlzuVZztFbvDEg4RzcJSAB9Zi59
ZkRDXB9eT2n+7VvhvnfX9uBNEuejBKgSEYFuzcRnMT3S8+v+Po2M6gOLS8rTfIljOMOySyXnFXNQ
vsvQxsau50h3ypN7tJsuqcjcqZ2Pmqh/vGPmHrEKPN73Ef6cDp78Z5UWKvBwu2CgBnZDviO1eXkA
79R5rLTvL00uko1HzjGc3BGXOtBiyR8dwUnhHp9uf94H2zcKMOOq0N30NJB+OrKUdezflqt5eBib
uctIdYrUVkoaDUoO0JcyiEsj5CIwGgrQiDbNDDHxqGNk5gAMkZE9jlA9zb83SSfipUmsIx/avCoc
fUjpOFsOWXt6p3oCIjS8CGTYaip+FhUs/RwdpSGrNdhMBg8ARWqWabX4RuNByfNOTYogeD+WYNaX
GFrM4HysPTY0MU2L83bUhqjJv8Kc2lxf3TLdCoX+mFjshWtz8qaM6tuAxZPDs87i7cc0Z5e3uQ4W
/6X4jL68fdqUulYfmbwGYoDEdqAC3zuuNr3Az5v9chr+lAbTxL1HF0/JVmCCneIwxhN1bdHgLUpP
ujK00ujc1Zz5NP8jOMaOxIaoNg0uXFo/rIJkgRzKCcWfah+lVMpZXDwInawF+Ee1qCjlxH4Tk0ph
5c6Lojiw77/rDua3m0mLgM5V6orVdIaw5PMZ3a3msRHp8/7051QKo969KNWCVD9U12dEg9hHxxcm
UhfDpcXjDAf4VD2WBkl3yNwLPZgJfvut4MueOVNa4sCB5a1zKlnDabE2sxtQRTx7SwtsxfuDrfd9
k0FVHjwc7X8c2m7ZLJe64nyPValnCFdhi1lWd2KOyVfp9K5gLtQCGMavWPWhT/DUqQn40sn+JEpS
sHJi/SO8GS5+jTVf8zWJp7Y3whnsoldYR/qZQl9Mbj6DmqY1/1Ps/SMngN818QAH2002VafQA6Qp
IkLrI2W0EQqTgKg/b2vYeF+sXwOhzWsgUK5GiO70lFZonhvs7+FxtJG93dh0NAxfdgQiGM5oWTAJ
D81YSUpUYBbwGfMhqZYA8ZAyeHG6PsNmjrLoq5J4D0aGARI3wi8USDyD9xmA/bYXphJXpcyyAOI0
mO62EAMcEUzFlTTA2icqWU2JsTv9XdR4K8JS6ZSLPE5lgzia3r/CZOmb6YYb6DWzohod1VMtaKlK
oRbokbofSu/05b3Qmtr3pByraaZQ1X0B4tor8SBdEaHoHqEr2nv+r5D86A5Y3NI7CykW/Aw2QLGG
mG9TBSvcw6X2SLO0XTSscGtCqRTTOseuj+XvBGkehvwjMcM7az2xG4aUM0YViTvOyA9957LVkdK9
Ak2lG0w3Vxo2PWEFxVOFIoXjiNunQOApKtejCsb6ncJLYOT+0GVkJKYAXem41m7DU4QpDGOElcoH
LUDdwF1KoC9BPbUybwa7ZAh9t4EwwzG6ZUsDFrU1/1SEnhYjdnZYAmdRdTWEAqPe7jmdLyX4syXJ
iSE5dK38rRvYfBKpMfEgBgTWbfv9s7BqvNHfVfymYIpKnfTm8uJ0SfRRpqxXOWmq5a1FGxKq56BG
28tKykkHVMmDdci+ZBqDwRemH8Lj79O+7NbHKTW2FTueaQPW29ihdO8S/B50t6MyHe0yXzszjwFH
mpyTTPHOibck0epJk2YEhr29PDuJ0sNnrdn+Kjmv5B2qqGi2rMm7oH1tuMlKMIR6NiuJyGTT3XyD
FbYbvh8fe3sJJuupJbJ7K201bh4xUKa5ZYCjkbbMdtZS/kKwemjZYSL/994C5UeKUQAc3fBEzqLa
HlOVL8TwihxVyGfPPinWSTuISxwkQBUdI0/sd+TYgbIUebFYnpT8iypHyKc318fAsTizwMaLoo62
bL9RrbAFzM+s+WaC8kVuyOpAB7qGSnK9z8i4BLgdEzoV83T3gQLmeeyhAqWYV7PwSmb7ourW7zL2
acIWchyHUUOCAfxMoAyVfsQcKhkirViQ+Qy1LitIfpGXqIAkXUqYMo0Yypc/3jaEsbM2uXzgT6gr
kxTXYyNmnfKQ7LKwHp2W9XTl4ljY68/cUhEQSlEIs/YoHfVVLpl+klYYKONmybI/mr80yWtrQ2yG
KIqFjjrKcP7oZyT3ZO9048qRF7GNoKZuNmkoR/Zr9mTl5rKNWq1uneOJaDVyG4TXWear7pWal5+Z
bYlrGIhqW3SYOvadsKV2r3MU0+O7LfhNw+aDJxAvNhz9q9ONiaVdiIpg6TRV9coh82ctknYdPFdf
mMWUnqwnrQCaGCAdIrSBMjPXpGIePzP1JtSSWOpB6IkuVu4R6QKPeur/vCR4WIRYFIthi4YkdWbl
pAKGOpvdSbGhiAG4O7MX35NxWE8Pf0CPxeqSnrmjbrcXGyIKh1HhJ1WVbkSB58tftDszPqLjw3Mb
SzMMC0gwa5ynmkYrai170l6cHd03ef7WCSPUcD4upfe4rlopkTfEiwiav8P/cmgNj6J25URDl9qv
I63MKhdOf+2p6vIt4BFO3CIF0gEGVnPMtkiKG46Wo6TNf6Gil8/WCRC4ig9yu8KeaWrB5bngX9dt
XE2/ig9ao1VoBUaFXGsQqA7/YW/7rAU37Aphe9BShlSDqfWIlci8rBIDycuXdLJRaUyQ50N2gh+Z
VMI+SZXr0K7+NWpSIQtQE0iDSwAordN8WklajWgNRzKnEeQXBgtlAnCEFvfD/F+tVvH2CGbDDCVw
xTRsSFiUSf3rtN3djf7z8+hmOIVseivwG+QdiX8rWwjVK5sTYv/arRnenTybe/Pp6vP2/onuL1dP
goh1VQ+HRlP/tk/OwkXgdOXhiEoAzZ9bmIHDRK+l78HilNuH++lC4hRepRcLqyEp4HgFkMQ67yOn
leEbzLffuNAnIRh9qutrQHY8vZobfq3AjItMTO7owsFE+jkeN6ceFy9PKAXgeiFOs0KDhfimvP28
p0qynf2ExKcK/TGSocwFAdUxhHXL3EiZiPFuLN1TIu/xC6mAFcqCp3mnfX8+MUGMVlw4AgDRTcRN
dld5qi4O8GYgGbPxZ6SkezkCUVWD1WjxbhVcy+aDcIHBgTeoDqiPV9avxDDAZxG5I7zz2zKNruc3
rzQjCsA7n/K7zs7z/71ziGjR9pkqzNPyPS/l927yYfK5NJIkXZti8G3p389t9sVTOpxIOsZ4Bly7
tP5x2UE3p6XNYC4g5B6ZUxFH29bZfKgFoVA6n2rRHu7HJ0/exOP1WDeK1UW22JLIjXphsqkFLqqa
UXMLd6S43nK6Zld6CaukBoDRbXKRzorePumuBTvXWOQQM7aXJxDO5d188dwyvWfboqwXspVckPvs
U/tsGknVKNBqB4OxCqD75+LzHFjoc1aX3FziH202F4c1F0cP7I+BtNVv5rNfVrnETvcHwqYbotvm
TrcyOgueovmtBk/RENxDP0eMrAyHNmUwjJh0et3hOUE6++sPYNW9HDjs2sax6S/blVJykGo8adtT
vqiGCVbTJl583OeptcYwWeJVUzEmQRpIYDJX+9shWbCVfNiaTSwo5kFn2ZUm8oZ6h9eN7UJp2vnT
2iOVf0DsWWckNSoI6EkRrdDE9yHQvb0bVhfdD6/3Po4cEfJ/xBR8RBAboC+gHvJ3VveDHXmCpQK1
IHNjbXzYI1TYc7bZlz9WqHIbblJSyKq0optoXwb5HtjLQOvqcJbFyrlbbGlwyBuw0lnj6RAiEsI3
o/Rk7CpkVoNwnKrJBfSlJ9uuT69SVJur85V3w0NdOmPykCXLz8l+7ldw7gdePmPu/utBR5UArxAP
wwkxY5vbD6/6VrLkP3ZrB7ApR1rOA+GqZk31Tq6TjsC07EaCP8j3M8l3vwN9oeGFrrfsV7k3eG6C
VKk50TMr9cNnRx+CerRnXClPLOIydd0yZUVEBmyLND0/B4Ee09b/xPIyEmbd5R67T5YMtWWOrtHL
L8vt4YtI3J0OzTrfc50xPjO1HIG+QHX4HAMpMFtrTLMY7uniyYvt4r5x8/ahsB0nGBMesJ020s84
noXWarMkrH2cStnc0D+/NsWTg9aNQ2uV+Fiy9wvrIByeuZiSrqSaj0gUazsOVjA+X1bWCYd92SaY
BFFaC77n4dlwhH6/5ysxI+t1r7GxUPngTirdQ6aq/zp78ZJ6qOiHTZ6lUOekVw7+Ov0xv2qEyM35
RKzIORzU5QO1BpHpID4SDk86C+bwRQzyhFj8f+GKQlQZAJf73X49mrJf1B6+H2gbk1xACP4lEwYI
IZZP4DyenEtdpjx7G1+wFiftAW/yGgHyvVTaU2G6klivfAHKWlO+7hzJZjf25/Klp2UczJ4rVKbN
gl/11ncL/rIMa9LF+ZgTb6H8EVCqkrxBgcAUSV6BXjJqocXV+oeq+ThZ0/jzMBpu6RnwO8Cw7tCo
OTmw6NsT3uG0gW8+i265hnFM1wSaOU+/HGySxoick+V+LoxJQpzf5swiVObAx5pkH+x8cDoFNIal
Iv/8yvPcCfXU4tHsnqNJ1OkQykRV6lGeWVVH9jxsR1sqTU6FcrS32vbG0am/urtWGzsp4fG4/F9h
eYHJkZSKjuQ7uDS4qoy/5kvc6x5iqNsbgpl1AjvDvPT03LaNa6STD8wGFtjJMcuM9zoBC9lNq2XJ
LLlbHD8VOHdmWzwwBTfjzXUmP989Vg+O2duqxuKMiUr5gPOD6VcM21iPcFBrydsKCwjOxg0EBFHg
XnZ7JBnz0e49qX995qGuVZawsoL9C3s/RSq/XN3Nq8ytZXvyKdaX9XcmN30vJWoClKQpAMrHT1V5
sdjw58E5GnnMBnC3CM41a9OIJEOLHOdJh87qvMBUGjh4Hhsc9yVEVINqtZq7QHKOhasrDIkLlSxO
5LW8ks2cO9EfjvPTLKq3vvcmR8rBbGyJtDt4G+OpOIgurcPL7WjNFiBkjZLnzGgY/Ff54SLIgLiK
I4c5o3iDsHz/8HHcOjjLBg1CHkR04+Zzp/R+8XSfVWN0kOiaUbVKEa1S3OL+29eR1ndCZS2D9ywM
UbEAn1EcHlbHSmzcqjCvIh2TbeXiVzigjYHlT+MrlS+uR2kDsLQPVLqpKE8M1xQd3J/zW7ST0FLV
YnSM8JUaiDFo3sO7iQ3eldgNXh+g5KkW+FKC+81H9Ll+RkJ6b4w/6izam/yolLK+7EnTIhxiy9go
3/BgicbxdHyG0RgHS5mf97bvWgWePKHQMF19RkKp0q2nL4UOo6Hbhj3/WtGdRc9ppnIxikPc/PZM
7Q3QhkWZhosTnzWKOQgtUJbbp1dYsV9tk8EjJaRSldctdgrsu223iQhOw4e1HoXW6D5qa8PiewbQ
uAQR+oQpi7jBzm56pGb+KUljzYr6R0NT42EKMh3iRrxXo/2fWCVbiw5FV0JHlBRLIyPkHgdLKW/j
KXLw7OnCHTZCypvkHPVyvQiaytDtOo1kLesFpotopPKvpAcSNgH19546odZs93b25y6mmAual1k9
uAMXL1MByyMDQqORum0sTtSGZ7bl+V180r9p7TdOsdbAofHUOz/e0FoJm+E0/VcAFoo+4MqTnPwp
6pvBtthFchZy3W+37Jc3HIOkrdCa//SLVMj+sTWq6FnRcq1K24TFQsEqE4+Hz+4AiCzWQnk+61Nn
9Oa8ICs7UGFu++cuA5WeVSIMMsNivSfWTU9057sUkwV3qMuMQ9prWkYQsuZThUn4MORnrPxUJQn0
BEX52ZJPA4BizwN5Yx09UDDmNgOJ9RwrfGjlZvj0Y8B0IMFGMBMD3XgAmBzVTLKSxjayk891eGFC
9MLRWq8CixbYQMiTqrVu7DfKxHHlBoGeY12CTD720yQIjKbf/0Q4Yj5fOnWRXGnY3Rn5Ev/UspJM
9Uqt31K3B2n/LkhDzZzy3cqfSrgO9gMgJ8sloHeeqvCwrLovY+fXqIyVQLkCB6y11Lh4/i50K95s
17lZRxLXywu1k42BFCvtoSD2W1cNXQExlIA4jJC4pJ9RjjXm94mRcZ5EcbOvYi1Rf7b/sSnemkxG
hd8Tz+8eSO8XHCdacdEzUsLVIsgPBK82s8E5Kzl29ysEzK1wmi0czRugqY3MQHhaw5CF8z3nn3At
ZKe0E9U26dvDNKyUbxSKinMIlFvSrNt3uMEOX/py74wYINO7GLsf4epRK6lsVmDGf3OCfX+Juw/K
owapV9xU8JoiGhsIR2ys3ofzYW7r4Mc2iEfRSX6wePtcLxwmXhMX5U+5jESLy6NBmXMAHyuR/6dn
QtsHheb9wdqkwDOhhMaWxUKwGSyLtSehug/SiyRqamt/T1hG1qjhRo2ZGJO6R1Og3ddp5MoaRXBw
pRYSwmE2tjvl8wRVlQpc/G7lQeryGqMQ+kg9hTzZSMDW/NiRAFBp9D4wuOFoSpWlnTUtiaGsiDGg
bG3+UaFkcOvEOIfYESn+g3vE+wPem3IoLR2xVichlpWAE766D3pk5mVi2nTMNACjfRGTqlhEcBZ1
cSX3jdJeTt4UMdIVyHpDFdb+mOVdWg5FWj2S2MMcJY7IPsPB7il3DX+IXJD2e8aaZMejqv4U7Xbm
dDYXRhf1bDkGMvgkzPXJ5ZGad4GTox5J+UTR/vzjz5Ix5Gl4itAbWMdj2nNr19uLtJNk60QXQrsI
FSnsvOgS3buB+DQ1fXDcNquWqnohr7T5BEUvBgAjqHl+6hSEisFDObZ+FlDoSQj4E7y2raSasCXR
s/U5qul+d7DYo3LuFrDjn3LAc2WuKhqisAdNkTxRSmEklQlihYGIz7NH0+4/togWWP9WAyTzTNg0
qonZkeUjLZnlFEoNdGUY76yEYgIquqteQXFMTup+d8L4JeSHuztvQZSw931Ets3oRnHfFzz3qGvQ
ZcGgcH0WYbd/ZqX+GryIYC85L1KzVYMF5lno3MRDIP2fqnXOP+2CyQN+cOU4fiAGMFV5brYzkv67
gKti5gnCzqBUI911asOgWCICRzjCvW3F5b84k32PIn92w9qA5jRJvaj/gjcuN3O/EaosT/bYcUir
NTp8Mrx+ccqmJcVDQ2/4lQhtRH45LNNrNP5VPLfr2OMTubbHQ0A+YWd4h6hMKO+pKWCBbKej1VUL
hqN5h3GJrcNjrGqxbYd731GOgkitWhhivUmwmY5/1LPOBPKZbZk3NErbZIGMVtrCpMy6E1yuEEJs
Lhen+R+eRvqHbVp9SwT9LFddki2MJjbINftQ/6lg7tKl9hmghJ9I//zGSLmFJPf7IMWf/sHGCsZ+
KOx+o/DIQ5EOE1i4TjQ6TixSjVAWNX/lUUy2c1F7cSiFAO7uPE0+bVcr2AnZ0XTovGNVL6iB5ySW
ahfcaAdbUN5Eig/cRjSoFYdhCuHhvGoIJpSdLy/xNiFkWwHGlHaBCRPQPjuYl/Gyo+/wGmP8ypJo
R1R2mtFfXdQ0nGqfxS8iWo4jvtb7Bl74x4jFoOpg4Z1ypX9SHtW9nVzdM/vxwXsNZOyBfeSUPzxE
KMS7o25b2bGrDsMbbXuXvxb7C3A8SL/2pUH0REwoqDGHZifBwa/RZfhHKsYIBKVsu6oFKm9AHSCU
2wdLRub2X2wOWxAdH6X9G9oLr02+qJXqcqK4iqUg79z/g8tXeRnTMlAA1m6Mk8U1kQmEh/g78dDn
KF3agpWH7w/7NqI0h3nhvTUCgX6KJC2Lcz055kQ285RMfH8M+wE0OMEftams3wvVpVXiDM6bY+q+
dmiR7GwwaxfvYrQwBq8S4uVFPqrZ6zvj/3g8/G0727cOQpbXesK3/fXWPwqrgBbIRB3lGgxvwIri
/XwCgC05mJE+5MIFea3phQH+lOVvkE5x+3IPcxxvcipUNwgDEAwAGlT3Ale6dvD1IdHXwfe3JmUM
h88LY6nE/wgZPJqB9S52pmG8+5KGj34FWzqUIOl3Q0WFA2dWaOh1gvt45qn9iEIl6RosfAT86lI2
ECA6KLCl1D7fwUpj2WtGBVjtNh+erJnMO1kjm1pe/n9kP0zeU/m5GcdDAo6HIgqOsKaeFGXc5UIL
9qq5ODbkRaQN4WbPqFKoDS9Y9Jj5CpGmk+2Ty4Hy0bgzrkpGy/XJkB9GJa5rlKkMoHlgFLGli1F7
5nIS4ILXYMVHpA7JHlBoX0k9nMEy1rzixSs7x0UZEIKrEMb8CX4zg0TeHFYNvpscPdIr/q/yd+Xd
Vk9kA2di/FehNf719jMCep1PKNWIUUGuzh4VoGLS6Idl6+hXF3lp2rxddTjbX5/Vxc6yGhgF4MO8
uaUxnQdYVYmA3UtDCLRsN/8HXIB3Z6s2DLn0mofdaNvrbyaWqYvh+CvguHk1CvzthRojBdy6z71K
ce4aZ6HLWavBmzIp7PrEH1BWYtis1Y/6DEyBtwrdYLxQHBq7er37uJHuOOjQ/T+wPcar6JdFuwqS
3am3MUczsGARGuffENcdj5LQxVQRqRnLqRUR2OnIb6c0sy+/jer2OzuXA7bPIKLojjsYSTihXnCL
8+qFowpNkQLU/qKVyecv7vpGEK/2pLeJ9bYTrRhPrifOdrunmUZJ+SaXB0onS+c3ABTnyc+L0/YB
k8FhKPHnnvOa8fPiXbMu5uRc8KKSfVQDoNMticNxJ02cbekJ/6iJyAzIe2vaQE2mBQVc0J8C7Sse
zXRsS0R2GkxVq8oZs2xv/wPk/FDkAkPL7KB3TfJu7aGlS8XkXCBbjyALuiYAItY/vKN/MVnVM345
9x8EAuBfBfFB59GHIsu3WDwuI8V41QDvn6os5caTdj0F5DS485R9KGN0G7JlkGRHpVVzmhqKldqt
byu6R4uIUNoWLMfTsC7JWm/xD87oGMqsyy39p7ZnDeLGgz9kXs2p2nEDQPBLojlaHfB6eNt6SacD
DJXtINfsGluwK9094eOjIulP7mI2YnB/Z1FlE6HzSwuQ4NLr0Yeu+dQ9XNpDfZcMt1FdngCEM+Hc
Q6BV99yfK58AdfRoMWkkS6+JSN7mpjlBdu+dJQd+3Zgf/kxk62in73eMpYHwbuabg2HF9Q3TDDPf
0nXrxr12wmiFaOPo9O9BWHRWdZGRP6TaWyZbXksSvUoe8JsbK3Z1rogbZuKvZVSGNgNhcAMd5wZe
zE9Ci8IDGrLfEETaNC+l5nRyRaTPi2SNvztCSE/MpU7HdpgBxPDWh0LMm/L33T7z05CVrA9O0ALr
u7CywnPTJ/05Xo29l5JZUYCWsvVUvf2rR/IJiONFWR71KDPMkYz/fzO0CxS5UutZo7ET0AylZVPa
eEY/d0xl7biXIT4pneofGtkik6NFyDGOn1xtG0SXzJwJof5RDVz/NR8kEX9PO5Soc7GGNhofgvzw
pXd/JcrTrBaAU2SJLq/2bKHbNaNwgT4cZl+pJZjh2Xkk7qOSAsB2FauthBhLmhyn1EqkHU6o+UdE
5NvHYtrQDogAVMvSlyG+Oz3Lpew4KJ78ZKunafuOD2p3zQ97J/yZjx08rn6ceFLzjEAlwBs+IoW6
72eugZjYKpkD/DYe15FmkCgAyv4YvoW/10J38pXqwBz/R2KBfAVCpcIndgv8ZqIKTJwpmfKJrkYn
5pKlue2nZHwqIguRO1JPSR7RpM0CQJk4U6Ag3RdNyE+cPU2+gGaNYDiSbnsCQi3FYp162e1RgUSd
6TsaaxKI/rP+uv0M7WZIrRX80R2zAFYUE4sXRk0a8iAf4JFedfsRVYHBE/Ie3uPk0ZIbuMEH7qzF
Hse7vldE6tHQnxLd8917NfN5eV6mYw/J2FcrW09p4HxMKe0smiymYjTSJ/k4HbBpQv5YfOk+S6n4
bBZsMvVz/W0QLl2i2nAZJCxPfmRZMWZcX85pN39EksSkrJuP05I+lXJ5Ey/VWTbJ8r625ut3oU2p
AsoC6O02V+7QfhBLos/0TlqdsB33oLfg5N7U8HczVfSujdaTBt3LK9iKkSwnKBuhi4xbM2kiBsst
+awu3vzgRDfBOHK10r3cHbAzLdf0GxJbsrnoZV8RnIgyzBL13v9OU/I82tmRVKJvS97M51ZAAXme
PLfsG+H6Yqkv3xcrt2WY9NWPO1cJ2SC/A35OsLmGodDDFPfLReKEE+jPSiqGWD4y9bHvS2t4AnQz
/zKsFZ5qJkeVHK+OvkLLbdK4oevnFnUizaF18JH5l8oxHy/LXBBEr8OJKB13S7NXiWxIMGZaS7PJ
J8LaZ27ZLD17k4dVPJnNZwvdf25jBZ/CseG0sB1rpccBDC+K1y7fusRuWSvSigzqBvmclIMyzt6c
vquNUyB7iLE13ewDbitrSqkf1OywicHu3DByTmWoyO1tCPzxUcSA9sttXdkYgO6rNNf96N1Xhd0Y
f5XozoAIPj2ONakBsDaVyO2cuSTqNzp2U3nGofegPD1DXLgZKQujNqMn89yqAR6sEOO9qHgdqMMF
MwMSRF/NI4911PnFJ0VtSpZTrxU55/K9Y3UTVmc0tYEuSOcYWhPCr34tT3KehtFmEaDiJEKi28Bu
A1F4Dv/lPRIWI4UIunQe3B4t7cD2jj02wdQSxcnCxw+8PK+QILRhTp/Lhcz65zEpXGZz3WiaUS8a
6M24brmpOCgK1CIil2RK+WBd8AdbI6M8hcn5w7pth0rMdPV6CfJRWEPNdHki08dEaOETJttdQmYu
uYoOfcATGhMHYLlTGy+NsRe2tRDSXHLDxF7R3q4UDinJF/+DV9Ya/ayrDs7bA6cQoJxpvIsuCUtE
mbsDVeMNdMIbOvQTFFYGRPsgSWCUCAIWsUkLSRRzkJnO0JQSwNheLdsrk7xSgz3bDk0fugVMlaMW
NpWyKIl2d4hnnU/Lp3Jz9HjFc17MI5OoTYbo3yi3pWLfVHEO8H2hhq/+Y4/6uOGBIaJfSEGLSlIc
BVOdRGftFEDOVe9xaFZ/M8ZFo+gM+MD5bsviVoTPeH4x5tK3fQALLUj5BoU8cPaDzlRXTIIdeY3t
Oj3PhrjuM/NBKg77p70Eiw2x87N0i+Sf4iUQrNblc8D8U6W/dYOrxnsfaKRqGrTWb+MpLc3cT9W1
gLzeYmOuB2E7O58HwpFz/QBQbCnXRoJm6mA9/dMkVsri8+NqIftTqjWt2gjzADvfhLoFyWOGj9Be
k028Yh/aNUS5dLub8mY0DquKrGbbGjJvrZ6V5rgyicPQP3krKXaJNkEmG4Ro0yh61OspBMnjIglT
gJNCfahFN5jdP+YNMjk6stbdCwLSQ7/yEvTIJNbip4+0g17iP+6uWBdD+n0qe/SAG5J0Vvf4ySma
cYijpBtPQ/3UzRW0Peb9LKB5evmYHZPJpMeaLf2tUWb8ORfYW0a341mQMvOtwIcOyJocmxnDYlm3
Vq8ttGVEQT2Usmy+86PJHGJmhmgPIQzYpy9ZmNbx2egJYD0GWM5xo8ZmpX81nL3OL8EoXxlncwLn
6nioqMj8nztb6uy5g6o3EOrjc5GHzYXJT1/0upZnWgAXpMgwTxf9oLVGqdPvxykXQInJiEl/Uk3z
3tH3wB2KPsKfEC3b1f0lHdafEdUyvxP+nFhZZa61ol9AVCroOJ8A/KFtAZN3iGoUqZcljJWAUxC4
bwSKPhLVtHbhO4zgNaKmBNkYcXClaKxHDY/kqtDHJdzHkz5y0XqG2sBUyGnkwpGb2C9Y2fInku5t
rENcPbXj/qO5b/MdafxpJpUwsi9VHrObuGMMS3kxPO8XIPbnCHt1uhAyWmXejVzkp7pGId6JPWnY
o4MKIrf+tLRttzsWU+nNW0c1tjOEQ1ccs9FhdNJaGD7oaT/8ShZ4ZzlBerdyuX3+sO6RnrNeYQmW
rg1zSt0q/Da17wpWKI5OOcO6J44xXLzQCP6eEZF94yKyceD0dR5qN7l3u2rX6rglFNQYywQ4YsnL
sbg7ctD99XIkWrJFkcZKQHVtL3uKau9IcRNjTt7mNxCDqTIe/nSFMEygeCqNxmyaDgy4TqavNAal
UL9Vy80USX/ZfWiwJ+7xaOV0NN7GtN+jD85l3ZyDA0/9lDU0TJ6sNLU4z40dVT8XCfytXh1VDco8
mO4FPEDB1+t+RYidpDKv/ig/rmFigSZfde9oGPrlQjmXhEV6zXGkBXw/JKMP/I0R6iLU+E/ELWk8
gZBoi9cPqYgU+MFiloAVNJQN4ZhyTudQ3FwfuY5v6nEm8isTButDmZXm/hP92ACyUyvsrzf9+UNk
HDEqp+Ufu1UziQt65BPIcIp6Dx29N2HcxKQMxI6HRF5/2d9h7uGPEgK9gsNibA+DjoE+iEFhKii1
KX3+I9kLikchJoy0viR+IIdte/M8m/OykabM0wwS5jRm2HgrhIxwna2GcsA4WSPzO0F3iPek9soI
L1NdP5bOCfg7v9Xr0vgEMrdQFabsGeVytxW7O08ySXTXVC7ueMyi/4draPqW535LKs+CX8zPenIG
My0gM7Yh6afjOxX+LUDNOlfOgtJ5ftT5Y2OaK+r6qS5XqP40i3oTk8s5cIs30buBUVSxG7nKY7+J
f9ox1UWDU0ubxX28g111/QDROauT290B1ya06mK49ehz093OIhPlziI3cTWA78HXNAnj9YTneRSb
EEBiJO7XWSueyhavlc9KYoq8icRVuRHQ85DHBKIsE8Mo6SQbBorBUxt9MyyZTMScfNhRtZUzJm+V
KgjaQ4NzILyRa5Y5/a8KsdYHxLQh7LQ+nJgNGn5BHMnSe6Mg+A8aEaY9jPoWLvqe8pcarTJ2gx/f
xICfwFf7N1OdnvNFHRjmagjau/V6NrsEiVZaR4CQf71ZifkGpYiRpgt0oguenUxD7Fo/EfvAllVM
6utYpTgzUfClIo88dqtKi4KaRwyjZtJtCdDCON4bvCbXWjIlVoegxqIj9XCz3DnOrfkL8FeDZmJu
LMfvZI7ZBzdaIHfz4xbH4MZwCOCLw+uTxgBiOSnKS+wiMHK3ljGpWHRahGfZIgTguV5GYc5eYp77
J/sKHWWPDWDmmDan+9llkLx61I2uB4awoMlThZqA1AsfVT67DZ1sgE/SApTxuneOv9dII5cl7zh0
2b16sKWG3v+lwkzaMdblvFXqKvAE+YZfDPMoytGJKS2VAI/vzu9tIXyVD/oqonc7Uf3x+r4LKVzP
AzbfOv14+p6Cm96OEi63EM892YaHoYTrZQYNzPwVqsQz6qn9DE1uWXS38jG6ab3+mWKvEdlGHMvi
rXJFsiaGRZxgCd3kWTkODSbE4T+KEnjiJnMXLjqRRpRbiLDqDjT1dtuLq/NSZNtCY08YGy+WYGlV
/wIIHvsyW3MgW8A1e9ulxYSLNnQIwzvuSy4HS3bQaJb5MBRJXsCSRSqr9wqSSQNDxIQ9Wf2tH7uM
MjorRxD5IK/XFxIKTl7doFrRJG7KwAqRDVU078aqtOMlEE/EltLl2l4qBVfDdOteULmpjTZ8uj4r
YKhjv4rdZL20rNAqiiZgoP5vNbuuRCYflho4Q5kH02qAkb7hOEESAeId+91b5tl5c3NIscITmIvp
8MlpWZSVuVSDrqtn1iwMGSj1JT+DyHpIJn0tTXrAUJUhCcpKRAgntAqjDLxoBnNFam0+lFhFbwo6
u9WYJDZD/fSiBa2TD/ijG/4gKYeMh1FJA+VyNbg3VKuxuvwT6QPo2yLEdckFfCbCZ+9Yt0dQp1/9
e1LnfJFrH7Lfu+zkhrYmA+HFDRe0svnkMweO5g4bywvNMqa0eOk5ppUBieIaGG1ZCPJWiRWOJDZO
JtK2ne//mvGoIt5Zo3DRn6H4PQz1kRrUFKAZtJ/gZoK8bomzVP5/g9avmMpEO9V0Fo6xiceQcwOu
q78rFrsbLsGcbOUCVdjR+2IuHrTo72FkTN+lWnq7KQRzsMiuN2Sti0huebavxKAj0pjxQK8U28H/
vvAwkMRwdbeFS7/w3q8RSbZgxqn+S/OjOyK4dTttsRtd6M+YTHz3M8Vl+aI/Byp8HSbUSnj34xdX
51j6etxGV0OSolBrpH4kIARIKveWgh08oEzbYlsni4jqsTHaEFLB3ItUtGrMBa7PRjD5c44myA7D
a4T76rNL2gdFYKGRtbJF1uGMQ7R/kqnd2DDdLDwJtPaKGRqHLnAK/aoOBL6A+ur7CuScfVOYtGxZ
8SWF8W28oiFitTjLKn6+0amE7XRG0vRCVqUh3IBRXUsycZambDhqfA8qqgMbqpoJGv88SnM5Lv5j
NtvbaSkDAjolPa8WwWmfFYYI7zIrqb7SOiLrPhFvu7hVERqcc9yxl9CN3MaR6RHgQjon4FUb6cpM
DKDXYuF90OirrYnB7/zYs2k67KPpdQTNleTcZb97NinJuafVSVjM1WsD922UhFAwCOYGLaxJhDvr
0zXZ7MRhUQAG75n1E9D10Zm9qpBtBDecf/IyCLIiiCXpjVo4FaytO3hlGxMewgHenDnJ6GW7QsSM
G/4BheE+sC26rCckn8exBCyUREL4TdQaJfB1oIrsLHK3kb3xPTCC4HqMukYl9nZFNFmz0bJ4n8ud
UodI+SYeNIY0ngegXo/AE7kcsfx9H7ksw2KyjusmO457xQczLOm/QUcsGlvTa2eebS90K8ZVFwMR
jDmgxPqtMRy8noaZvT2ujpvr6CzQ8qzKLAaTYVo/bSC5sQgCnH7kIU7SNUWVui01W5JtxQqrj+tk
17avgmRVlCMXxsXszAVkW+OnVY6KMTtizHJsjQgQCC15kTbL/iWpWcGc2CjtFZdVaB0OiIuo0vJX
C/iK7k2CQ/bVSJaZvPORH+Tpy5cCDl3T3oblh69NCQIVE1RzuuaFsAX1eXpqkxdm6+OwGNLPzhlv
U7QEhl3YWrV7E06+nx1+taFBj6vNycePyZO5yHeQS9HXGaIm47rI7K+kR3IgvCgCwFWfP9v29Plj
bUoNLTUOxoZ8d4/i9sCT62zKD08QQb9pDpxyEMxmap57R+53N4uUWgzGGLiZEALlVDbfsuMRz/iu
h6GL9/DNyUyJMg+TmX9E/PJiUCDUiT949xtLJQVWC8ogxmFv4i6HY0cSkXa1w3DWYpgGAXWsofnR
Dkg7sFpVhRpEHMc3dlsGHuO3LNRVT5QohIUpvgLw/a4EAoFZ5LNNbEwDoyHlOt+Dyfjp2cSK2CXt
H6mnrb1/kW9bv7FgaS+3kwbpucLy5JJbvJZmXnR0Z9RAW13LV8LkH7Lfn4ZTemqIB6z89brVqh0B
nlir+KQfIiaTA25VRHmUVWiCYLkp0waFyBjfzGjBZCf5VWCbOCHxI5yzTjTEp837WWA4xNPkXM1O
Y97w6Wbu34+vnYMwwSRmqW+7GDHkANXvYDTyCXs+QGGe8tBkJbRQIAiIzRAJYgUpAUOLb93QUyIe
66eQkQAkgyRpd3iLNVWs8Lo9sF+OwohzIjJaqcNxceBEm/yCjnuHwGz1wBOJnT/ijZ/O8KpbitO5
nOoGsH0m3zFd3uMgzcIa9bEcG97UzdVDD+HrxpcoUHEHTB8zGRKImH5DXhz3eI8u8yORLfKPV/pn
PJ/qIUvQ36Gb9DAQEwH4+9qcm+pzSMk9JTbVcSg7JBqVuJTYdMyGy58cVKqhEGxTRW77GTpY8XL6
6WPrPyPnYrP9wTcxz/rrAfZ9DzNURVx4jMqWdsIJlHtDo7YPXEQvRIrCPmIGfCPCgk9YzYDB60yM
lETj4HCF4tGYYMSHaGYYbAriRIC8WUZeDR0cQKYDkVTXWXma6ps5c7I3T/JBgnnF/k5nOBbsylZm
TgL6fyw0oDvMipXEbO6fcNIy9CFSvolOYrxmWocW37f8A1QpPudOEVxd8PPR/bZk8IvLtJ1icXVF
jylHw6dQDBsEBrFwfHfkw+146DI0idMRFxHiKmNNK/EQyi3wBDUWl04eepfdMXGw7GTs4gXIM4hg
2XznTFwmtljU2zR4XH01AzYR90cR7mFKk321vs+Vyv67yuTEvhxa4GEQblpBIpoehfzh33bFKafd
Ldo+T8UwXYw3Uv9X0M+iu27ZU/6MXDPTzpT8H9NbANgGS01ds8vo03SZGmrk8+0Qa7sfg7MlebzM
VUcviaosLIElt8C1Zdynf5Fr3ZfSMXx4MFWLXofCHb9/AM7Y92l1HMpwYtpOwAAeIV/D++CC2lfW
JbgvquRIz6mJiyjEktyqxO2mZ6DEWheJ9AyBAQwsRtZZX6/9C5lQzloczF9mIuhbBcx/jWiseK1B
78YHGfcGHGRvAyGkjGyShICrXFWFXiIXEz6eKwO+WrXfcCjvgCaa8MeiTj6NzaGO583qUp9xtpb8
R1fmfJssEGIifgBO0SjuCac23yJ+E5FTLKW2kHhOHTw9PmAPvWZE1DACuUU0r2GXRp10HPlAAYAe
7Ktg5LCPf29qjnat6QLLkXA7ZgNh7JGMtuhob1u0YTaDtqutCLfAQBN6eYMfkf4GdSobxTZabIiG
scc/XLjpmiVqqDOhNl0Wstp7bNmMpbolrYJeNh4HHTu3LSOBPSICHecFNMcAS/PV1ubbg3P3/ukn
MGqEStF/pjE0h2qGsxH8o+THdfHtJSvkd4AhvOPEeloOEWAQ7CocO3YakxHZlL76rAVSza5enolT
6/jLTj3Ip3AqRNoZD8zDcm6fSfjNShdAn0+JP8+ppTi3FEcGgT14pbj42vKkF5GNPQXOY+pr/rqm
bW4NwhVDZdY/Q+AbA1CXNj6iUsnblJhVmqoDuAHiUgsvdQPyyLD/XnBQPxbj+rX/28FRXRV0c0vm
lUdm+LZyLTkC9EUHiEM7m4Tom383nmfZKn0gMD4xVjBYnki7rrEzT6BRPKROvjyirkMcpOvNM6oa
q7HPDsH0f0SJNBQZOseBKkz7FG1RWQwauars/rrGX/6DwvPqGFUMesVY5U71qIqPVMZXCgY9RwsQ
IjVchafu8uYiYneYtMP2JV2fkmB9MGnIBw/U6lR+bmE5u8n+Eg/fokg7WxdyQVhGtVFwVkrHUrgM
aHHyDhXuhuPnRgN5IPV1hwGE5thNJ14zoYkPeuG/0cOaDz9/BycE2lgD1Lav3AaonzrJZ40XW3uO
RaCyrWm6TscnIAdSLDa/o0msVUeF4f4pWLFcoMHO0JZoaus16f+Wk3RjXKZsox13k4w4OV+/EMou
BsulNFoyBGf3KjpRSfbVComOh4hKixBcMOd4A/vG55MKtrZOBvyORQUbGOwowQKxufsXsgaXticf
pjxnMnB5omHvNhRad0snwT/JXJ8KHp6L7In+eV2QmydRW0KDBjhrhtnqFr1dbZ2EKpwekyvag71A
Ii69waxi4QZuiLPs02hsgPuu02mkvtJl2gPz1OS4JxUJRKYw0Lsx4bB8fOyDmsZyoEthJG8JCpJV
yGYUM6SKkpMN9TSJBYHuoH/MLm4lqF17DNTKvQ3FdevafXFvzoefla+hJFGBCWV+RdogsKhdNGNd
3AVH9iYHKeaGwhWOiIs8gce9gfgTurxetUee+7t7Wj+5m4mCW/50v1IphM8mNKd9wQJFWzobTHIO
zxYse9MZszA8b64Jk9su0EkOFfATsVR/BWFCI55Gn6sdB01kud0wm9VZhHHX1RCp81FY6i49/PXx
j4sHn6qP699cOaXWyJFpEXHLbDO/Q/PC3eLpxXkClsckupL2eqecWPKCSp/izOXD+ihOAOcvc1fF
JQGr4fU35uoeoA8E9CQd6lubIf/zZI6WeqgIE8DJ1s1HqxtJ3aR+R9joWbsZtLbEZz2GVVAEssCr
0Am0PcjwJx7nnXFNE3WPD9O1BSA3wwMD5CTpyxh20ZltCAhLUon12GkruEASKImIPRzGbCgscJ3X
APuK5s6JccKZYhLH9IGTm+ZsXKozFbRp9PD8GvSXggxDyvpNWNlWm8yrspmv858qzFHWQUnIzaJz
DdwfJ+STNISngEV4PKIKPd46M6GiX7z7Lx746LykqH+Y35LF5ZE6O/yF0dqnXkbthgGkYINk4IuT
spnL9I80swLNPBMEoMIWshM7hvHtXTRoUDt7kdg2dXaOKNBV8Uig0p564EWPfw1GYIjj0c4GtuMb
Nh1bKxcWFuYjSd8WUG5NKugLqibdqQ68Bg8K/WZ9gM01Cb56IwXFrg3yJnj1KoNdSFO2OO8xW858
cBs3+//4NlwTCxiEQyXpbX1Q3BQPACs703a8eio5kPw3LrW+m3QmomJRHy1v7Z9naUMYWyeNXiJq
V36smTZ9A4vJWj5VjUAxqv4l+haMO9K78kbKS3KQVUKoktGJpCRVMUYHCkBqE+MsslAlW15VTFgm
gkIE7LCSZtCYwXO6nTNQOtNj8TQhZJSNL2ZSa4WtuOqp+BvapUgS5SqY2Lzw+q5D1nJkFga6jf8f
k4TreIH4x2kwA/NH7k7dFoQO6hPcG7SvZtNQFp8ADNdEURNaMACNAwxr36zO178dy9yFaAuoUbB8
/ydkhSDrRO7d5Zqcs4kII+0HYK6HOgznPBtuW7ihlU3LACwLnF8bcJQnlCfBsl7YDpXim0HUQzr5
OHOaJ3k4Obwug95N8DncX/Xb19DiMVW3S2+amgUjzpi+umlZIMJ7J38gfDQTmoP8++95UY6WJueN
Lnj2c2Gx/JJmBU/XGmS2qitjAR47vYHmb4oie25MI+Ks8++mAnhLRb/OOYJfHg6b9qOsmXZ/3V6c
LXTYIHTCpiv5x4E0hWXvNKTNJtCxAwYZ0WizI4c78ZTHi1zQ5etQkFOFG+uJLDT7oikDcVuV5t/g
RGNUVooA2Rn5vkIA++RkHP2siDffNd2B0mZLn3k4GGd8TjYdADRgQjNQW57WGHHkxKldTdp+UBEz
joWd/X7MOMi7/C9oRo7pyB7mHTxZnkuNtDDefxUrYgJwyhsycRYCDZLPEzAYZFQm0RvVrQrFkHAi
0HYDRojzssjSuJUjkLWr11TEaorYSJsqoNwMXSchv+WKGo5NnqWdhl5yNTIRz9/9yUIOnNdf8isA
3bRuj+/WNPNP1SG9VlurhIm/FjBfwD8bxvqYEfHEbaTuIQp94C+3fw3VDo7nyDUQGvqzLG5g25Us
Ca2lzdyurTj84E/1MKDx4eN0VernoAOGxt56L36nd9cdyy8PEFveREsqXpB7czO06jFWLMwURX6l
eGE/PQ5t2UIeVFfvbdGl7KesBV/k1sR3AuRRxcvy8XX4ebRH5I5rF8nPuarQQCT8Z0bJ5qu4HDsZ
S9aU60GIMSYYc4LQVRqNTDKUhd8hymPnGusYBqDKKsjYmxR6j6fJCvViiuuBLlSdHngnGN9KLHRa
UkNMBIL9aMfTDsKdG2Y7fBslDOA2C3Op04p0fmef63Itu6o67pWyOYonfrMq1LKUaGrb6o755WoV
EewmKpHePKwJQlqOh6C36UGqyZO2SupDEW0esxWWCzqawzF+FXQNP1sOtQS1+RqXY27bfGPMgPfw
vS0POLeAeiNh8GVobmNNJn6A+YZKtGvkiW7F0r4zOQgS12unykik8swtAfoOpJEMpmkrajyAy0Ui
Wm+JIHOR4nOp+t0uA+nlZqgwx9uJ0uHm6u6EeN22PrvNYifixlUCdvRaG3RAm0EFj3QJkUtCHxTy
wORhLdQwXggSFnQQsX2H1ffAG1tNirGn1raIGzToyeY6gA3RXGGV/05LGndk+TE1jNjethRmGzsg
3X+4J5naUC2TbTbUZY/djBBuawldxlHBjDZRbf6C497x0X4mATlO7O63hzyMUi9BT4M9yko5BJMM
9sGLvUHozjeWVAHI1VmM5ZGZTBRkLFE6zMACCVzqofRFrc1fZcN3gpNdBgT7utTzWBZtqmmrWsiP
Cus0sxEEqv2IRJEaKKPq9ooetDUiuOjv7uv91RPb6n5buq6I52wEsJ9DqUSv/LWXaUISNIJdg9h5
sJjTxL4PtSxOvEs0hlG5TIzJdish/T4bLEJlYjmBLCy/464iSfZn6VbKp3f0JI88oPGGtVILwIbD
aK26wwGfaXyxR193TZC+Mt47bdNfImF1JWM/wHx6lJZxkLrBxR56NE6aJks6uwKwUG9maofrf+oN
B9mPE3ko/1xTkF/6c5WC1IQ2FMWouucnP7lO0dAYlBCKMm9nPXdEWbs1/RDmbAIMcfHXJo9MZa3n
Evh4txDauheKfB3gzEHcbTnafHvECC2ZiZIv2AJG9kg0PXzc4ZyD+XKlNghk6uPz5A7TzyAklVzD
M3uHeEu/tOyScKHh4vcq8QWLRwMBOtLw2wWu3GHgQ6MTCw53HltU/NuLlerOSLl+q435pP2zF0tc
1fkK1u2mbT7IqX+6qGXrLBUUM7sCOHDBLL0NEIQymkFwzu4xUFw90hUqBgxBhdS/IAd7llYFFDcW
v3UY7BUZUN9hxrCzuIWXAGv5WQW0kXJ3PtBAD4bJVEqUeOcSZsPKwqECu9iLHuWmUuDWxEt5qk2v
qEbedArdp3T9jjuUmI6nka1/KCk6DKUWVjDNpuC7ozkPQTcd2fd3TUFElbqNxdJ5irOCZMhQv/3O
JyGaFq9bPfemRvuEKEyIRNSOtiOMWRHixLgtUvZ0ZubyIRT+CZ/RN/bcOe31smDXeilOFMTtjeSr
5FuAf459oUGJ8Dg2bUnV4ulpgdfPzyHq1ixcTW3m3JmIyrewMH9wSu1hm6R49p/5ht27+vMOg9Ji
cJUkEvFR8Zgasu3qeDrfmQqz7sDXiQOX1lO5fsbJZdMO2osmTJjZ9ZC3DpxzflRltDRuvxTHxuvx
Iti61fwYStdJw4VirxpnD9KtDq+shjJDdElfMzoVRT3VZpHKOXZ5+sOclO/cmZ8CmcqDqfPLNlfh
v8LOV+blP1qp8VzU7tTTzFLnLTM6cc6AaDh7WIsZydTLGvcODJP0wwcKpvLYS653oDsWhaDDvZNN
9vz8LZ7ra7jZ+gVHNKXHXdpmDESWzjqXrfNnGslo74RtkXZhtvzWUXHy3xKYFv2Wo49TYN3fC4bX
XHFlAueMPzxpia4x/rhPkp2JpX+PtH09KLi2tv5qwLdIJhXlrqPU3tDDv1HtixRkdjHKOKAWQAav
vqlGNDTfI6brz9qTwnLvWHHvxor7rBxabygmimzju7dTqlrU1XKIH0n8tnCeis58mQOPFrch8Qj5
xl8UU/stCtb6ae7xHonrI3XnBKaPxGNAhMPkg3zf5KTc88B22DdVDQa7k/x5sDUpgrVXop03nZLq
ifa08Q2nkScTUTniOjyT2DhwKjCBqL5hxov0zHQsewekIvx64FTTa+kq1KT9qGQjzVKZefqKUKi0
Lu6jc36GfICY23Rt7DCne75FUNQm3ODIiJyeBiypZd1THzCIaZiyqzGtD1KDVYWX3Vhj4DB0tdyz
nGuHni385LKJhFTZJNxQoyjm3ziKyDjFscVQKNXXEB8aq0oMtg6FRihF5/iJaMamvLkvk+zKhspY
72xHh2V28ISeXi9oHSDpi7j1Uhhh5KyWOAZ92uwn9SIIPrdQzzvi9cH451FF0fI4dkbng6zArEJM
0SDpFpa1MT1ndgy8LneZd6FLwl4Fq+HLS5Mt8Rq2sBoB/PMCklnVR93uEPBwztMQ6JviI/+GKqRs
Y68tWE/XbcDtsZgl82QFzJJNMsRj70/xz/RT2aX7A8plaeBv3pkPaWc1stuEhlxiVyZb8QujX3/x
gUqeyZC+HPoj7BkqrM4zz8jI3woqFRqP1njN4Sj9o7zTHvUXZcjaRvirZZ9H7OF/jfjkFbr/8nbY
Ea+KO1yhIn/VwWcJN6sl/MGK3V5OyQYJwIqLYCSg6UY0BCov9Y5O8Smi5fNMMSpqeGCmE9uZM406
FMecjFtLgm2OieN9yY1itrmmFvDaiW8EjweJUQoHopXdIPZzbnwU6fUFyfkgqfi8gzq6SzAM6OFJ
g/eaqqAmT8qH+N/zeNItqJu7y9e2FsfS2ceyuLxXDLVsjTiADFtYP+rm+AYHXdmKseua5DNmNiGd
uoA/DRX6XR1AajnIAXtj0AWeKly/q4ntO6uSZHJBx1bdCrQrVDgWhs+sxuegWlhgZq989wgxXQva
+kqef08Ch3e1EL9hu5i4I1Jnok03KzE4kwzNfWSyN3LmQU/yYQugiCUNQ9asPkwwYTjM/ZKhsKlP
mCFaQfpLy2v4Wz6dlLjuWn67qz4tqoLy8L0YOTvr1h4YyuqQaHpmteCHuTQNACuuo7d41MoGmz+N
4oRz27bgqcDL6XRBH1RGtq6UeLFMFLJr1HOCoz0c9XI3vDrFiKhTkMjm2PBACaHOOUG7qJd1D+lw
SqlBmg2SpIC9bZG+cz4UGdQVWrLC7D1ZaH2ksxyI+xuTDwMBPI2lt8D9CNzOcvk1MjdQCsHmP5ue
dqCaOGcrXXyhYlnaTh3HSjm3gMswy+Fv01XABVdAvcmn1BFnSYe1hTWLbLZSgY6n72CCC5bSVMHX
CBKtw6B3hJ+sdr5uqSRadtTBvTWSurNMvGg/IGOinAKYc2F6rJn9+2NmRQoPx8gwKHLMUeXTrmQd
VPQx2fZ+vC24fdSFaesqBGrNk7Fbt8mRQQRHAOdNje7D8uO5c8B3CTkcdNif/vOvUFz9JpS8lvAm
OuYckmqszzh1j7P8QhR/dywZpxqn2X1z7F+bS8ZMvzh9KdFW5VTIUGK7OCv3Nbok2byZJpNnoqqK
wv1u/JLzgOqiiVFVxmObTM8unqgY2K2QgFyPMc+fNLTZ/6Rrv3Ko7qYIAtuL1UluVqyO53Y1PyFz
wDr9VGQvTu9HwDgYcBhxKgPcvw6/taALECCqcbw1cFgjTeds8/aQesoR+uTe49CQZg95C4f2TGWq
FDLB6HDSBMS76/JJtd919mulrdoBb/bj3++cDsQF5LO5Xs8bESL0wctgYWCwGJ2xjqMLg/y2sBFp
kVcl65JIDa4cB1U/jxgZi8KSktoM1FHUP7DMTpWcL3f5zSpZo9xHvQYo6XttMuTSb+2SXB6pM/Th
86tn8AYbT9CB5QuLUP9IN4rj4nDESWIigJJpR1Z35pOKzsdkJlvnx5QfgSUphCUnehMNdfK09kSQ
CYYLC2I82Nw5Fd1aNs12EkwxH+RgEOMnn5tbtU/FAACqfbWaB1F3SqMQP7FpXHg++7Rj8elPpJgG
+rQ54ayaji0Jw5PPiphKudr11Ng/eScxmVTbIaPxbFtI0u0rccrRj3vUtHjF/OmwvcXjKhTHSWOv
oHBQfSBysKjBlfv6RG3HuGiWuCiKGtT0Yte/HLNuDAwP8JYxiIU1ZQt+knjQXpeOhLVYm7Qz4uUM
554REJYNNdjiH0cWv+lLHPm+KlJDSpcWFvbpDDxbhfFHz3+pV5gz5mP+DMv0u8yR0YM2VgqODfR4
e2zqe6+D8UoyB451HIMqbEG3+vZTro8n/C0bDInjJfLaMX4pREBGTLrdufTIMmTkR4zWHhefljKK
rkPWjJixy7ZfDnQLH9ZYHbg+OxpMl8mJxC4qVNkjmt9HnBDmUSeiOXVuyTIzVcxKJEo20skdikg3
JyXG4+Kdi0/vxR6NuSm2BKAx/gyppmBB7POT1OWS1NT7W0mLukOAhF96Bn85wTpNWAwjb1L/bPEY
rXTZxuNzHf3CbVanL/pY4dp0vY45C2UFM/JJc5xQYvSH95Oam1EHM78+z1Ia8mcNukAFnnoHjoqC
7CG9Tj030yrPv+THTQAERzZhKnqt5akHSI8V9nLYgX464Ie98Ui03pwBet50bRs5pTbMwX2B0bxP
y7+d2vI/w5uaKz1dnyXhOnvMyhp7D+soxulqlxi0hLhzKouBRRVYT4Z9lTR+OLpjzXXT9xRHy43r
ID7S/GTBw6TJyrz2Eg4UCjFA7gwadH3PEnF1/qGcsfdFdnpaXesfKJiYRqIvMONWG+ol4b+wzjGm
kU/VWC9U3fpJF04KSEBD0ElKXkL2TJ9n5+53+I+COgvsgGh1e2Lm/2A0cm7aeuZWC/6eV0uQhmMX
E7DFixBF5PUbRjlbTX+xwvbgA+yD+o+JRnccKmEGUAwxNVSNKTFTNRqR8TNUfEtSZEkvv0SBMU+U
WnZuOYQ4NUSKy/WpljVLMv2pQh8bZGDok7/IVWgy1oPiOqC7iIerDACUJ7xFGnMnhOKZ3W1SmiE3
eiVgn6/j1brp4UXN2wVOtXYkTzpJx2rUtLj8iRAABNozeQjdT7vvarFzG4eev5lqK2rWAq0dTDJD
FdtvwrNfswmIDnqPMo+b8eeKMZ/i/iW4Q047Qn90olW7rwgVBBy/QldbJU0a8fa83Yc+fX4WfIvv
DY7Se8OQSaIOlJkv8a6V7rzuyDryRoNNcVZwho565G44Nsx7sCkyhXXGDhdO4lRF7qYv9KOeekGM
B5yORukLVQBoy/fgpxxqvaMqdeEpTdrXi1loUxj/P98XVz16ltII3gUkkDmJf1NB3jMxbjaAlE9e
fK+ReQzWXuyMA1x9IHBcNWg9l1FjnV9kqFOPhYMaMBt5G1vG2nRXqdMKJyXcYgXXpiTexCjJsr/j
YAdhOmovTx3TsyRawsHlV+NQ3U4LvazswYWRXwtQy2sJVjZ3D1c1raMmud8zgd48kdS0UKoYPAGJ
veuCzCLFoxhgl4LOA9Hw429umJWlNkAjGJLZ9Z6Srs5REWyCyQSW+/2sE8D47XfCkcL6HiRqEzif
8S1ffr5QrAsiDXTo7S3JThKQnqU0SRDvtWBJ04ighRKY+IZdb9oH1KRdnc2kEwdZ4S/ceuNgpkeh
hywZjqf31hZCfS/5gHRhe+xEXCLeiSmPoSU/UMUoxGzg2div3XxAz8jXCI7GRwBHKXVZKNr6iFUx
P8AHZCYTIONpLT7w3SFiplQqwjip4Le7SwXIh4dCTkFtf8AX7P1WF0ew+RQEJF8aenTWrMFoZ+Il
4lnPezLhOv0Y1mczZi01dgto+L+YqjeI+kX+J0BHIx2ylKJ/OH1fgiWVsB/XENvuJQCpHy8t3agp
Y7efGqLfC47xcXPT9JWJM9zXUepjzMCZ9p5WyERIuQ3c5Ok8E46DbiNNT/H5YCTzEefcDoBEsZsc
CnUV9xFC/FRdpyxbFCGnsx0IWFAKd5PjqyCDxivScQuIYCCSm4e0AAxwKWELCAG1LqwfYfnu3X43
qGqrrjuN/Qc0iAxjaMI0355arhCGmLQWmQ/pjhtnIL/9IZpk+qf9EiguwJWx5W9kXA0alAesVzWZ
xbE+xEtjw2FVvTmGScdMpE4riV5RqB1q1nKweaSzEsZW4Kmqg0Rxv6aYrR6L43/xgSqJHNCO8VqK
h7mZ1G4Xht3vobVG8XWcS/VdH8GTc7hmNTawkRJYt/syRjKFuNyVaY0fdR7rDf3ZTDpZk9JgOMmV
e5j9J5J4ntky4M0ZWGc8OSbPSZBfcJNjnRNO9JR6nPTzw0bLmXszm5d5op/72dyOFxMt010PcnXb
YmaTLSzMALyOge7rgnnGpVSAwRS5cY0mMWQ/lFWc5C2AOzer5RqGEdx28IKbJVIRx8IOCLN8R9Yn
q32egkXOp6VGRsOpn/noBtfNcdbSfXpYfV7Cik8UaW+qKs4DDH4GKW/GcwaIZH/q82diKBbB1rTX
Be6Uuq1QNr7KJRM0jT6fQ2iI5Afjit/s+vkY9kXgGOQokNeCTfHEJe0bqNAFQCl01foMZWumfEnM
uJ/4m7nsQEpLHzUFgCsl6jM/1yg3Cy0iUeWpDNVn/0CWvSspCxG/+raQ6CePNeX3buWRdse2WvDx
AFziRxGTXhH2tpv9jyNQk9UsGcQLTdJBz79lEridwOGPY9vCiKK/ig7Io0gYxwjBZpncly/xFbOx
G2hV1MB+/P2pNlRA+GeqM1/CUpy/pApQmNh4Fg6bsrndQp29MYMOOD1mf3risgrpC/CvMDSXEdhk
1bpQM8YpoHXtWL8T+hLJayCSgEA95PN+jUsWuIVOx3/r3zJjMqN9Ntz5OwIrEeKOvaM3h5fipO3J
y0d19KGsYLmWtmwW2NqZwK7t64Ka5WYIOqN5KDy7pPhyj0OAPFVSY8hhRDWNrswdv+P7ur68G9IR
GXQroi+KJo4bzYykp+d8mNe5oZuQHulMNExG1MZD4FJewTSxUs9eny04EZGLtrFcAT6PxmOM8Smb
Oaob5zOjd5plJSxWxOomEIN2aldRJULYBTMg3ezT+nAssx6ALLsC2DP+DdShT4cHj4G5fy1Yf1ZS
Zn8rBUbeW5oiZoif5mBQrLkwiplEW25G3jOF+uABYDiN2Zb9L9JxPRaSMjWPinQwcEaTvzMIaESy
Cz50xWkSjdr6jLFAxK1Z35gettAuhFi/r8vyjq8EDtq5UHDErlSsHap2iPPcaELCmwStqpWMBfF5
KFIgbA5Qw+EttnPUANkxobFeUN7dqQdZI5bLtRiWiCE+MC0qJrv8ZFzcfRLhffXgRbi8nQflX8iL
auJ3Ae59xzWQUteDYZ/tk9p/FJxqRTWJ7TRh1RtUFWIMqSMa8SiPjexOBoUeQsQHVO8f8/ClRonY
Zwqw6WZbAMCgSkhi/jIqiKd2rPhCulWg9KfrWKX/SUrWn0Rr3mloYoOTKRLvuA7Wll9uoIbB91m+
BbR1y1biTWH7ItIaLHwZgP7YdqXrSBUtGOhLOyaSJUMu7qtuCRrmleZOA0CiquVKmITH4BkGENei
dNap1e+W+euceMxtCcHzd+qQbb8snCFPeKv/Y3sYgny6C3u24PvL5+Ikq6z7g3ZqxOxmm1ml8Ty2
aAY7p0FPGppSOJrtt3syswZ216EB4K9GKYLpBY4XidoLdQKd2AIyoE3aVpxj5kghxCHYgFSYGoeH
IIEh5Yymf6mxNcRgRGf7rje06Nj81GD3DN9jp0iZSeUU5dqzvq8ziYUKeb1bZJuVFbbworUKMoZV
oKR6wxlbGz4jHIpXrdTHCW9inJLV3A3lSJ/syBUFKp6ThwYNuQxOua0/yo9ifi/02drR0Hc0c1xV
VmxY7t41kqyqx8pcX4xAeS56p27ym4cWXkwDgTVzQhP5/U0n5NV9TAExEumLoMs9Sg/CZCWgY8iP
xWYeuLm4gKscRWz3eSTswGHgq0w5hrDMkxf9q5s5rOxzT0c/j2II/JEWujywlNXUXzSyh0m7vUvr
xnxPX96l2P80t89i9dz/V4klW4F5rQCiT9JQKUu8dYJeyaKapcRBXmIXTz7yZrc1mk+dGXtfaoI3
EKYwD3u8HxS2Nva+cwSwk8c6KwhtV5FfskghfeySbiV/Ydhaxps8c6XMZ+5OeiPVBubLOOfhE4q+
oop3W7wWTtQZTHQtzITOzAn+E4AOOKdiwyIBweVK6O4BOEHiuhPWx19bf0bHDo9+jDjbM/JIv4It
Ac22RuJhcwN1OxIB29JtzqvAaa2j+v+Wch3haiLUMoGiPWz9Cjwhw1Dnhf0gsDSnZroO1cbWn/B0
SozYbJdKZDvpSeqAqe5OVMpmouyndDl9w545GCPKceTFc3l/a0dF+h7B2LhkRSgrEj2fvyUHTdlr
s80nSC9rElHg+fDJgQRsFwsxaGClXUngOEwnQ9j8gPxqzTuZM1aXO6S+BEF701wsaSZWO0Le+3ue
43zRwZDUiO798Q8e5uZeVcEHwuDlclY6svhrvDBMFWUWS/ZiFm2XRopXeTwztbJshhi26k4Ss7Jl
g4ZhvcDv8HcO810YcYI5tnd6F0WtvOjSCmACXXlgmaAxeKnRqiyzYfuJrspvBilmNmL8Mmu4MRKn
3nCuimWFsCzhaF8zyOi1ZlfvHSae5Jmxpt2r5nmpkEXr5iQqlDKNkJLHzPnhJxBOeOVb+rTaZHpB
vDmfIkVn6Sx+4Wo3RBqKkVQ9E81N8p956UYE6Fft0lqTMCekW6oygzjIYHDOt0CKIQ1FRj6a+8Fc
Asj5HQyzdQvlXjvfzRrCzifIqfe3NSTGVhLCn23dzJ1v1Qith215JyWMLxSL+BJFfVZk5ch4hOow
4mJurmJG/5NvkiuRh03cyRyapTNPYECxqYyqYeGJcC5dIKW0a+aecMEigV8qIAMao9hfYnWwSy6A
8rENHk9gBMwNMo0V5MqB6bzijjX9nptSSNIaWwfYeEB1XDIBDdPFHfV2UAiXmIcTFp0huJOvz731
T1Nlyn3ZzAUMznvG8iZbL5Myb/yRttl9MKv/04Wp/bBWhQfAfiw6u0WeaAVqmQZlU9k7Ek7k0c5m
+y/zW4ZjfnW6pdwMtNaqQXFay2Y1YmsrzmkvXoLMSBJbuAj0VTA08PzqWs5R2aL2rrU+ahs3vHob
6P0w8Y3Wha5AHpR8yvkXLsikwtpfrHfUhaIbFG7fFzpvAdlnWqhywY+ih1AzSLSj8QhdiH9m1t/C
YcY6TmmfzHPP8J6XicKUk8NGP7dvjkXHjYkiUDunvAa5iKkfjhHgUzvxMlBJ2xv+nJcd0dSf0mmo
BZM+w54lWdBjB4szStDKL2DfTbvOCRuyg3eVdzPp1iUyUTkyLwlaKoxHJ9brUHXAj8WnoRLdHVnj
kC9nqe7d3WGDVvwYQm60tJ5P6c8XxByxlmxuO/ZQuBpNO6VptFBFVtvtm/Tx5m3jgCEG2P4OXS2t
L3LVN6gKva0AMv4bHxm15Irj+WJ9SFv1INmogc6XSQIFV++8Dlt7A72AMPXHzONElS1QTkJKvtbw
uwKhoiX6Rl9R0nYMfNMGqmLaMMltClkugmxKplzyAugIdBMJXM1ct+m3FbBAcdu4c/JyMIGBNYlo
FXBpJ34TdBLcCbWJ11qXjkCAZx8LqNgyP0Xnk7Zab88cLwM9TusNUcdst6ubU9bBN624naBoutBF
Uzkt1XSHIV2idPkZluOy+WbwCuO2BwtKPEb0GF3prs90akqjouyh0XokgKFzo3EevbFDuFXwL+xT
cGASr5AkaaTf5+/Wgps7YLT4sOXHN0HH225sSHr4XLVnR2+Sr87yNowOLXeTNNwk5heExkFk52Sr
1u2vEvQcOoJ+gVVdPWzzgBzm2CIEwfNuBBEUvxa6/BwR6z+G3wBOQOm7P4GBWXo/pIF2aPJiI1jO
509Qk3Acp9oNoiVQjR+eUlzLF2EC/wps6jzwiy9ZVYfVVDQYg5AG1kplx7bu89e+1QhUaFq6t9l0
oHlRYupqrwJrMyzlwPqZom5SwJTmpkTXMjFZ5D+Q+s0khRJl4mb6CRAfoC5h3CGb/Oic6VLdiRWJ
hpSGbYEzoQK7ANilIp4dm5oDW/0V5yU5X7/LtqnmSOETFfD9u5C+D7RfpktyCGCGE/Nw0suGBbjS
JdBXN7BMJH6jSRjImNDD4M41jxOqrHFMVyWW9zXDuac5hvhTm6sIpyWUJ8fUzusKSZJ1B2iSHwIO
h2kUXhc710vZqODa/lqaAHYXlWSU8rSfONo8LwOwXfsMODpt09gLcSrbCBLK5dgHEWr4KfXiJTq+
mo17ZGSdyGKGtLEx2b1+WWp7hqa/d8qSR1cenxxifJFl/HLv9021RVGwuJGKa8N+Ii7/x6IcMCxp
Zmylj8xVRZXRsa1/0dWOxqRLqTVQo8vi7LzS85APNePpwWj0F4V4wjBWw3hY40A6a7zliRJKcWQp
4BdDhGVQjx3A7fssvUyAfF0jQcR3cuYgiJkRsz1BWlp+UI/d0Adez7/R6NJxMyrWERLToWyTK/Ut
Vn/dEqy+UpEl4TO58AFA7OQ5t91vVxW7kVPkKMy0O5Bw07O4ydpx0Jejm2Lvo4xM8zjZOedMh2yn
SUc8IiclIWtpnryclPserbmWwEvygJTDO6u/G3a1VE814CZEGKmBG3Rs6BlhkhtLNGZlFxMNlw8O
kpYHt/PagPWCvB7KZbStzgyl8Yv9FYvbbUcI1m/O6DtFS2Ft/LQtsbJ8Wlp+GM9d9+h5mSUfZBKg
3GL7cc+N3BY/jgLGNRy9xZLaR+CwofDJVxhTbWlMweByjliAV5NCx5TKqGPTL3Xp8c8Ik2K55Kyw
B0dwhvEowkth4pni3ctzzOtCX7vT+Fa3ev5UUvlGNPdoyaSLUHTB990xd4lghUBkgQQQC4/pryF/
WYDuUuJV60nrvqU0i+qNttB5eE2ROSw1Jp5vwDenWkvtRuYjL+oSdpSCFoXScyXJYwd5SKYg6c2j
vraH1NpLFV7Jlw/t2XdO22GU5Xiq22MkZoINOEJqbOVpKy8DESAZJSOg56hO0ivgQ/+c7wetzIVy
zlTg+be5WyfQW51gfVWlRGHFaFj4SCpzqbqrFaHlYOO53OzNWOGr20mKODy8KDKfu021NVGVazkQ
ZP8Sd4kfP9cLZHQ1LQ8mjDfhae/9wSCTPdXcpMfOA5ITusIjpBERUQfvl7557ogz4OTz6nydHCVb
2zA78s+YiK5TgTEKIUjpmQccBadW9YnoCMZZCBicrbbgUhCqYvjpb5FeAHRBMO4H5mml/cQZblVK
mMVUYSWgZyrK3Ol8h5kGWe5g7NLZVCw7jvg+lIfegfNH318DXlcIQGlw3Zotjpzc0/ZiEFGtSBSL
WdinRECC2+CgpFPsHS1u4ygUtFISWJrKTH1wNcgYqNURshK8K/BKbQrX8QkEWukeS2HLGcR77uFq
l8SEul1ImbpICnXYqXW+JVJlydLdjkK0ts6GxwK7ehaBjx4hj2T4jVFbJvhNfVkdz6B7PGptUntw
/ecWBAKYaDuF0PWd6rbg/zjeMEIMrBajcgTfyfOI+TSyjvWyEG6ijajJkRTzgbCYQYmFm1egFenU
yPvzP/w43P2QGQ78lxXIdXZb14BRA7Uw0ZPDUgKhye7YJU44u5geRstTyc5V32PzwY1ES4mS9CX0
IuMkmZUNyxWr7DfwqzeXOiLUqTSU5bDZXZv5Tm+vzmNDqlThyZj9hQX1Uste64+ih5Po+jMPXzP/
RgJ/uq3t98YwpUw4whmgOaZlg5tKlbPfnkfpLJ0oyFHrWenVWKnYy96/mJIpji2GAdKO3CcGz7bS
RN6vByx0512qZNZUcmTj/62XrPbrQuzVRNDqx3vVYZZPhjaYL+CBjWh2Gx/dZRxiMj6qpZ+EzNy7
YvadrRj2+PchI44c8go7JEXZCrSgGYwOJH1+GAQcPi6wHrLnT00WfAKddKIxtP00wa1mv4WKTiLz
nvL+vrfJbX/RfPIzAJaKNA+ph9OeHw+KCIYHzKMr1kc0ilv97JI9o1NSCi5Bz+aP1HSUovSFSWCD
jZhecZlVh4ELayhOgFBAUAMHmwhTQQwJfl4IbXLGU+3OYla3SkKnlXD8st1ukefUPhXmsMMW9dB/
XLoKEDd7IHt1yXoy+52IzHbSmWDzqQfRF7Nvpbawk3v+ldfDr1HYYCtvR6pA4jO6t7WpNOxFU2aE
Ptl2rvC5qV2k546OdtU58a6qAv7Czq3xIC4oKi429+5xk41TX4ilHbRz9RESjHZKuoxdxu6Tr0ce
nBRWLx+4TzH3tMFCHTlg6wCSRwHhGQTbtETJt27cPbCUKwzxKtyIHdWqMw3dihW34FFuyLHO42dd
9WL8ib5LoY90lEvVV6QsKgRkSMEfWHYa3mb/IHGfT8oVeXVcdDrJl33UwQlJUk4/tPwWSYKmXnQk
mUh+uUBGVqxirlC3G1laSL3gmjz1CxUa1F3AIJqWggXE6b/PG08XopVvdxuxVGzfxOxngKR3B1qv
QYgBDH2EJ98M1A6EL6rrlDa3blCALp5PqVTyFhuVv0qZAi65TUhH9AF+YNltk9FOxsk1OtjUqtB/
AZoLNXtLqJz4att6alAclBO6HZkGyO5ZDQNh4yWU0YsIBTF5bjqd46mG3OVjMrC4iuV+b9fnzCgf
vFYf61Yb6+ULjFX6JrIBPIyDGzI5Sj9m1At5GBDNGErHLn4lELrRTiMUNY9v51eGqXdL0Ya76Oz7
aOEiQJsxWq9/5/sIFEkRQj4SYigKyIfqNiCFdULOUm430YT7hD/U4OSe/Rmc/dPklNbkXl+w3Fr5
pReJyLJSv5HCY+McngprLQTE3sl3xTRgOw+UZfq+UGwpDy4mEh7HzDog2u2Oeo2bDOgLENsOXg+4
mdgOUNG6iedB9gsPtbViK5NOorXMN+AVN6Xp5VKHPCBeli2zq4jePXL5sgeg/v6IjldnYrF6cZop
a5yX2DWTD11sNmcnfOMAJTBozxf5rmmhXKy6/VKbZ3w0EsxbQKPcLg6CGwpOIrz9Pc2ihtHITjx9
FbMSjtyXdUH1XhsmXsv80pYPF9Tk2ABkBRL+BV64d2xjYamQVnx25eSui7CievBz0k5aZS/chCRw
5u9eqa4EFvcKfRIca+BPdRuRggwcWedfDdrUBa5XuxslvLB15kkVrVS+tToOIDEEAIjs0loLCqmf
nV8wqlg+owv5CLQUT2a5PZbA8WjoIiMsoIng8MyLt+Y4n0au9VaFXIdAu+X6AvVL/v1bvFZgvrGn
qoj/Wx/IddWTnP3vHK410k69agJU0/W4x2yeRQVk/iZOHrqOcbFZUS/gFRDujfAwqYhoM6jvRVYu
bYrnmXqND9DR83Oa2gZZuwGsaNBiHJYPZlmL5N4FHgGPiC8MOzyDfgfJhhsSEDFMAfmqz8FL5AfW
ibG8HRyIaeOeDP9ukOFfAAMFQc39UDPrbklLTolfhctysRx3q6h/Mx4LI4i5HzLA4dSNC+ldRTHG
xICJRuMLmpzCigzSRj+Yh53F4tLdZtpTycXFrxwy+9oNdRF9TtN4uyRE1XMngqK8FLDn/C25o0LM
3fNt+4D/QB7pP34aWQEDZX1YndBaz5zqZYaFMoG06Brt5liDuTfKiJiD95wH+2niOfVn85Kb0rwy
L8rJ4Z0x7EwyBtN3zJZcx9V5U3TLcfbsj+tOdC+wpRgQAm0GRxmof8GNSWVYMF4IH15/bKE9Z78u
LlHl5j1sv5J7YV5a4oOAc6xsOlhZGN5wRvQq2o51Q1qfGHBUSDdkgJC/KO8q9W0CoKeCl1xj1A/P
CPieEWm9W2kyvRQT0U4jtzckt2lwPnRXnzOcCd6WIbXY76Sits9PT4JpQt+Uz6nc2Z8KzFhDo04K
2MQtrP+2SAty5nNBIHL7Z+FxMakxZJqCrpxF8WQ6i39dGRPsTq+Y6BV+bRrMmtzOhtJMhNdzEG9k
Mdyb99hfODd5nUCjHwAy+xSJbgzWGWCAsrGTjua/2Pt2fjXb3bMPLlw0jMLCClN/Dihb5sGShoVw
s3OymypAhwzuwq1oxxsAou5v0xAgNpSqYpiNMqdits9w1WzK7YrJyfm2JL2qDorGONCbAxXesFg+
zEZ7zH3cEeBBWN0aQUdpH/thRHqNd3l0KCXAU78zVEZbXHLvb9UGly2XvrhbgOZjq0F/8kr6hn+G
RR8Si7ByX9B+1Zy8DXU64sDyva4EI3neb+NtytEB3SRVj7x4OVi9mZgbNiRqhQymMfccmsRA8KeN
Nzh1FkhlkIXnXAINa38nkg2khrpKU/1wnZmamivLo/Un6naS+oJfPsjDwgoSN1ej5ZEmEqQcXHZS
y1TJN1YeOIp1EKBgx342v37Bia0ar6Rejq/uidSwO3163S5Uj7orU7wv0hRL/5QIe51jB+mdRFxL
mKiACO0t8IjI8+fdHGnJrWV7UvjMS/VadNSri/lfS5zZuEDc+jP3XVHxgkkIIgg2BUnKwgQAnkgw
/08a205pS2MwucI/5HuWAYry7PRiCWtLBY6pRdZgMjDqRrwRd7/a7T3ZLQYK/+RPz5/ZIUDF494h
v8QKvfOzeDs3JzbooaPRFQk+SjWKviOQVP5+xkuaBkL6lHMQ7Qo0dFi0SERElmdQWdXhIirHWlCI
S/m/zWzNL757zRgx2rU8yiFcnC81EO8J4nlGSKwslQ+SR7PpyKz6w3TOsh46EndtAakyhs6lYwVV
PPxXdbS28vfkqKTfD/36hYQ4kawAybaa6HKZnDKkpUog3auURvVYGzXpoSfAXXjsihx3BIkBfVpl
wH9Btf/prG6sB1M/Dlya5m+f1psLwc/lPm5YFC6QWcEyG627YTY4uvzs7FKpRukatCJ8dWeCnL6A
DXkjDvAxAUWF6e0BD6hWBvL/Hft9u0/kXGMvRokOjbkf/kIXx0C79IQgEqbe7fsDlp6cv74WaTXc
DyZ/UZ+KIPOWC7M2ZLqOvwBboQgjwQuqymBXRRSvJALjioHEfMAV5CIZ9jEfs5Hmju5FAPhA7ZUb
5mfcVMudYcieNkWbY//y09f7XTNEmTrF8Ut5hWT0sFV2vE5CzRKOobtPoG0RDoYHH2OcuItZ7Dwl
0XG3yG8L7sq/vOPuOsBhYNQJ4KF6SiRaX4NDFe98fw45xwCReLxWyRAB7T58eNjaNVNN5jSrJyjQ
sBTPGheIUbPPmjIlwjlFu7/kM5oZ8OIhUJU/V1ZzAZiMwgMyWgPNmoNGgS8V6SEIKKYucX+FarSB
xXRjEZYZS5wUuRZ+sVBrNS4sX26kvsUv002blfQJkV4wy7VGozQYdwreM5qHPGsuoiHRX3eSgzul
xENdDkS4XDLEeSk8rkWMgUblkNBVtPIIpu6tqKUyBaIRHZCF7KYhsgqnjHMOUJMettUhuM3No9/q
CqkZrRg84YRfpb7OA6Y47jitpySleV78ty0OSdOJju5hXXkHpMvwDKvngfRY6VaeL8TjU7+vFhu9
OKtIyajXq3bZICPiASCcjFQJ0MUkekM8czkSX6Iq+0y4HTKzc83SBQQWcZqzkq4I4N6BYNzEzAIR
tPR7jh75IDIu5Ojrct098GifgwtOTnx3eJGPkgPYUxLHT0oU/Fs8zyRvqPo4jogyLzAuzE2V2MBD
dewLBtWYF4Zbsgu2tM2CnrfDdOTTD6iAf9ZxTCj6VfFmVQsthfp153qS2LPKiR0NWzq39AQfENuy
ZCBPF0IEYtvPBCznu4xWjKQM7G6ntiuC1qrizJUooPs3XwwGvlO8R12tA+JyriQxmrHY/T2n6KYe
Jb68ml8SyzW1n5H7TnYn27Kr9i9ahPLdsrNRjm7ClD1IWRNMhGjFOJghQHz5bKMumG8QAtPXzNJy
Ugzrfcn0geqdh4yM3KlAV7efYBcK0XKhpaOikmzuOdX0DaW6WsmUNJGfIEw5AEc6fCD2UjUlEkjc
+PRDiuvAo57xLi8Dxn5bSkbRDS0+u8L6ZlaAm8cG2Fr+6xNm+1wjR+xVmwqpl0wygPhFfWKsc9TM
jayZP8NVRXLhvIj12Yixq/yEQP3csOGvKy5USXbjCAMKE+DVKSAHd15LsFGRGRDE1hBfn/b01zrn
e5GW8q8LhK4tCSETCr4bJ39DcAsnBYzw2tG0j6nAfXnmJkidcbeODgxAkPenXw6ijoHmaAngCdZX
CKLn359Ao46FVRCoHO2iC4fO3TRsPsk/Ui+f7aSoD14Qb77HHVxfxTYMv4fYitpDoDiiev9DMurz
zE4P31kROqykib5VRif+FIMBQXrFSI/6D4PrRMlvCXNvyzn4BUNMFXON6krpAAwEiSaS5OpW6A45
Mhep6fj610pmUzAqYthR9ubdYMrq4DOX5TJQAZk5y1b8/j2Oz8HZvLijmPJ08/3KRYfNfdlJuvpi
lPqZOKkncty39fNx3tfX/B1AeT6O+Yfr6wj0MonrPXfmw1UbVSk5xlMBaziWIA1XDkRkbBx3yBHB
4Hzil/fikcEcuMnpaz7vSMNM7eWfXQibBHKz2uixsWmb1qq9mDllUMx+EZG0lfZ3bjMG45XaJARc
wofACVZqKnbiuow0wRP6rWi8SpfZh2/WKLGPrrCoA6CvlSmbDWScKl8atJSmiAImYfZlBPE8DLb7
jN2w1NLQGAbiqCplfzJBaSlQVE397HDfnFYBJmMpjUPRvnJcsGubwKrBMP+D92x5U/KqguuRirOh
RKgB1aJnmdU9M3kYCvfytFcXhIAa9490xR0vbvWbf3My41MRB087Y138LNkWJ0WTqrqMacsanqEr
vRE65XPi7bGKRZgnx4lG68S2n9doyaIA5ryLeJdzdL86jRgAz9SzUDygIjG79YTivbO8kUny1M4T
eemOMJL7akh8cBLy8QibBEyJWjoFGIdHSSvlg2vrb7WN22QErHfzeav7NjrHeMv1e1l65jkKTIBw
O22ZQgbhTI2usm22+q9342rKZr4lJuNKPffYSniP5S6mjQ/64Qs4J1tlur3umXdd7llb4hBQSPXE
VQ54YdTf+4Nif1qom7WRxnNanBd1cDysBwN7mkMj6Ck1V4TG4VU9Kwe3ydKfVE2GbxXgMjzZ4nkU
gCHNBcqoXrkJnbnp92jFqTvqwm6NjgbYIteKtdFsSp3gCTeXw3c94nd8WEhIKapFweITuNWXlKNJ
xK05AA1ivfj4v8IZ7G9U9VOYCwoMrTpgXuFh3YCQo/sPSRKWmsGRYRlBPpWxg/eoFPKCPUt2jmQw
FUjjAGT+C41KJuEw56Ggokt1lliS8/SNKCR8oebeEKgqlPP/zCKFT3W8mexTrMx1WAoxvi8wbX9l
PS3ZDDuO72gYgMw+TI22OCD0d8O/hWUHtJM11zXbp9F2h2tZDlqw2AGAwABmsbEsiwHUmwAD/Cb/
zKY25BJ+npH7GTnNFtFdQEjDN7SKqesEkaS9gW91Q2JufymUu+sKREterRycLat2PAArFkR5djJn
btfPf4sEC3lrZD9MxdbVaKskR2jkZpP03EX4LfqawgaoKTv+pynUTbtigTXDiy/vpTtOt/HspoNP
8kqGgmXDNAp8FCRbKife+NknPiK3AVm3Y7b2wF7u5Nd87KlxnlupYtODOyANnRGtvTsN1zMuTyjf
bNdUOo1nHfSOJ6/a6EqkOel0NGCNnIzl+pOdGjmlX5Fu5rl58Gi3wc62Q9MJ0DeYdITYujTMftqn
HE9pRizVVpr9oRgAyBaJXOXfKxNl7DKeJThGxpxrXfOQlNQ25HIHe8RCUega7VlBxbsmVWjxV1s1
xBwzFUk2QmKHjyHMc2hx579s36xeEy9RRdat0EgJu8eoszpw605u26xzVpOqNQQ4mHvYVXuTwzwA
rb9TSDwwtlMUOB7oZK9D7lDeVMnzDFB8uxqyJZxxxL6UmZhF2A8ChZAQaRUjB1hEx6JGsuM6PM6a
NVrxWD0eQ683IySZ/A9ojmCt1QGDa5pUkELIuOEMxmXcRBCRK8DwKmd5ZBjudwnpjBWpg77t7yya
ecxSu1KGQtQ9MnZilEymKb9HPOAoqiErDGdj/T5O3hRlYigEa83xqtyIj2P57LBz8j9jER/0Mjye
j8e+4Y9IdjUdcGS1rEAIEeJ59J1tG/32Ww81Vt/9KlrHyutpP0umVe6N4oSw9sqXoZlPfptimpcR
lce2tgd7A1ouOjBjMlXVZLadw3Ea9Z1/fxsVPjy+uB+bWMex6S2uTaM0yQvGrelfjO42WwPvCQOb
bnQsDSBRmFsZ6h1wom5xDf22lYcSxjpBxNRLrgGpzIyeRtTiqEKcMdtTnMtUOKwEKg3OF4kxmW18
FbNOUAb8wCgoKnmWLrvbR+b9ae1/NNxxVyZaghWp3CN+0tzT9Np+b7v32N80FFZvdu0TGIOkFYAn
Li6hFxK29+cpU83av6bxYUoE0jeT9hsP6cO/g7U3EbhKJKgTM7Z5duY+pWtCaqE4xf62bujHy6im
4kIDpxaLWINHztBV9cAXJPF39ezuD7IXfMfZpHha3zWGmPzwwGaG2VqDHJz5imw6yQcYY+4iwZX7
HrUQ2f73jtduLrorLP74lh5EIWa2RbWLe9iCuh0dPArbboPYKGf3aeGn5akZY/Kf1keNdQiP7qwq
2j400zS9SqBGr5mBpppnE6vfiJqW1tKu7woObrPWSmvFeCbSSlWYO2vp4uuJVquCYOQu22f5a4pp
YFDlqXHVqTWJ2EYXE2tOppbczl3QDcy19qaGMG+qftib+Y8fqo9SP+oKCv3wt06zsnCST37rs0OM
kHYFfpa+rQ8dU6WQB1X7kRNzJT2D6mBtoOyg1TNjpCbSd2sJc1TCIOhMKDj4QzqkNqCboRG/cwKT
14wSt7S8g8dmDkG4xa1FRjG1gRLtIcZ9L9mBGeHriyJ0JEIuqKxl0krWDCFygFSb7UsnK6CzNY5K
NEOEQCEXd91sX/B4Q2uvP9BlhCthjZiL3tBWoBWq4VApi43lBP4/ETEEmmhh2m/0Ykmmr5Y8jVNK
c0hsXlP59eFuxY5yGYJkCjokTDT0S3AdNqmpBqj5hO0sTsaN/JYVzPIYOze1kejOrAAA+C47yXdW
0DbVrj8L2BeCol/mh8QjaeM/hnXX3SEB0Vn1Gm3OADaem8JA4nXe1Cqx0UJg8q9kwrgqIvt7xKv4
TcyNlpZ0NffhcV7fH1p7hcOqq0DJTt6jmsa/zz1DzP4Hq3yEkiGG35kWMMG2042MKVWMGFxHbMW9
RSjmgnaD+pxq/sjzZFsnp0rg6298BifV9kjV2Vze0UjjzpgJPj0x+zG/kY4zMkkcKzhb1sJA17/Y
F+IM0joClBbRjvs8uaq89RNRl5hwbMvTVQZJ1fuw0612F+Q5smzYhsiyxfsGcqFriTdN/7Ksdd6A
5hpBMZ2COkeIKds5N+HOKoWguWtlrHjP4illIkj5qQAM2YSPW1FQXHTSiR1nMomtddEv4KfVugwH
3rLqs7HZVS5Og9XLk2A4P14PHKyulj4D4EwdPy9BdQfQPrf0IIjxupUH1an8+aOHPERqEkEp5DTb
f6J7nzrkbojJL0SN1yeqg/zsWiHL7YxbhwZ31OYgM574OshI0ZHwterse/OasT+KxMlLr9sIzDC9
fSp99Y0xqUDmjQoj/87cKDiV0Q/CkA01K8RjhsvBVbvhW+uGu1xHnEF/dXdNanWA6pNOd6qYoJGV
HT/rDAevbLUNHlGuhXetLfWz5Zp1XrP+YsV3jK8F18QZnYH/7XDLba+NXdENmb9xjeVQ+Hc7ICZ9
5mgC5k8YqiTSXJgtUMWc+r9yMnqj05csJV94wL63/EYCMbwLWG/7JyoX74118unK10HbiNYBgQYC
1AkB+u2g2SH45gsz6YzIWg9R5XXTs1akEfs1xYFHchTtsOwyTklvCvDP3qZvoEO/L2IfakDFMMk6
sgOplJnVi2i0gP2NUNN2tPoS2DIs0NPK2FuxeYjGmbG/KrpEepBuCjzQq0egOdlQPI+dQqNMKQWO
hCmTMBW+3o7WKQoA6aGDUk2tJSjqJN1bkxsfoHBjgeAazZe8yU9pnKre41s5FA7efpiFnAOIz7fr
xqTC5cWFXVxOvHC12CWDZk3GrDvSKvx4UBXLWMs40gTOvyBR+39rT8/Q+6TyGV7aqm5TluBP59rv
C+wtKWB8CaUMKa4MpNLe1XQO6yUHt0u7eORmtsAy4MhFUbTw8G/g3hK0c0Co3vp1Zm11C5klQpiI
pAGOHJZ4bDJc2yjVyMLoi093txUzLo2K/MiPc8aRpyaEvXADSrucW75oXFsDlhNTx+S2/bTVm/0I
eQ0I8XFyT4EXWcJh99Ac1CeXRBvmOr3D+t2p/gxKQvRBuEy4TuZWnNZXtiz5cirIxWZQ0TgZOAmE
ALKAqbx1gKWqxdx7tmDs6J9w7cYyEcl5ZJto4lfHpw9e17zjHfcn16rXFWIkv+yOhMG0Ky7Gcq4Z
oiHHUHVBzT/eva0Gpk6s3Mekk4jF/fj7V69r8b/iU2GLChZ4JHCCtfjQytX7dZOQUtiZiPgOWhQN
/RXvOoEkXsru9eNKXhg31utZkJWjIuhLRtNvX2IPdcN6IVXDdGrCvpMM235ALTNIq1ZBuqtZ3bj9
OVzCU6Sah3MlLP1KCejJCQjMEY9JkfaGqOvFNtCzbzvo4auRS5l7Lx2Jbikq78ttlhGdZ3ZRFVG5
xRnvHacXwVePwR4vgDhzwlqrN8YZZM6V1NnPi1fItkcOYTp88eUnh9IuP7UAa7wbY7eF1laezIPY
iaa76q2AZwvPWyaqTieYTTouz6MZHwjw2KH5Mwn7IHkNgnIPkKvJhdVVuFMJaJ/VdyRkP2HLOkxK
RA405Uwst04eqJsBnV1yPzC/JYwx2qK2oHOWmsciRu/QchfmYhZZU4hd2maS+XbGupDBFtmcTuBH
bMIuryq0aRkdN9j0KnDnbPptaEFyDa3Vx17m3uZRO9bpC7895+TvNSe6P/pW89IwZHja8sONz9Gw
AH+kS9tQDOiHLvQh7oTHnMw2167nFxKUI0VnlJY8aV3OicRJ/3BD7ClbsAScZKvSipByWlMNiqOz
R5Dhi9mEq+48jGdFe+Zv/6J8E9C5FHVeHp1szlqq9V98gow2IYpQX6cGJvzozFpErP6BEsyTME9m
9MuplS60yqA5Ayb/CwYHgLC9GOe0myh2pJJKhynagr78oy8ylqw9ZpYHAp4MZSTSbpqpHo1McSJI
1nIEoAn05gCVkom18s34xDukrFJiIPQ6md7fgs2TVbBXJAQJJSNHiPNPEuticT3/buD4CEZqCiOt
GaOt4yQt8E0/w7nZoLY5WwBGalHrlkswBf8AF3l/fjuUozNQ9aHJI/g1BtwEB3rnNefbKjBvmVDh
PFtOu4xwwWDCcJdPfZ27fk2LNO2ZHC8f9OAaDUmHGfMi3p+5cX093Oji5I1Keec0LM8hQh40pCxU
mtgIKrpL3bNgeMBV0W8/7aA6UfocGQsZrbmIgwyKPf+USiiRvz21OWUsDjbGx0ls9Wlrwm5zA+Tz
AzEBk76k4/ADe2LlXwB9NbQHAiYtqd8/vng66c3NoZn6C9BHLn995qhuic70GlOBnXCrCg2SLTcq
wgljNzX8z7PpAFIO2sn0uspJDl4Eh+lzzQ+PC/hPD8cR2M25aJYiclrI/4dBMCXSc5+B0R/KuuPf
hitZnyNJYZUO+aY3VJehHwl/0m2Rgb+LoQ1WcnN2Syokfna6vKC+gRuqC6dn4b+cD5KKsndQVF3j
KPrAtnqCKMPQ6mDxktnIY1vWw/5fyWcJMrcyMynUrKwv1ZenRTExaOIGHIOJJjNnClQYWSH1ja1g
WLdkaEJMMOhjmHtYPiUN7E6UY1C6Ooj4G6WNqMp1y2JNN/TfWq7tRKCclf6a37OxuMLhXsjQ9Jh4
yw63rblPsUUmm5nI5AqEqiXLH58oTPWw6K/OLx0l6j+OhGUORvrV6ofTydGQ+1ZSUjafMK5ghsDi
/a/VctwY+QEaHoFYeUXFD4ZgS0oNkc2w7z6NZcgodPxfQvBlbA2MeBj60OcMu2dIRBNcwfA7gUiG
QJ31oGkWy1pZxhDtsQw1scdmctkipzEcu5y2e4rsm+BL1TJjukJE1wy65O++783y7wi4NdO5F9kF
KJJlagy9OWMb4Jzmt+qwSWyWG2LSPAwkFuv6FjdajhWUu3UoKxHM6+ghoMeZiXimDXdoAC8zHQ5g
qegS5VngjM56sIc4/l25uB828EqT49FUgwt38wXy97iNfZM1UIHOoaKyD7gyR9MJsXZbKZX9YDk7
A2zZ6O47dCoD3iCOI8XwO5WXukyhxO0U84xRPYqgy2KwWgE9RKQycnqQMPD/zFAV5zxO5i+lenAQ
v4KV23+GmhXtCce7nNCNrr7nv7beQuE5MYYHdHV1Ljj7xBZwf75AS9DhhDCXIQsBwLvns+Pl4tVl
9B2fX3/C5lw4R1Uex/RRMEiuy1+ALYTD6dxqzjEIFGfcisrU9Pq6ogpcZOLj1auZk205mDSuX4AH
jqGLVpyJBef0cRyt6UOV5G8Y0+XdfkX23XX1FUpah1/OC7jMnI8XsXn6DL4s8x7Zx2dny+67VqQz
O2BDDe2VkzYYSqDqJvO1/cCmjfsXc373+ngAPC8KPMlawci69f88iZ+ZmiismmC1j7fTzgsqLmE3
vlni+jG/AW3nGLGVIHo+/Yutnk32YGd2NsYKanXTwAMePTyF89g5SiRmza33pgdimIHDuKb1KTDn
eKAnu7SZFkeLyhS3l8zSQ40JMaH9i3Y95eyhilJOIts9wmosECVONtO94i3es1UsgRdfo4a+mh6I
2Wnas4cLj+j08VjqAM2QhoBHWhedukV253OmwRn4KdUbab1mvtbB5pLdMGlHoOKYoN3CI89IFuBD
PKUDNLN3JTQRSe49yGCbXgZ+31VPXfEaJf7VKyE9+b+30lFixLf69FtkIK2HoO1KE8OKpYYOaJWf
4FTE/BUkWDq0JuTz6+JbRflBISWqvjL4bjbWAAsTe+RBuxfGw0er4NxDDCaDgpDkIeTiTiSVMDP6
kZeuRLcWSWAY96zPzeUanfaJGtbDQ5VDq+felKcWjvJ5w6Hqqb/qfCLe8ByVyq4ftFmKP/zWYZpJ
zYSrs7tZsHjRVRvRlDZVH0yH/oSYXMqTvGsajRLkYYD3DJ7dSpRGe6Iu9H0mkgxQzyOUnpeD/XoT
evA/zzJ0pWSU5KaFNiGG04zZm/8idZ8wltd4+3U2cSzTE76PPMj8a0QgoWK/11X0xOiDZxClwoSM
hQ1QJblY0ziKX+tRelNpEUyw5vOBMyHGaj/E3U9NLwDNe5nox5br6rm+5toZyqPMBZ3mLUCeGeoy
V/68T/GtLZGKnCS5o5RUfu87KrlFQN6fZSYMECgIYQohkhiva8RJ70NOiPxcEu1mR+2nBhHrxDFR
C2DEQ80sLExzCTSq99sxjFY4c0ig1cxCk9PM/b1TRwXrY5EkvP0oOcWAWhZ0/I3JBwcc7ft4cKOY
USVK36dvwhT2PN4ydqdafmxq/e2bhXH3KfMbunWC3ZthXcpdwHr/SWpHK/d/49aUVj2SJeS2ncQz
QBH3/Te63m5DpAqLN/mWPEXwc4T05X6vjsG2iQPzbN50iDqmmXoc8oethkjiKRukrwMgFi7ILd9/
nCb6F2eCUTObQNWZ9rAa/mM5knOQLGzMU4n2nw+ucaggl3qPWV3J3gNet7wRsu1dxdB73Q+luCbQ
6eqQprBDjxGp+uKxhiGQlhK3F7rGIxvAWMUjWeKya0PhfLb24YbqN45ru18ahw4VN/dKdUplOhoE
qxBw34DGEdp2oVia/0AONDtvC5x8HTTYeqNOV/JKHyVp6BdedlgynvM8WKc3qWMNlVH65BdBKNuM
BgRBLuVw/d+2ocxCVWwEbeiadlStmnX0CyjRMIoF8H3y45vvuZEqWy0eOP+2tGEnBr0n30GOgFvX
YVAJ7RHdvDbes9dEkfjsQ0X5QiA9QSDxCmtDrFh/JfEksx3nJ0irrbIWqO91vOFkXbkYEkk8E2Je
9skF/a0aT6XrGNoxUjpWRQGx+tPSwjCkH+ZB0HIETkcocApOw+kPeoiC2+Ovacf7o8RoNjDcQZET
GjheoDdactkZG6cBu6peeFIqLqq87lBnPqH/yP1pCHTL62WX5igU2We8H4/Vz+TzBguj4kxBAY8p
bvvlY5boyg3HSHKz0XoTuqa1X2Qx98FB+yDRLhXcDDBG+JZablkNeXs4sfcaGiQlkpKLmHzvgZbu
5atNVhkdE2ANm+kGEmOW8RvMHpOaAqyBwqhQWdfSZKZBW2Hr76BmXUJXJGpaXAYOq3ok7pqX1dVK
W1zkD1V+aYJPjgW4PW5n06DJjWAP+5zfJeDy7A5QTTXm9ljAfaVYZuHVn5ttL63KKUd6wKpJ2hyZ
yZNYy2yHJnwhp69q86QNpxbJJmS3Nc+EyWfAYW6TQvzCovZohvvOEkGap2hTMW4rSGQGOq8G38ak
S92MPKAm7EcsIOAmmlc16MWqA/d6PBbhzpF//BW61hxpMDOuZUUazJemPdS+FpaqTEAexcPo0FNi
YWIs28fjRxaRbHtRz/Og/DfbzpvZy1q2edAHiJoAyTPh4MJzuq+W+t9VDJ8YWnEVkhPpnMD+ukX+
HQhUMof8+aSi3kb/FSWbBDt+3EW+/qT3M7XtQ6SiNNQCLlcETI0gvdBLkxVXUctkaJg1bTkW0jw7
ppf88WCwoOZ9sOqkg/ug3/VOf4wQmLfe+Ub5SOzNT5smpCJ53qgIqPyx5xuxvnRdsTFqgf8raZw0
lFYhDcKNIoKJBY0kv/peorEg7gjcJ0Y9vprpkPLu5KpqZzAJDCx4VDYMo1Gzoxv8jgRNp9GnNBlu
YfBvDxO4/PdKdWPfcln64rMHegZyhX/Ez/B+6D88sJh2DFj/Bdzb/ZFAjq6IljGJ6t5Pw3Umm7dn
frZyTuPS6nvvsceEgPkQKUQ5/q3LPjyVf6HA829NqwWeDkf9Ih7ztlEsACKSf10sKbHGmCt6D8Ut
An1TlsGQf/1I+PCA/mpUaXsSg44Ght9TA36giky+fZ0RfjRbmO4oKx7WKczJmlvxrVL2o0Rl3B33
XTltn8Yqx+WCiU+ZZ6BCApXr8sGqqDQWUN8kQ1pM4zxFJFL/+QqgXozoJsTUCV+EdTyZ71TBBnhU
GHa15O0xyKEE2ee5oPKO3DV1tmrN+dEDz3/PxBU98/6CnjMiG/n81nE0a8+gdgp9Poxrdzw+m7uK
Dwcx8LrJOa5UhRpcIrShvq/27gQS86ZEKXWclDTEh+IWvYPYPQlzrG1GENUpWWsDkl1B4Ks+SvKA
EC8ZBNstas9vbZ6vmmqm1TaKwkSVT3zYgPXiINRJ1n+vppCS1uXo2mCP8HgLthT0TEUlC+ewBaCq
+WcfNHUVvlBdivtJ6KLG7ute13CA51HYqIM5lAgKZO1F2dFuY0tuVpf5LllPaVyLAlePydBeSrAB
P6IVLx1DFYrfkZyixwR8RVu3TZRlP3UrvSxJ692quCDU//b9pvT0P5R+cFD3QMWx+u0Yv+CCHh/z
zxifEwl8/jOOKHP7+rdqgkXXddOm1f7kxjcxLW8Uq0M/myls/XPZvEjs0gwAwOPcHP+QvbTEpAt4
lvdDDnmDrlDxtuZ+mffrDA2Muw2X0v7xp8WnzrK+3ML3S6kH8FkFFaQ40evUhDdEHfTErGeptDrZ
GMN8OjgT8Ly5TXhZKmR7PEx/tZC0gEs+ev7h8PCTH07uTH9a/DS+ehDKkHhZUG+2nQOxvMJ2E65K
xzdLSLlHR3mGFRksAC87/V+GmmjWSUjOlf5mUNO7PEnakL+7bWu0ielAT6V+nNMX86oojyVLnIEi
9qgGu75Z7rRmKtMQTMg1fISXq4cfVhHizhnNZ/ruK686PWM4zHnPvPtrLzpAEowcdpj3XaQj2sLP
eM32e/ECrtQX4vRzHPiY74zLIMed/zAqsovmRaPRp6G9vEYnKzZUMSWuA/q4TBXDIoNKCzl30rFC
pWrLJYRGLhNIEI8yfT5Pu9pFq/0HPhFKl05ueR+YVedJsIwgckF52wRftSmOxXv3jTgONsV5l/qx
u5644jnoXHi5e6odXLI+osXokaC/pBlpsNEaPxQFW/BpgzT+dSj1Qen941kyjMwptOCU1MJSa68O
p07O9FxWx6FHJEh3eICtpy3oghVQaoV2VMEKHjDd3C9cVnRLCNerqLPpdX5mJAAenn2vsoXPqAHx
C5oso89wYyuYPhaCBPJWQN0YR5V9LKbzJBp29aXbk5cQlFD22/J1b7xMlno8y+60+EeHB1b0CXyn
SRd4nsRl3lbO9JgsE1uTfhvSJSUqCZGnoOJrCE5PGJck5ArX004G+sqRpIwK8w+lDH20eXV3knPg
ei+LBbyDAPl6/j+hjjtvpCfzumqP7DWynG8sqdNQbHTHLj2rUZ7Hvd2Sxn86fJEb9Q3H1vkvJTKu
t8Pk1wdy8M5ljFHIh+vaw/FH/+qV02NrwIqMXQUAegLsGJjU1tNhqN0Eil4l3mTr27D/EYUf5xln
/r9Sp9NoQ9UWX6Qk7Pi8pb24Sec6I02mMCKmr19UMmuHY9GamE+bv5Jpnz6HTUo5yziDHBpnSTen
OGpVgSTe0xH3vKDN0GW0Vm6Yc1V7ZjT00uOf81JYMGlQSxACKKpTs7mBCGnBqdAIDbvb1FhdlBVp
RCQ2D7j8XsemGXpMb946mmnu7DrrmSuWUNTho0PS6UtvLkFwHvtBJf06wt9VW4VWGCp1D6N0SZDG
T4OilDzRRDwxCUaXfFWSFImnRklJ/uqSm7N4tu9vbvSxujfEdSyJeYQAwcNEIGrP5asMiG5kknMA
m4feOF0Gp9i+/u0nb+gHX3KKnJkEBQIaYOUUv6e22HjqGPvGOIHAiMhDg5VgCih59ng2BwdjjR1y
m6HHz+IIwtHsegKi9cg4o2omc/DO54ht6HHR3k8pHXa4Q4/WXJKRCDUTrqSIGm76OlgteDNDKNxw
tUsqVI2NKFagHmNprIS6q4FNhNGIc+K7uBjeuELR/Sn4Dx98vVCJd7rnq2v9N05NMmayIMebfA5b
+aop95Jr5KtNNyEAGgYLuE1gc1wq34KeyPgfM30vEPfGi98K6czy2DXjco0d5Lz4gDGIuSSldght
MSekffg5Hhxzuc/GIMt6HbAaHtY+DwmlNkQ3WfyNUM/MEWNZK+ff3UMAwbMvLDjR8Q+Ekob+zgkA
0GU7uGPRMjTtXKhS2FajwLDUh6FdFwJim0T1bdDuaxMVTqXByyaW+7so6vRkUncGxT2mlurNgj4V
xaNI3DPdN60tQiEsx6CnUUluHDfIinwrM+WRuXQvwzbHXlgBR0kGBBQTMfIH1Nr4g99LFKH7dAh+
tGpmE2B2GhaTxFctoDBpniEda/2kW0u1Pi5nfJ4WsANcQvpzdksp9VrxYsDg8a0sduN6dR1ZrONA
SO/aIVPR2QpESrl895dXUTE+C/3gOG2QVsFgFUaNBMu3Pv6GuqVW6h8QGoJDGkyaNtcYof+I2mhG
n4Bc8zvLnsScCaLDwAcmoMLgay4uB+WDyJeeqssACnmkk41sW7iCb5/CWE244MWJmTMBqPu8Gm5W
pCqn20mZSCElh2IKLtLicMrlU/x/WFk67U4v7FY1LKrGAQPyFQ4NQSem+ODFZL6t5s6pTKIvERTO
cY3DCXQi30CH0k5Jj4O7et8yAvktY4FMkMlFYTnlTsUThf/XAMDYIdK5iiRuZZ3Mk5rfL5mEuFrU
Ys6ZsxhE0QLf0KtTeehqATqZoitFy+2/Nz8PtpxXnKvUSPLQD/N8hbEM3B2792M+4N8617Hn3EU6
smUeDFeAYy8YUyhiegYYXvMycLwpgIqhDVDRfBPBPEoo2mgcaYgMzd/rKv0/wofnJdg6td9MTTUS
1CTJ5KwM7fj7Xs99D/dEAt/OXdtDFEqlCmeaJ6OwvD5j9dEWJZan04Cm320eKcGvW2SGfM8PaR0X
1/sDae/2F4aVEc7TSeG/AlOvU+6SYTIVrrIts6O+MIVF8Uo8WTWPbOPNBryH51lPJnGMohAlZ4c8
YBMer8VmfCt1LzBqV0ImVLgDs9x/XH7ckm9jZj88yO+g1/oh7s45DhH/1PM7aYxYjmK/F7Dw2Bkr
qVGM1f9Ss0UyxkRGpDH84fFQFzoa15e+XPSkO3MhpsX0tQ9Ij6+NKO1RRt/9Belx0dJf8ltqbO76
AQwy0xB70U8P+cqINTwawUFkkhEpG5BbMU55B+g9bJgxT3MgEOv1Kymfz2y5/sMbIvPxdjSIjFtI
eyg1ukC0d/zT/2lqk2cAz+XXFxo9gaZJPs+RLxVVqProzoMZUT0bImUm7cA9sStKADpL1KyMEZ50
H175uM/1SIS5GBOys4FvqN2hytUhB2QrVmoJKGz4XN5N11Ff4+8l0XyoM/+US2XwQZHCFQaLyerQ
L6A90pMEWuNrn6uAEREazgpVrrw/2f4pOfFFF+swMbEelgz0VQYIEvffwANk45ImUK95IFEc458z
9W1NLNy3lND+QFwcTGFLBjNv/OmGbLw1QRo59JhR2InScHP38yqIDH91TCQmaPFSUA7Tzxrh5OpN
JJnk2VPV00FYBfN4wfF1VevtC4Shrc3Z41SO4BsysA7vEMNx4mNrOjzUgO1x85roFS77sRbLFKli
YmXB639CYAa4Se5dBEpb4klGnpEquOdMskG68q58FuyYQyJOXegSNhgzauRzWhhTD9FUZtew0Q2z
gaeSzHvGY0X1fiIiJyfc769dF/3rg+onecJFuhqX9Ua4QZloVNYN8XRYKF4TAnxTiZu5LlUBk6Xz
nvv4etW6ha+3P2PgMc/WiNtgZOri30cweN4gxGbIh6isiEP6A2hPoOKH+tP3n3RRIyPYkt/KrE9a
Szka6DqFqdYrbFgjmYMpvkWAdxYxLufiIrCRHPFeKxFnlKtBNwVY348iQkX8XRyroQhBIGnauekT
m3cwtovZZNG1gI1MGzCLHqN4aJuRdviRBPhsRrp7lIToi+c25ot81GHIfiKSfCrvVQtN/tGQLuQc
XertRYAfkQoATV3q6scFZmGw/cn3YolNWYMuJmIp6uphIeSzEr+db/LnJa0/lDxMDb/DzqMq/eMg
aKzLIEKZ14xKQmq+wIKi4AZ6C4kR4FnvC/+BHeRa9kVPVGRlMBWmm/8QyHcbTPDpAqNX0gZHX9d3
lH4IX/l18vqcG5UDbqGq1gHuDKeveh4JOuQugMGtqSxsjoolBJ/iyO3rSG5It3lqJ+Do8YGI+ndk
PtdGRm+6gU5Uk9rYjuSFOOv1mIXkD1Kyk62F8Qq3SRNMH6fW7m+GrOhCKrNTtXz83QiuCGlkjrZw
epAex476wI936fVOayjp9PwIcPbwJKfTB/8knDA2OLgoWjwQyi3tqr/jjQFOCXkrqu5usoL6jpIu
/DXJYt1FW84uWwAFrFwPyqVbhzEePDJwsW+yg3Svzh8MZ1g+8A6YowSQIrX1gnWWMxLhPK/DF4Y4
G7wHgQx0zSbpibGAdomp3Yv4btc7gCdFtdTMUugD73p1n275MvTf3CfDNkcFwJQUHKDxNkypsgFh
5mGnINpsByqGXUELNcOSvoFvcfSTz9TnZpr10/jKJMSBhk5Eh07+qt488Hwzm/yZYYCxTOWmUcrF
ywOJJLwSI6OG+spqHsb9GZVDz/fWdPsaMSmSZyV04s3gqlyZ8Fae12ZsEFqG8i3Bil44xWKcBc//
mk44ZzwtmVROgJI9VngTdBVgeTL3g3gBFRVB+CeCO5SQ1eQWXXHA9c4uDZW6VVkRWN/xhrOr3DKO
TGkM4zykwC4WdXUc+0PQ7v6bWj/dHvoqV1kSpUFGjywc273AhCUhvO1cFl7SXm1cqCm9cn5Ax75J
P9cnsWZi1lLV7tp9fVBPQmZM/g/O5LRlrSVQxEH0fLQtRtrvUo2ANyL2m9uoEaeQWh3HFZTf4RQb
hrTjbZT3aG7tdKeQvXkMm4BZptnQH0TlIylu/Qfikq/yVZb20ka4JXgz86gCDUIifo9uKoH1+ZRR
jzwLS8BUUbSWymqvftFAUokDFLjlgvh1dIUoRObiFCbF8kR1jeiHBA2G3biR853wL5ZTNAbzpu1P
fc1Oeul2bbS7V+nMAkdg1Z0g01awZ+9EX6v6hTwgaB3RGbhLPOKequxQZkMI5cYY9YBi/7RCP9XB
vHVlaquYOA0pAChxgg8bywEN4Nin8+FoXEB4VD+ghO7hgvLCLGXhMFfdBpDSyR5rdNYaGpMx+sjf
ReEL7AQok3+8AniR7LFrDzJ63+7GMWEszScw63HRAKkhmpCtkuNfYmrDCFpZa17WypHVLkYGcG6c
kyPn8l6JSQYYwH+4LLkrNlWVIBqX22oU0sfAhdAwpXOIs1S82hS5E0oOy47GNvK4I7r72ppmw8Bs
ahmRa9GczM+WZ5POybDUP7QzwUpLIo6uRJV4gkNohne0BxQ9fkl3fzV/vdrB8S6vB6fz/jm8NA+e
Kuc+we2nUWTkobBXPHNYPVtZOQdoz2rR0xfoQyvXxeUbYCcztQB0Pf6+okNnAl6KBfgIbLJ/5Dq1
uLQ4DCkw9IQ0ifYD7/7VBVSLQEWM7CDg3sEtU0nzR6632AdKOoMyTOURypdNMc9J9+5tVB1QHyEz
JDH8JR1qO/Awb0mkw/DD2RjZqCv72xmqTNNEwLPU0Tgyqngjk185NiVLyQ8bhWbhEgVKb+TvRj6Z
ll7pcqd81nOOgiQhncvQZr5kJzsPQKr3UEzKnUJYF5K8tAcm2daUn1oIdSQGLd5S36nAcKSYhkcK
2Id/4k1nWLqn5BntlLSccQyuVwLT5F4iBYrUs7n8g3mDyFK0HP9qAnU43ar9eW/ahcHslXtQ6R9z
z30aAtTWR+JJ5plHUZAu/CK25nD/ImUSRkM88i8oDKygy+xzWe5wnlLzr34aWo7c+UOhd7JLaXmL
UbHQHW0WLn26i6gGaaHXFPTfcJayEJz8St0zkXAatEeb8thsoxA+yH6/f0eS3UKuZ2GZPd+7dIrs
PottwNggnoSuKodpy2BI2JLHZuipAgQTnC9WQH2ebxpqS9NPj2PHEF7TntU85yGNGw1ytDczOJrg
v5lYPVGQO0tR0x+aK0HYn8+eRwauE+I3b718HXR3WYG4Z77/EQNp2f4TnlS1udvpu/8a+1FL/j5z
q0M9o++SSdUS9GB/aFG6yVRO2/Ac3OQmlDH7OHqgNYzpKkdLmo11kh6G49ZxqGD/JdeGczlKEdzX
EMJM2knw1S23bZxzCy2lrBsp84MtI0fYlAyB+cbT2EGO8bHBjyzsPmzrgrr+Av3Z1WnW2UDLQgsY
FwQsBo4PlEIEO3ZNQ2ky+x45cMihGLV3GrIZ30Vyz0yRHtB4064TwTBIN7+hQG2Zw7PRBWlknJeh
/vCLS3lxocf++DEqJN5M0efmeN3ayRyYb0gTMhy2ByrCMo1bRbzaJYVHTIevmL43SEAk+EndBhia
shwHPQwMAHRI8W19tn36IsnW+G5LtJcK0VhrxWoMQimpKbyNc9RZa0vRQIun5PcCBEZicOwfcRrB
SLgg0p5zI2Ty6NA3fmH97f2aJHG2vuyi9JDizl9IbBNVgw4yWFCVouMht4QG9lnN0OJ3pSegBDsG
vG0dD0jZ2qQf5kwnaXIHH+jc0HaOk81wsSZvYKGwwlsTWp8gXwo5bhEwF531u429yIe3eS+o8JUG
aGBPZdqj6MI+uDCgwxCFr1oqod9N4m2IEO5QIBtQ6rQxDyIm8NrazEHPRHPKWNCbycWc50FAMyu1
JsJrO2jBej6fapBhVTbGKRrHmPYNVHb3umi5oTIf7q6sqQ0KSBA9dYIcrSpiW12HbtISi88ZOb51
cuPXwiHIZB+ciAE9OZFH9YhRl5uqyRMxoWpvh0dXFkGUQf9ZB4QsVZi+J4QiSmgVzUCiFKftaT5A
SRf0zGX9SZMnGQVxcxEbgmsTAn2oV5kzkMDQ9LTS3RBRqmLXpGNtoAmkhELmVc4YzywONJglzp8f
ZWcevpZR1Tde4q2jx9MWWEPo6Jb4bVxN9eG0j4hH6OKnyt90H0PkpEBLnBEixMLgCGtKVGCMp+CM
7Y/uf1upP7nhMV/emMe89blmK7k4ADwMBUROla4wtCi5oKnFOd/yLAaEuI+q1DCegeryHsqsaKe1
QKGr/sXQ1UvUk6JJIpkvEUhN6B8G+zcQNa8RyAKl66sT0tqqrGuDT639cZX3oiooia3fUhg8+1z7
ojFPTErUbHaJn09+3nA1C2sKWGheNYBVebzF1XhgVtg7eQcra3jeHw1NHaPmqsyKhNdO235AD+lv
tNbPxyAkzC0zezf5U03iNkdJUkycw3ZIKpfxr+T2arxx0GKPHMHI3uUZOy2YPCGhZZpJ1ruPfDCV
FoIfu9NEJcfLV4JhFUuEPuAFuvPLg5qQ6BvfbJzJ6RMAusqOw3IeH6zoXj10Ri/FHNPVTK4FK9PY
wrehWcJ8PBcux0q69YH/0llZQdQMrO5Ty5E3oR6OtpPBAtJXOiLOfeWYWOjWe0FOIptti9cJSPAU
zToBOw/e68bnIkd2pEyZwWJl0DeU6CLAca3SY55r7PYpWgAFBH6cssX0K/rbOCYV3i4w8qU70XOp
vB9hfGqvX2SNWQ47m4yclk3nHXjhNeqS3Y+xdL0W5q4XbCmRjTyppDsl46DqoajJlpKoq7hlAl1I
4K/CFXuxyfY852nYc0NzTgIj9o0rp+0MVdKyBlFq6eb5ucIwDpdzrTEpQC8dWkgXFOD2EKvFzJN5
xC6zUjIi4QCzzVpoJkWg1FzJC2X5lZg2bjbS7ev/nKdU5/njhNp42mvE6m5Vk0D9VNTRmHF/ZG/X
yQM5+Y2SoWtmRjXYUFe2eBxB1AokfYXcSiOjgTBmCvyl9xikKPdLXeGMpYtg6s3QWxGjZYui2Ia/
Znp+pwWDj0ATVlvMKIFrV0YLV3avNTnRUjob+AlrTuhK++ti65o2mju05t73mKW+gZKVUxMmZ+h9
MlOeeW5y1eyMw8R96/e0N7FtKj0pLbC2ttpj6DEVBVQQV/nRvzLPZq6gpS9jATm834qZ3s87EJew
8v64aynMXi1kxZ8pMMTiKSBYbqFCU+3xoaVjCWdCB8HkAXd8VALXbIym6PN2ORjDUY2adDplz0TJ
fceeToF8efRYhn2nRq4+JWGde9R3F7QXD+/fpJrAgSSp/g+hgZxKTjjw5AjL5jv5iZ4XHbUXau8u
h98kJHnYw+z7PUQNEY8aSIC3vuJrDlpAp/M7v6bzkQq4957oO+TPQlDTY+BWO+yjBdNfZQ/pSXhx
Zctq0AUwuJ18m0VouasNnSQ+ZfdYC+9W5GmHrTpqnx8znbK9fL3f3WE8Jn0YpEYh1Oct49F1eirK
jv2FWqNGyQX6egMzQQX4PEB/fq9ICbutz7YOeZ8m4wI9SOOJ46v7UJJ4eFFqX2JiV/6YWkZL1s15
WsfMZfesJmjqdyAoWaas5ZmF4X2q7cikDhi86/VRNVu7sRLfJuggZrYh2dfa/7RhNNJL5/maVEMD
1S6MVMHBaaGIl99SoOgXvgaaemaGShFMA4qCRbv6mT7JQOdndTk7p2lppS5WLWqlJq4JSq5v3HDh
JFcO4+MzVzRcguU5noL6MUGUyIAOyVCE/SnR+VHEKAfIe2Scj14+XcTUlfqY8RRKaLxpud6+YOmm
WefCI++UG/Cmrs0QMs38xJOkSBfZT4gU3zS+85ChF+w2a3DIlnAbH8GHwqgwIIYtMvTx11Nmj1wG
HCEP8Z1YV2nB0dbokaNHBl7a/u4TfmOkPLl7bE7pm4jtc4lrFDxx9fX6Z/VImmrv8702/k2XdPep
K2ZhbDJAOvNd3g/RT/xf98lxxsy2L7ZRPcKL5OY3NoYrjW3Ylwsw5NU/g5uoDvO9Pfrl+CyO0nMA
/xtVGZjvoq/Yb55f0L+d/TFNIlE5eTaAfbdLauJ13yEhFiFCvbj7rnBPhv2PykRJwgsKzuJwTJbd
pIuCUnvW5ZC+RsQjplsD4BqqRW3E4aorP/F/zSV/Mus6oSisCjnNmYiI8iv9u5tNcOH2TY6HMCt0
zkwGaZu4/m249Lr27HR4hiYTC98N0hp46NhRzwv2xXJaaNKxz2WR/F06+JsqyrxkRb1qU/+6UTVd
cCQKzDY+8fkLUzxKNMk31s7D5DtrxsGO/Doz3J0nsjAHwfT2WHEymZE+HaL0o1R7lG9Yqb/3Ff34
FiIdEOBNyq79WNJBhjtNny0f0bth9CAA8V+9URx0awH1CsM0rnkzrNHNtslUFSYv0EeJ612ZKKLL
MhZtMLrZYHqPUI6nsPNeJ+M30Yq8ufv3Mzy2+GoF4wQsoZrR+dY0QZP6QW36SPk50uyOLjUBEuff
MWXGUQAFibsVKhyOEvS+UEzQPvhVB9gR2CL1ySjbTlJMKnCu7YKbWcAWfisWB2M5oSCRDE477MtF
mOKDgkqls+JQlWJA7oTetbftINqFN/twJoNRLbT7k9IimEpnhKAnnc1blnVb88KzY+sLI0nilT7f
66s/T269dE/JTTxQBhB87EBO1paTI0ijDjF9BX7LpG3Mqf2/ZyF9DJzyUNoTdypgci4m6spWOrhS
sJFGNbbiLVrR4iHdFh58hm0AAfHx+Y69fWiEdpD8n4I5AcpA88E2eNvkHshsq1LotLONvhbHgFmZ
+Jq+iOOqXw4sHvtiZaVqoezmIEkO1850f2SyP0FIvtQtM1PicMZHW5YJx/s6xUtLwcpiftmR1IKu
NQgOdpQHTNJIRrq8SK57BbCwfAPl7jfunRB0u8TqTzNSm74V2AufpZ8rIjBw9REIaprBIRW0CeWB
Sspr/UBo9BsQs7B2BGEPeQ2wjra0s7MYoHsjDC7DnUH9L+N/V20Wm5/RCTPwAcAt5OkTWUOe52fS
wP+Il9usWgMnQkPkK2LRuDRtYK0OzO2YbukebPHDgWCm1CCLhDtwLTuTLCdGhSmWlwa6GCrGjx5p
pNBV9JvBcEbjvIYA28hJxkjTTdeS4xWdMoBpiq5ij3UdpYzfH6YBcFIauygJrie3iQGegdjfyzF4
QJeG7Hu9ZLLDAC7gAb3yfWf2zVyC8bjpsgCXXteKwxTZOtJoQAG8zUlwLtbnYqvPv7XCI5/iySrS
in9mFV2TlKwy2D5hipztVjA/BPulm+Zkak8cgeU/UbAETmozVC6PIbLPHgHiwcb+iA0dAWm7o3fD
UunPw31m28XGd7RjAKLRObzyJ6LQ91afUAVQHfMwLUsV/xjnwDjxvDR3Z3YJS8DADXZfNW2bec1+
cy8bTyX66h/aDFJvUcUwpghd52nHEs/bn3qALQJA9d3pFXolYiSJwux8Z9EGjjMwPsXnKxnnXg2A
MYx+bqV1A+7+Ei47cUYs7Z1o3P4kdeIJ6SJyLUbnYqVBD74/MvS6O/yuNF1EkVr3sjHJHG++gQLu
TWcf4rzWLwFv+pUh7IlY5ZXW6lly8ISIDN6LFxnhfK5u/QCjdCewNcfQpLgwTjHilSKWVVl3DeiB
ab9iihaVScB41prXdymmZW96DjEIvm3zEURjYK9F4003qYQqX8vpSDTXtlixbX9pkESSZ4iQlzh/
nE1Eeo66MPzs8ANtuuk9htEJMduCTLMn+6h49AHiZh8+6MvgpJE7BnSBHmuthCQoQBMqk4AXkKCO
jF3QEZ9mw2OwyfUArWxhxHWLG1N/AkhWT/qAJ1dngIJFzj3Qntx6fhtZY4YjDU8i8sy+OJBSoU1K
eUPnai5ViFelCh8LA5AJZ9onc6BY4hr50lmagzuagT8ik7yQCDszhBcaYNAtXstHKgP1VBvuLECR
0cp8Qd5aEWgs+8I4l+3b/36VwyN+yQbe5efxqs9EbSOXr1jcGgNAPQSdAcwAwCYn8PhZGH1PscZn
4aS8vMTQn16rbsfJCSl5LcASbuD9CPq73ic4qqHLa5E1QgWDn3ZOkmMaKQeN5iwrV7FiFi8b99tN
ZEIdIEZM7+ZLMJs0phZi/aOglm7OYleFlKfi/iZrZItnvZrTh2s8sDCiFCCeegj17wnAbc91RTep
PFIkJ1abrc8vQZtpj6fmRO1ITgEbYk+7A71T9cznY8iOBZWJUuSKcLb9HmDAhXlVJjMjMZ8WQ85H
ZPZEk8FmYlTqku86dFHpMr6WZbaTe9N/pQydSIn1hHvUoRWo96Z801gqzdjTgex1H2eMxaOqs30Y
trvYSPCfqykCSndCdBgOP+AN+vFb/qRfsSECRpDFSSs1OaogIy0nNzOvBs0YcLLNw/PlNrgy4mnJ
+0l0YJ93ORFjWERxp7b0J734nzczPSAcGvW39d0wjacB1XKZRRYi5PaOPqwQlxyYtH0raNr/Z9Zd
q5SULgocLJq+yAQmtr/wkgMM2iKjl4xsdBxXZOSvOeWKk/2vE9hOUCPUAxLuXKkY7WzcTYrkoQpo
kbgaTV8C7szHK6eNmG7gIkuXr6JRGrYjXpbwptvp3rlucN4HyAJFd8z3eQ346uOYVOQ4GSVPLFDN
1cF5EU35l176F52e3YY6iOrDV5STpXg3XPIBthneyI80h1pU1euCYUCbRoRDA7CiAIlkkn1JpeDl
NUOcr2a1gdXGKm3pq0PhgIH6XYjbSuy3+yeMRHJ8MBugPMlyFb56Eopc4USxG7j/BFPDSVcZKAD5
Tdf10CPlwaNleg2ZID/cilYewYs2ltuqimQ6lPyQvFJHSWEkGMhiOKzg90ZrL0Yv6F3GYeLEl/FR
Wwk66h0TGSxfL2UDnS9KFLA420CL9uzwh7M7lFkeoO685Wb/8PkxIFqBKjjwH8LlqBRIVKeGXr3m
jf1DCGU5yg0VsozB8cBcvULdKqhwNb4ULaM5dmETI3CnGtA7D2tFS/Y1nWUGuiQfzKpokCYgSiPp
jDUqirNf+pWEJTjqSLGV/XeXTISCU7ZV9PT6NR+ITdPKBVXd4nBWok1T4Rg9/n4ovzWu5U5qCFZX
OJzAmDVfK1la/MIsR8P42VU7y/qc13LumI1OYBwW9Yzgy1uXWdXZSHNRyWYcckvCMsmGFYcpyLN2
kpGSxuPU5C5S0eqztxUJs1N2ZIjjRwD8gAX3xswUpt8UYJD366y6rs8BddXEZkGqLnyc3LXVkGWd
SIi5DN937hT/LzT6/T3FysWYSC/3NKcA+FsfkifC1lj4hTs5wMNeaw82gOelZjI+gmT2cHEM03OY
gyM0rY2fDFlKSBw+TXfQZIk8gzT3JMFAyL13ub3rBNTl/Vlg14a5fzwD2r2DlY94YmvzBNMyplli
Qp/0g/l6oniDNcWRWjTT74N0lIupBnXp8nuXSxDYEq5HcvtSAa4wA5JUHo5VNOqfLbtUw/GPtt8u
qm1YwwGr3D/aP2rI9rGr/vlVIMnJNAPMsOr2ZlnQNnKtSeaJ/mzCdtxQN7AI+JcNViai6mP+VKEH
gYSNtOORzKxjOqa6VTiHubuaWaKBgwQ6y4o2WFqyEPlksEDPyL7X888RcT1Mzdl3X+JypkYQC48O
Q8PBGj9GniJUrOPDTadrzRP1FkZq4zsoL4I9S+sXDB6jMoAhNHQ0ui4uMxiPK4RQk3LoeHWIarLT
wYJBf7RQ1tIxNagLBG595n/IULwBfdkQbeEPihpDuQtZf1HJYvazmsYLp7AFbDy1ZOuHLk7AxcqH
S1PcgtWp/ZNCVtktDSJGCrwYCrjip+jl4h01aBgWJBme7J9PDLcqw9H/3pmqKmJGSoC1QCK2P+Oc
qWMTXAbcJR4T+doR/WVNoCdrirqccRyS1AMwRlPkH8GKO5lo//j2SsOOcl9nq0cSb64Y5E6cUd4R
b5LCBuM5YhTc0IArJsO+/7+iDqjc5kmPk1PvgebeGn/BqHnltjU2cmRrKKZcAOYAs9JSSr5fUZae
m+ztql11+N9ZADPYRDXje6RHDU/cCgEasxfqFb4cK77Vj3dYgFzpHVlVr5LSR5duSBotwC42wQVZ
Iu1ghuwyJnL6IBj6WTvU+G1uywbTutlFPZmy3C0e21oeYhaUopZQxUwbTH2I8Uk0Lz3bka+IG521
FET6e3JXvuLLu+Pc87hIsCCyZf2ypFXBr0FjuXHyq1LhgFmAhDwUct0wpHvJPkaUnTwDWBm7k07Q
G6p3vvo0ysU4gcw7zZfhZ73/jKcutVCZAKYCsbAYBLIWGslorfJ8un8XdndyuPPkvIP9QtXuUqah
t18D+xPt+WeKKb+rgJDhZQ4OhlA8WjpDCsMsQGdmdDKx5OyQpAMR6cOPmwpyTacv9EPR7Lb+uZaw
4WgtV0h6xKTSOnyvglNh+s8zErLmdfHr1+22yyakvvkdxn8We+sqMvnzKbi4uqQQW8L/lMbVvwUC
aaTFZ1LTkJlj6uixLkliIgGXMaSsR+IRoyB1XpLO3PejsIZk5dYEkOVwry8+Yma3SyjfnWerb7w5
9oL7AwR2xvZHIruIoL5Nk9gr3WRd88uqpUPk0pYijTu0XdryBWlvgMdmGOuZ95ekxL+Bo/QeVlAZ
Ch9W32liE/LblNQvxYMnYv7ZgXEYvEkau+uS+v5UhfgDEbm3SgFUX2cl5J5gFOXZ3bqE0UYq9qI1
FHoxSrwHRnGIBoabNbDozSL+HIYXhJWuws6jsn7DOuBqSLcMvuO3HGxVH4csi8ZsDEKIb4XVXrVR
ETmHCCaGuwd6DO8XiQdjzn0Zc4OzToMtUAECHpaiBotm0B1/o+YJNcfNbq6jGe2n0OwsvuMKLoN/
ULtZ2fIz4+O/vK0Rojsckv7pl3EqGLsvH1CxkcBud2DVYfoi3cyLAeej8i6mdSYSMug67b1ybthp
3oGofeUEZZg8CUudf4cj/+nRF+WOXL3TH337yM2UWFMbW9hevoP0yip0DYxs9XQmiP9cV2Nhz6IB
LdjNqdAY3R1DsSqMP7X4CXKxeHJ8EfhLKLc1tophl0QvL+WfZ6qDMp+9LIWZ9pCDjOqqK5OUUgFQ
FV5hBXOXbDocTD5BydUWF9NJDJvI5fmWLJZpmsm1paN7WQSvQlpkGoH3F34yN8Jtx3IAi3r2tDSi
eWw5feto52evemg5h9ZZi6QJ7TDTlxvl24P9HH2lExmMGqFBSSXoStXp1BGDxdT1pXa22NEZYyTe
b+F5Hm3HzeU0h5oTBEepUsPJ/1vx/ETbhI2yQWgyZ7QxIZA7VwKIH+q+UlXwGNweWUnwMzCG+Txa
XDsw9kDlKwO/eEqF07dan3W32UVT4C7Q//cq1c5/+Pd9RTSFmklAwUe+jYwj7KnHCagkS1smVTzo
TN7ysvqrgXzRdpJ4LFjBqZXSblwFpYXIZjPiDJ1WE5cPrB3LBr3ZQM7pY+42OY+gA62Zwi0B99le
IrnNRwJS5NWGbFMfIyT/LEexAhYZ56n5pS5u6IWuC9HoicclISd4r3o2+FhBLxFZLNPvFxEDFomr
OF/eirXqI9/50bEWpNZt8rBP0oElV/6eroPHZApVG8j8V4WWdQvaQ0tvP8PCIJBg+ZSiUFGGKwDU
CNU0+9zoBG7B6DKO5Xbt//vR1yaQbVb/iVHQajieoGQedG4+SEfcoE0Cv96Pca4WKjQNUIwxhaCt
hItm+sl/YqYhWPXgjBwoi10n0EpERh6A3nvM9vxh6xcKWf4Lk+fepxZ0MUvCS3RiAIZzVyeOzf7N
LqvA6Hv+mvnYESjMctyG6WiX496MR2lFsuvCzY14nmnY5lc1cHLBeXT2+VR0sR+vcal61vjVjLir
aAjanUnVI2i0S1J/IGgS8GSrE/HFYyrnfrf2SkU52sDOfNwIthdOO2wnJxXAJPHHmLRyikrUvWGy
qPd3/RVXdTZVkSZCwuBvSuBwIPSOVWez2+DZc7DqltCJwzkJwofSH6OSTY/EWV8uSXwPAwV+Ri3A
iNUhnVuY387nywxp6HMaA6s5v61OYGPr6oBQEQ98kED5UqAahW2kS78yEcvOwPDOG2tcOEbESlR1
WYIQCPBSkHk9CCTpA7E5R3uKCmmP/oYuIzKvPGfdiF22+9VB22DhOfqlrv2rSAD79CoUlbUZz+6C
ErZCXK9zV8SUsFNhM+R9pNw8uaQGy33lP605NpfnllTG7YPmBaBHSWxV9MEbYPmjL1URXUBlEIqc
fR9J6kiDMQ6LAfJdl4257g1t/Pu0R8c9HO55pfM3ORE/mTtb6u8LkcMYrfPoIXDXkMP5l85irG00
D/SR0/pIpdUjZGAeyRL9yZMzaw5eKyws5iC8Ra78tNwb5V3ALIgHHPJfCTn4JlRrIvwCiusn0jyK
KJf55kLkELGjXAhfv7HPAGyKWFIMQCeHdbo+5RXboRegm4gwzIX8dLVny8xt0DUvtjalBP2djB1/
uerbw0eHg5E0m3jmPzqEGU9fGcj34f9KRGZ7ZLlZ8b9VXzTsbqsR1V2ORS+Rcp3LJ0HfDozTOKxa
hFxpDVvz3Woz7Rzzqcf/MhtN4VEzC+fEQJm99nKzWwbkQxet1z7hfR54bEfJw46DwPPSu2ngBoIf
g4gjRaeWlQx4HKBaTl+8yIBCmch7xyr8UYzVT6l0VPIlm8uTJ7ThNxtqWbrefWeeivjiIRnHGEU9
Fpa5cONxUY+FTIGk0Hjus6e6zhzKhxqklsItVq7lZosNE4Drh3p3jtemlaXaXw4yPoOhBn14Yodh
SOQla2YAa/4K0AcW9Nn3sjh0Jfo7/tws8/i7t+HMNzyK7fzF42zIRvp1Ofl7XxE2ih2pwJsv5FwR
wtgOxIBCxY/HnFE1Rty+h4qTmupTsQ2zLAZtlouX2sClOpNmXrLDpHVsKtpUrXNjnugZRgE7VMkt
fGdPrIOPt3LGISTBdyOjrcLl5sAYZ+y2H0qQtn3UbdzqekiPlTWBL2v7btP73oM9PtF9NKthfKO3
Xj6Cl/1Ol6KWTiZCnk2GOSp+9017PU8YvChR/7hMHjp2Ed/tP/NozDHk3N/VzxosDDBytrHezn6e
V8RfSV2cxXYXLkt3WaIrgZ2os5lbvtcyVDTCctjbmoLlLxc3NGXCWeCR6+JCX3xGsEx8VOFJDhb7
qIWuq2/O06rWrEz0VmA1gmFHCR686BTS6u+iHv+PyaYkZic5MHbcDM1nNldKtLY2mW68leQ1okXT
eE/GukUvKbSNpUT5F0x3IfmNfFboHRbCe9dZC/KjLkvz4JZcXgICWspt1M7nTJLEy2GtcgNR6mLQ
njtby2uUK/Ysvg1bzpC/yy2y0eYkW9JPPPMF8IQi2UWRihlb32qz+CFmk/qQqwFbXIEIKH0vJK2m
GrysBTX9TRlQ+CO1VFAjmBllnw+vUc+Gn7SPnWnL8L/Fm+ToacGOzDIDXUyzlFO4vx3ZRAdCrxxV
osEwBiVJb6QM32ASuiayXQglbCmVvIa0UTyhh55j3nuY/0yZIxJVy+P9YowSf73nz4P8fHatsyGo
ViIoPy275PJKWPnbJaLi5tN1l/chxpqUsU51P3/xCUOHEqm5WSzWoy6Z7WpBT/RDi4uQ2eoX0yFP
6LZhN2ihdbjKJK5eK5bQymU2rDRhJSFeAh7h05NSdhzYLE4woXWiC9L7NlUA52BeBI4JZ/DO95sT
M7UrgP7lHm/AO49gzIjkTyfwiJo7uHLh5DPDgfX2NUvkO2xt6r45Xk3j6ZEwkJNycXOrByoXBzxk
W5muWve/Xftx7OzHGOH9sSgrs8Wklfta58ZnUtFD71K3NJUyU/C07WLmhTtvaaLigqx5rBCekZXN
n70Gw5I+lj2Wi3ycn3GSUISPRdoDtWscb3QnUqkmLlzgLY2LbEvlUAwZkzvYHjWLkL2KDOx+9zmH
f72RSoa2o3vozJywuHlsnHN9kCFNOUJhlKTbcv13lbPFJU0wDQejS0qguV7MKPA9qXB0xJUTSPvH
YPPpntrGP0IYZyIatG0VWzWS3WwFKheQXyvL76iS3XMpbGSx2ck1ihqfZdgosXXW0gFUyxgeWqxf
IkBoquQb2vfmNFQUNV5oqkIDtBbZ2ONX6Zl00ri463ibxDhlvJJvL+QdkoL4g/swRe4XOQDkaJMG
vrGAa50mTTxukrgmnGKk+AMMfKPVJgvi0smwNl6oEQq48HgFUb6Swyay/jbJuDmO+epvH7DEs/MV
Hw+uGYSJqgS2fAXfkdNgXJndnZqK8xm/wN61kKTP9CypVc7dwKgr18+x1n9PX6fS6nz8AGnDiVIQ
BCuyMdxtfmIrmQ50j6eciO4dKoggmHxM991JzSbr7DqGn98Zi0xOQzqfcWDhXzOjS9lpRswMoMKA
g1E2aEYileuR2N9kZ+Jkjwc6yK7cSpxYK3wtCEZSd4Frpf5j3hk/hjR8nbGTC10vU72v7YuX6fOm
soVG8sIB9rfHXaSjeHCzzq7EmsvQ1NPiAKbYdGaLvmDLIFBz/iw8v6scYFhtGNHxhSEj2YjdPC5W
SK20fiT8NJyzimiKbpeW1BFVy+WaS/awYgQGkMWIaQpnRnH+sTEJYDVczNwostFmEFsqTks3DyVo
ODlLswCuVxhl2ECQeUQbwUqJfalob+xdGQF5mUmy/HyETLclPJElkcPzioXhy5pe8ReyK/piCSbM
ZfV/xwe9y924tdwhBCedjmVKrgTXoeyk3OKeWG0+mb+GZ6lj2bdoYpQF7lQIRcdJhEY6NvepJvO5
3pf4Wzas6lBgPLyOQlA2dASRCLM0yqpJn5Ofn5f/vfnka3LSJIcr/rIAPq5gQlUT8xwmBjWTJ/yF
TBrw4+6H9uf2LqiRK+wFuNkqENXhNGvvhqYjo679MLxuxKj5gbBlJvZMHmH3Q73RCL0f7iVa2Ks8
FFYsCgjfb5WBLEdL40PioOCpiV5TQUGxcfDCEUwaRax7rOft8VK8iqndyBuS8wQ1Q0F//2336os6
7dVsRLBzENFZ6SSGI8OTwR8Rp15zAfuKT1cemaIx3JleoXk326y3FCdtPUfWntjgrkODIq57Yj51
B0FOAuXHq1DjdsBblUvi4i92rtP/PZgeY9IjsttspVchXYnGOBSHATQm8mLbzGQ3XqODvNW/Trph
G1eAET9LmvIrvushuGW1R9bLErOaEBRTK4qIcwGnTbRENCOGFHArI9AnJUxxohZ1wwutoN0CtIlW
4wDRgPPNB8hcEOu68zD416g+7ZCzY6j+ZPlJ+S2RzHelQLDcKj8NauNuNv57pd9JiMUNsba8Kzcy
qTqWjuNMF+vjEPLaapPrQBhHQpVldt9pGqAueZH32cdI+0vwXcmNVlp4mNj0zFwTdVOLESH8Ec44
7Dj5fZnlQG6qhkAanzLtShPJsSDi65BdaP3g70If84vg+z187WURxBC5jjuVUVkfxyCAAZaDukNK
XW2DWpjo5uKQteSqNqhfxq+KlSTrqLoCu20v7fxj3IaiCGQvjivfCaSuGLVWdSn7ZDRnWdpWFyuO
bkxdLQjcO4LsCeMYUAiN+Caz9EiJYmFTNeT+remJ1RhqkvaE//DU5ZBsxPFTDCyl+fyH9jZpWcem
yxI8xzCYFly7zsWEicdJhfmLOPeFUtKKM9qGhxuR130DDMPJyx71pTNN74bz2ECI2Mrs5f1axMsr
yK0rFiBYgf1CrQZnc5FJKLSbM+Sxms9EYqoWOc/WlkWJvkIFpNQbzEqcKlHvkC754ntjqqq+mliK
MJeXw4wOPmvAQwAZ25mFtdO+XI6kINs2AOuaiC0fqE5JtQ+hApjiPXKziHXUL4lVfbzKRuzE1NK4
ogSsEh+pwSd/X5mH2BxY/XD8j3558l4h5xAcCDvWzPNL3ybcU8BAwoyb5P64rg6FSq7TcsLJYIRK
rR6h5s6qrYDMacAtHAzCYb2za0kIGl4gIn9WRvTNLcy0pe+HtPVUzAMv4c82uYpsV9UzlCaFMkJe
67pXEiMFH4OUgSaddcRoGzOqT8MghlkELijJ9jzk8CBK/4g4QKeSjkH/vzt1Xp7lQVxJNiHMwpjD
RCsPrfQAYnTy+6PtITRGO+TzP6xHxMAVvWRy/lqoN/RMRYXBUKhrdVxGm/gBh2IXAJMDPul1rw97
G8r6dE1QTssmG0cZsckNt7iC/kyriLmfnRb6Pvh21j88UVVychd1YjYlttM8I7oCL9WUEj97qsgG
PRkvbTlfqmhBpWG9OEF4/KnDbJK0rWnBCapTJ8/M7klAGDkGBqm+LIxA3HGWKFbOSAND9hAKOPm0
a0QlnWlqUbILjwQZkIVEDyDxkQmqSUEtnyqUvcXcEzjZ/HTww5o47/On8M7R/7S288uw7BuVBGzC
QeiRNnN75YkASTyAuGleZ/APNnSzVCxf+tuG/kjxv5HF6u7A55SCv4nqYbxGW57eOnjjP6C1ZseN
DpFrIyks7nlEnvm0uwjK+LJ5QXL0xjRi5TVvoNwqv5fl+yJoy0iKZpkY/gngUxvertjZjz+g14yq
hq21ZR4gES0LDUgddUwnkayrCdYxaSQFu7F9U2YJRFU1gabOQChIyKcDhRS+rEqLcTBeuvet48c2
9MyQMIGUzLBY6lfrIQUGI+J1Z62IYdTz/3Z1bSbmOT+Kx5ZWXflF0lNFlMLdfqSqOtDfaOWMY2fk
O+vycyMkwrt0vCidjGzT5J5RXpRtPQ4SJJdpftfLAYBvefgXiusVxDjESo0in/I0/a4O/8+Uai/r
NgeNsAQCtDGDj0Sf8iLO7FFiwm0adJS6Q0w5fzjxygTaZbUnPFPBVu6hjkeb+pRdfoHZJe9e8MpI
9KXqcuI8T2jEIZn9L9KCNhSlPzJrDhzBvEhE7fV7WTepH2H6dIGVPUGOxdA2GDz4YcMjCjtWTmOT
pVkBfWtDYynabzkosiwf99u3xLWV7P0t24sgklc5FAqlU1BfZd+34wvcP8aqqE1Kqd7M12q2ojlO
2aZa8ujNkWmng0pc4Icl3683zBZ/2pAD8+T0cPjVp/AHp+gkjv+My9wPKKucrJ6Bmk5teHy4Sh8x
861ccBfScbuuXTxVq3SapIoiJCWHCsFOhW77Em/xJYw5938uQZ9f28C7YjUrcOgQbc8uUgFZqUpj
ESPj28tonfyWIlvEQpYl3yvWc7pnGmhKtRWQo9mht4/F0R8kRdjp65crEFEsdyhc0Z9lZuAjplnC
LHeHgiRijk3oNxuAiUSMsfZPiINr7Ab9dhj/m9S+0VJZyMSWF4Q5Ty/lJwKWDqiJsAflMlDlv3PD
VKewYBBIiSnWZYKsMQyEYvR0CIihZGMT3zsbiQ0zqWTh5hRF1WBj9FiHokqIyAcEOuUFvIGuF9TK
ZuiCcIHdvpMFTS39zkulna5HJFXrVXaIGMIBhb00n/C/ObMuMiaCs9Wz12Cp6OWKR5VKxWwV2H24
SYavGfOuP2ZZpaBY6JVNUk7qHW+EN2Kp02GxrLXbkU6/vCe7Hh6b5DpeQ+P4xPA+oDxlPBveYQYm
eSXd4ORAN3MPT1OiBvtv3XHiVjtijKc8PDJUtlA4nI12cHKtQzPBMCm5Kx+oUF54odcdM9yiXf17
7Whd/lUIIyLyxz4t5oJZvEmW+pX3z6N6GaV0sP2k18c5nUJliBhII04Yjo8bQjTG92nJrjPmoD/z
uM4bz6rUn77u/YNwzvYSHmE8V2nj+mqm760WFEnKDfdDcY4xKVCy/LGttL9mAxnsKICoOyhPQDPf
lyQQ1rh8gHrFu9wLJj5j76hdeCNHu3UA7Z4cv8OoHskuRBxAF680q2/JqrmZVM47TPzqoAunY8P1
yy4nBApaeLGf0eeT1f/CORzofcphAcm9BuHqDsT25cr47zo+1hQBHV0XbmD1zPZxMYrXgPHq/dlP
tZo+OhpqsM9PN5QG36Cxlf58sQTMdLqH+bKw8+Jg1jVehgbtXH0H/hhoVvIkgooc9lvuJbrftPF0
gpIABOBmFWjLn5s6FIy7leZXO7NwHwuyvQQxjNP5aBCa8+UkqUpq8WsrMEvL49tvpJbMQZz7Vt5q
mCUrhBxzAnpcYgjzrmX76u8c6NT+rrBTVTAdkzW0oTimAuTRQk7r1TNzx3DwekP47N8uOLjdI5er
Mkt3igzeYP8PBG14OJDZ24PlHwBS2OHaOxpQ0L6CsbnMEkNiUwNZ/3Fa5pQ4ICJHuvL8twsioo0h
nsp3+qKm9LXbORuGST7T6tccxM4JYoS2OG+Zbd2vIa2RlTQ0SydEAwOzgX+ojeDI8zFf9QjeByKS
xSoC4fL2F1TwGG0sVepg+V6+yljd92uNYHeRIiw6HNWkI3IZc6aTgeomMgkz4RBIw/BOaYVa3UDb
NDauNLziwYSJAXbHMpXGJU+fZOKUV3yfLf+Bvk93Um+2MELe6Bv2zrw0qeXojboOphjmCveBcF6N
DIADCDqUhamgHdnCmLYgs6/JBH58uvQG+ONv9ATH951dp90yJY3bt689IBdpRcUUAvaMQZaJkaTB
IuTsW2dd/6jQKby4Ic9clNEBH19zLlXeb+i9u5m+YLF2GzygYwGwOyC8bNy0aNgTZplcDfeCQHnP
C9jGxVQykzPvb9qPjKCO+TKkiXAJeDloA+9ZE8ADRNjsa7RuUf1cwoz/5U6oE2vcaLEVLptr7S0W
hoaxhsx2xG4YPYM9VCtd00/uI/mBtTmcDKmG+8edzuj0/3ONcgqSZ/JVp9bYuEiktPJ43MBX6vGH
kLrnw7Ci8FVmE6eUiGy10RTUwGrGIGOyxGt69JikLNeCsAzFfjOXQ6KwKJlKxhmTuEmSyHSk+1XS
R4ip4yha04IWMDJ1gqN/BYvRNpRA1zCi96eNidVvk5f8bfzS9TL3lFgopqD6oH/HbGC7oEQh74a/
/qkgvB8zTIfDkpWV4zGQr8nzxtESeYlOIwpsNq6ggF9RO7s/8kSv+4jeiXrDGy7Ajsg5BZYfJkZB
7Ud/tNf/ImSOCFvjHgAcDagOxvsE+5DXrFPBeSfkHtqCHddAF0ognqzFTeOyjsy6AjAM0XOhmAoW
uQ5NaR6zmHk6WNCcsFPkOpbSoLYtnQlp4ZQqRhtIHuzcm93AeMIiLl9DIhq3FIwOIvhGXl8H8GUU
HSmKn9us9XF4GmyBStmLq54z9TX8VIx/d+6aBgFORHxhK8s+14epwwVn1g9dmtI+urqfdu9Qdw6J
JB0XapoeHPMHyCyxNWyWXtW35qLyeucg+IxUvbOqiyCdA4T7s2HWotMRzR+1kXMjxFUpvGqcc+Iz
JcJuNHpbSbBVgGOmNWh5HfPnI3T8rwdqK+zLWNOHxnWAVerN0DZQWycqVOiNXuMhH2/hi+I/hFYu
cvRlpRA7OfBEEBgeMsTYjFfLNUrwbWLLWXpq4cqbQJkJGse76fiyi6yXsBjZMS2h5dIhmfjmFKBK
sZL9TdExRMDj9FvivX9w7v4f2gDhhlCeppscakXl6jarFSrGpiwJaEYX6C2UYcPOnH7M72Qh/10f
zmLYOvQubxr9K1J9i47j/oD7EiUHjJPwSkynl2JH1yJeHvR2J/gGlCXLbrfDULxkP1aEHwh45VgD
E4BcxHm9j2ZbjMUTUYYUuEjRp/jjich51oBBcQWd68/N8rXAauiS0UY0p215TnZKtdlGHDibAxaT
dmgiaYS2yIEycJAKBhhx5aC2P4EByww6pFU5J659saglgfbeqL9gQBVMcBogbumhe7pkHdfdcjXB
FTtUqe8ZiBUhT+k+v1iB+Ajth+2eWz6K16Wsu38LxGGJOXFIbXAaBZrL+KlnJ9CSK6AH5y9xEOeJ
iQmUc7tF1dLz6aftIO+BUGGZOVHbyUrZdGwZqBNGtHkrO4KKu1U7lD9lWiAl2jGgwNL36Lkk7fk9
lQsm2IJDFjmDcsqSmd3E+774tjYKqqWtFaqclg+cB9qZoaZjuMY5yOasyEtNM50mW77+ncchlRyL
s/Hb83UHc1NvBSj9a8vvN8vQTqogBb7r1jxASIuCGo6nM5CPh5pkzwzmJl9w3BxgISFck6069A0u
k/yaAW4XZj19o763aDal5AgXV/iYluDfexxFrw5Xs8jIPcC5ODPe5HVb66c5HEihXseWH58hukgb
rpFdwuJD/hWDXSDflhGrB+4Wv5I/AUzFDTQBJ9eBZqIDR6XhHXx868sAOBffXXmQi+kfIqq7sVn7
n7n2JGnuPxuAfR9wh+/ywqgXKE7tLrw2x4ltbVIlR01tFEYZ8lnpdZ6iOCqUQof/dDL1TWKz7oSH
oEGhjCi+rqltv7F8lKy9qZS662TCdoOTkUmF7EmPDrdf2Rmhco1AixebLlxghbVpj6ZLQrWn38nT
1W+KbhxBkjzT3GiTvarYwxO9WVgO7d5My+LgPL8b5kiT+7IFmtoRGjG0U1PchI+0iLPQ2FOQOEFh
5IFvluPQKAOvd09zgYIqzMyIXHPT6XEcQGckwwRqFMpZ6GS8a+Posa5uZlmHxfYTemtCRzMGDGY1
MAOrFL2/gZUYkcTpTnCSYEOlK4C5nA+hdLKY4bnMgpbu6oin2L1gNvOZEM5dklcqDI3AM5nU2aVL
y0tVAhFGJcSRcjwCv1yydgxNYhbmod/uyn9NtQvGFDznzWDhL33CaA7YQK3HC17qwBfpQ39l+kXu
+0lmrvNA59LcRyTHyuqW7NSCp4cZYWDdqdavwURwQ1o0duQWkxWKyD2hPkGELPAaU9he72MsmU9U
v/WOc/nmomjxy/AhQd9ki5S990Vv0A8Yzs9NrMpR8gx9wm7uPKaFm3Nwk7LPOCk9+NCdmZy0pFL3
gFI0uFFYMpBvSc1SmUkOBtN7jtW8VftLzFRitAp5iGz5r3p4s9X5jeCY6Ok/39yi1cwNTYnDkmU7
eqb6JGU6CDhHynLGBOmCUGvPvfyLR2MdkSEc+JOUCfpKgHqifPX8YFsyf0LiG/ch5JyhYAP3nCeK
wN+JdIQuN0UkoxOLMVgN6uOct3KesPCSgBWiKrpy+b+NlS/VE1SjX37emS/2WQUxlq7CQ525HZ33
a3o3+BgaCGKB+KPC7szyVBoG9gsFuFDhGKFIyLBhqW+QlMWcF0EJ79h9fIPYj8EV4SmXXF1KiBRl
lODf9HKfAqULVbzWBqhXgAzWK8BWKvo9aaM05lq8eY1acUPt17sYpzmn7sVSXY65WRZYbbc9QEFt
6UcQDgk+cvXcdJZOfh4xg5lrozIEfZr/4u11i+50D28qI1LMoedzQ1eI7HpZo+46WWHpMJRFByxZ
6DQQkpO1ZCbMmyyEGNH4RhTzUhcl+/8A1xMD4CQ1QfChHFSSuwSnLvu8n7AXtC8w7+v8oge7Ba9b
TzquWqraiUB6Oj199hybdN5lCKh8akaazc5t7mzrZc4ZgZ0SOXZ+8cBORnIHalDLJn4+la8yyN+b
3vqewSGArQoZ3j5Mm9/K+GxQoGjAH99ULkKE2wKcnx6sIqQvKeflctGHYhOOZekYUek4QIYN77ya
nj9yi2D9Qg1lS0ghy17Rq7jDqhZ4t00luutoTXdMZwRBCySkyi+3htnuygSZHbILh3vtEMMfiZi7
P27/zI0CEwOzxSqJybbzo71uMqWvsXiWdLeLWC5czMHwkVvRIZKLfY5XtpRlITAkvQOZWv+L221D
n07xeMRO06CZf2IhxhHkbdNkVhjCaKRtRDyWxDd0EX6HuFo5jpPncwOaXvEiqGCpXPhuOWOTg5t2
E22a1fnzyB2K4fRMCFyjZInvDEr/WBSPbocnTRLmxvRNlpSoh9Lb5rtYYa9RdgVZy520/x3BiP6v
Z6s3CFvy0yubVFz0yE+orTXr3J8k7MpTN/3wraWMAVgDfCtSCpSBzAMf3K8P/A7NDqDy4H1v/uTU
eJfhjot1M0TjZyvBAMC+yhSYNPwIgkjJtvT7tD2YWVqnVs4QAp6WTypLLCp3yAWhWwAYAnKKem5S
NAM4d5tu+F7EtldxnreF0RbTEWvnNjRuK3C0uk8+ITrAlmlczBkSTJ7HHs1gNJ21brKzhKDutLdi
P8fL/4VhoXlYaVZuQ5AeMAPvxOJVVh1J9OX/kD6U4Q4CntJTbeQGHvbnVymm8mjRYUQAwwbZq17y
KiiQubNvEO0KKmSWW83EGpSRlhnh6PPNoTi5O6vgh9VWDqMtbSYZ48Ez2NziBFGLbrSi2pKD89PD
iXDSHzL5e6A3qPmtFyIVDIUrr8Gm+6WgYoUsXeVB12wLcfrjzR5OGOXDR4yftGwbiN6DRPZBqHA0
7PZI/vJ1WXWqNqLeztCzUJbGoNW5o7VYb9SxcZSOV9mCP3wB21hkBdTyO46vLRxNs7nlgpz0FWdw
RDmBTuI4CTO78Dx4ZIEGEbNRQuGb97xLdZhiO3mvPbN1PrID+ZI1CRI3xVBdhgao2kAT1g69rpIt
isjjDW39oOLyYK+vEkh+Ks9gYmFtte80DOQGBqY2hlEbddYLsOhLOxosM20ZCgRyrGLTvgt6xThL
AziDevJq1OhenKz/CrMuR9TQWflUNz0nXUHiAgLlYT/c7KucTGMg0ZS0JzhYArXJVFlHe1wiC6HV
CzqJThKHl9ZiLCkK/nR2sJV8d/hRAsVQoXP2AFlCvRPaN46RFENj7Mig42a7VpkdZn5nNE2BcwCs
Abx2QHYQa0DncK3AXtYEXNiVi2dXYFY/x3/n2OIaTci7VeaHPKOzgqeu3/DiMFrDLlYrx1pF42iY
RI303r7TK427v534VQtKFYRIyyiRAZI7eNeotlTY8SaJ598obaVjYQx1W/oiGZo8t16sQpipFlOA
RRUcpoYSE9xY2J6zUOOiCDyjy43lMIcBna0b7vcym3uiXY9TcX9mF4gjXCMUIUgQ4skhqslqa8qr
nBEZlDhkInHZ6eSVhx7JGvRx/TbiqDsAbtwg+HbbpO6AHVtGie6YHcIWfO9bLwOKbXKMi2IozmMl
qZNu5Wrd2LKOTiTkjXY9b6InCGfu5zw8MCVgT3oIdutq5F0K3PS/RBZDHlO9FWC7R2Wf5cWt+6jo
lCdLyAwjmwQmEkpDefeWRmdnOnYV2clMnDpxICFYVeiNJQnLJJwF3Ylbp4mU/ZAYv/Fp9lnGJZN/
yK8xWr/vRcZpdur2zn+pQQGQ/sgXAxkcritWmA6yv6SXlhljRLxdnQRKOwOJQe0APNq1Vn6wlyH9
GF06M0b7V0msd6tltgo4ktAHyf7mQKhUnojsmsKN4M72/O/2UBjW/xvlA9JqoBnzQs0kqp5mbAlv
sIxgEMATB3YaGXHEjHTD3QuK2d0bbsNmEyfpF3i0vKcYMxczvXMU3/d5mDuoLrLxzB9XUNtknMKN
nqjrJScGQdhORcQk2WlqwQ95MXZBO9CuHoBBjL++BDrls9JC8eiTgFu69XnhcNo8N+NCP3yCLjsb
wP9LuikRjpVXY8q21sBDWnhf3gSn4yqaa8d3620ug/stBTlC2K3BV96x2M7n2DvTEFuZOTdpYoLb
4i7Axpg4SJPfVZ7yAktUReeIG8P1Br+AEnWz88C/kP25B8iEGKhm+nnD0OzrIAXObd2fys2wPyE/
JuhKlmPUAF4DeSRaocKSFl6EGhgHClY+fXUXE4/FCYkX0YTLQ26rAyyYypDgQGe1xl658CAPXA6l
/wNCEIHi/x1z5O6F53o1rpK4Qgo4RUijBeZSsclj8R+50K+p1Z0/avLlzolaplTeQPi3EyLcDkAs
4CBehs/jOBuIowTWAezqX9Q202uSPknn6XWkbg2nj1e0Fci0UumdP7ASJpmhNFLm2mnQeajW7TiY
fDTIh3wudNW+j7GYi/A18ljJ/Kb5FdEEDTauYlN1Q3kIT0PWalPsn2qs+MbvfV9/GGxfGDj+K6ka
qhClfokH/2G7a8zbuyoxb2lD8+gyXlzMXUpXgcY9yREQR6oC2gDVSqn9RA7T7biqvfyjrz3wjsAG
FfM12dB7+/PI66VuGQaRpPtnO6/SQY0AAEy38OeyQZs+rxN1DH+Edqaw3S4PCgEEvQmxuF0vNdoD
5SffJRbvj9sJrQ/NLHejil3oh+/Gh4cr2SpAntIkT82SBZcSxSBG+31FXHNmERT72a6jUcJ7JKQG
ydN8AN8bDLlkHZN9i9M9o6u2IIKbc9RivjaLMqdxtAgfHXu2zR0VA7167t/SO1hRCTFd+DQiXGQB
V7ojFAcChhkr5kFXwxoFTCLngAq4o+AnnHxTyVXI6uyjnLMpY2wx/khGO+HSkoX5cd7UcaBw/0r8
imSbcRXcltSdAruY86jwDj1kuE6w6TLii43HbRsdFHMgXQHoWJ1fa2qDUDHROb596zpZLUhQhGS8
xvouVvH9Dx3inKMFGvjiR5j2urAXEjtPwpkSUwEfVISB55ZOum3SnAhtFxBMKsgMgQtS6HG7Igzh
8pRgjp+kftA76lhOcgAYeIV+j0629D476BrbcPErZkh4TA4vlnKqPo9bJOa5xHijnCyxgr9T3VbV
sbgHlUBkUW3NeE5tXaZte9+9WpK4PpvWPzjxLTlz5zD5H2UuSouvA/Tyf48U3bqgHNzmhxTvNTbB
JbRTTVx3C88n9sm/BGX+TUpTxDUzIhjfdE5I0xGzuk6VqhsSF5YtnJM74r6F5mV+IlkGIRjC89/b
ubCqOPgCruTPT/DeAnoUlpHkBsUrRU2dymiQFe+5OJdiC/7r/gAp8fTiIQrWlxkzs5fomaqpSW/G
K7eMbAHo3pCMmzrEWnEUNDZ/e5qbzg02skNnwCAqFYodMJKlqkRKvS721hRs/bfVrJeW0fnOQydT
tGrwsOd5cLqDIWpmX08GxfucXY7HdPEfYkajzidzI27lOpwskAMtjOrW/fIU3njWL2yYcYNZnCIg
ZOh4dDG7+lhIU5bQDD+iaJo1MUH87EISDyZU0QkJdfg1yXIFpCng5mF9bvowpr4NBjX3d9NqavZi
CtuzNM/R3Gxmrw+VgtDV6Swew7yMDTzlvoIrciY3U9gjqLTZoNQRZRt6UgU2crFFwIfpN5qLC2Ma
lNQ6DGaEQtRIVqZDMqTU49yi7aPIuxKdFvPoTSb9RdtcV45zue07BHS27ZqHRAiflMI7SB5l8a6M
bsyw4eQh8/FktdKJ8BfhgmIgLBjRBelTfCTnIpH9WIpGgz/fdPo6WyaSYX6WgPgaOCoZFN13EYxj
FWVyGZHPkE7D+DkDbmnVDdqWDjhWoHJH1cQIorc6f0x2QkEEeN4Xq0+HCnuIzzKy/XauizTNtzJe
E3L+Ym1SY4rcuSPX/SFPgMOdK9txm1866jRV1SIRRcVKbRW2jsN0hRNQGNmtZ7Dknc9XDnZgXlCD
NNUAYOphvmVs0PbxX++Eu7tZ5eO/+5YqM9BraXFYySC/v7R3jf/cNik4dMG/JaIpjkEkSy0/0DDJ
3xaLJoDKpTxCL1DXcCxsysag/CF0vtiDz3n3ZXI5zMNKoRTzSrkHhp2lkeHW2o5Q9fI7M0qw6AVN
0pu/QRo17l7DBCRahq3WFaQgIZC81ckPTlSz1lR/Ips5g+jktbjnhXMc41K8E8pvQpCSCpmhrVom
JjLvNdsaKQmoJthHxcRgCICcpqFHqMDyzPdp/KoDwhOh4v9+UkQlvG5+gci/Qkqez05T+h5CZUxH
sxWWS99G47R4CTjiuz2XZPHA74r55MEZKy0xDulgJWiheCWYuaDuFghksxiz4LcE0nmhcRoo0lUo
FykvtHP4QkdG9vUSKBfLZzIZSDo66giqtZtrOGVbi1l9cjPkJQCYTc1PEv3QBs/142qnBAXciwKX
L3kLNAoh5QnWoYPOQH5AaasvPUVEQnEKJ5WfnUp9Bbvmly55pFaJsJn40L6nVVxD5NsHAMcq7h7u
T1ZDBGhpau3IpSoOe6xFSQJszeoYT0kMwuTN6W1hFvGZ3X0wiK1fPdqPGmzyWWu2qEjsVpFF3cS0
shC+FYLJfh0VeHirct0bntNr0fe67X+SDGhQaZ9CtkStjZby93neEAMujJmQ8dB00uEvXJ5uYt4Q
2JhXk8BgZ2/SrQcAPOdR9u/A3aU9isPwsTgLTOfFgrkIk75h/j2dg5p81S2bqlPAs7qBexOJ2FLW
48T9Lm3TsqozIR5xQo9uHqzkMrhIoqPIc3+iuEHUcdvRWBNVk8tjdt6ZFYFh0PsOK7xIQYebzx4C
C89MB4kwbQ/zQoE4kQa2TSw2FCdnHFi2X4I4T5SM58rkWn5oVwTQ/5pImoMD1MlvBliEtCBn5IkJ
ljq6VQyz/u9RsF9jR+SFSv3VC0A5B0lppzL4S4s94siBPKGPfa47Pw7ji57kn48hkxrBVfGqWLTO
/Gjz23cM2OiYwDxtvL8Vc3ITPfRNlvyJDyu/c8wl56T9YY/5ClVy9AaDt6Sbi25fkcaCNGSlBtlE
i1078fj7YbmKUAlsz/rdM6S80le113+6SXXWrgmWAnxwcvHeyk73jPJWppmUeku5HGI3Zo8U3ysH
jxov2tTjf7+F3Qr43Aj+i+nybFhKaXBRzCQBx80ZTJP0i4RjdtY1r2IfvzH20r1TI6VoLmKVfUAW
wwvlj7HSAutnd6kjmJbIoi1bncQMyhfWgq0lNfXqvYqs98oYhHrGchZo7q25Krrlv2uF/i4Vc4mr
WTw+wpobZ+OicJx/5VEdtToiEx6YwxWOanL4FS2GimxoXB8a9k/7nat0u0/rBvAENh9k/4yAhMl5
S+vM/Y2SAMYqj8Kfy9hEq+YfG5aKgJPS0XpAsPIEV42GWCSNKpRU2/5Of78XDQffKdN6wdH+PbXB
jlqIlz9K619rMJAA/ZAQN57XUBGAY1DMGLOIgXjv1MctLyOZ9TtNaEakHiPXsQ2PUTPsYI0af4oc
ZTEmz9kO1lnA6nOrUZI4mydkqnMkJQ+Hc2o+/liYDdgmY6Ms4z387d0d23JwFhvAL8zRfwqr5ClN
AxFQWCIwmtSStvF2EIiri4yPv5iGjV86yumgNXZVeySy20fG2VdQJafNP9kF9gNsXpy3+xomnTD2
IxVMbFiN2RsMhQL/5aVHd/a45Zdqf0L6vIHt9lpFvYAuebEw8+Z64VydojGq6YBOjsaE8DQ3kH9H
VFYu7mOSOxagIqnABULGdDravgamtqT/iav3IB6ev7XrGUnG9ZmTBYCbMzKmvwpTJeVYObMwRG6F
7aafwNonzb/tGAGwuCa3xv6CYPJc+OLXQ+9uwXm78kBStIQ9/a2Ky5EOikpoxc3oE5Va9Orqiu9d
EiQK3XymDjjU9ZY+hQL5xPE9Z93vpPnuulolInjmUxtqv1GwsqHiN5dWz70Zh8rpGYn/0dW2CjWO
q2BOz+MCa12S5z0d8hVC3Nr/Iasu4a52zMOWAwx6U4CeaM80LZ1scOKiZQNFCK3/SfmuA1zy800F
XU96KYXDrCRaQtYkUIEAtzrLF3KVMvLx5WirmPMZEL1WPXODUW0RjHgiOOiG6IKHigvSWUA9UiOI
ZP/N40D2qK62Ao0tQj3Qai3qc+4HCbhzd0SkrK+pRybsVWiQNxurmXdmhOBts0L5WRI54MAzK9Bh
GrlRIX+ohaMc9C5WfcwH34Vtx8dIT8cwF5AKMQL8MExJyKSzuTpm0kPGRkUVuEtWe/7zfDGziUux
TO4BisRcTyfm2WN4YOu24vP6axPDVWGOz3bLgwvMN6vHdXpe57ce9eEm9IiAHelnlB7HrniLKzZj
ux5AdlcIbWswmgyBVFq68Z6c6gXrD4P2IXkqfim59T214/D3vN0n94ci+Yhfj/2q59halkyZ4sy8
LVLqYJ4yCPHlplYTJQGfvcut7GP6h/NWKmABb5KEGo+HZSo7OABo47rVFoSKrlWSgD0XIV0YfZRW
hPMXuJS95xpujcYWCnO/1vJRyvjK4GzUIrtkY3guIA0saukQDxSGTCJMncITBUFMwAXmD19luwTS
BoAs7fTC43LDCu5RrJ6yCnH2gj6jApfinfauNvP1c09TPYPQlGX4u5+1jCiqbW+FSRYXBoKzIybH
9fPcUU78W06Z4gtkakwAw+WvLJP7Mu4ZHnEIwU6DrvNX6rgnoZIrDbNHXenHe/dRvVKkF1xf67c0
i12ss3cDpKnl66P4WVCay5oR44pGAcZebfZUvtQn3RveZgXtVKXsU3A9xc9TFnLhj5KMXh+kYFsp
NVX+zYpYGn/L+up5T3H3wwauRQEkyPSfc8hr41cCM/4X4RvIbUzocWqjHnjfBOObrBkvmvBoLktw
r233VGTY6vx9DbtKOCCmZHCVasBlXZIuQCmPActCWsS37BDGKOnd8VCoTc7VPqPiPflWyoklFMqE
/nqr3y1CtCsqvCD8NCz9j8weAGlgjQV2tg3abtaXWnX+9GZejiOx8zVvM6wONw1l5Vi8OEJxxMzK
mvVPfjsIUuH+dcBTO3AUa+UjxENLn/i/m3m1qT6E6kJ6OZpnbQ9iKR5kNokBIA9yfdtIuTCnBoXB
bhD3Baes1iczqlCldfoAWW7VNIwqiLsbysOW4AGW1d99dK3S6B5Y9zvNzb16uxM1yBvqQI+5n/KC
hvmhhknC60s8FFziCyK9kBXLbCcwsdE28c418MT9QyxKbWOo85ZtniyWejQxjpt1Q4y4h1awe85H
pjWKeb2QolHVUmZwGB+cFCjTjg8hBQVr1E0ihpOb0eHCSy6a6pWrHqZ4ibMnfXIyaV391u+NXIWF
6oxtg0dMFME2KpaOCYpxWvwmm2cYV7POy185qIDHJ6UiSbLUyU4vVHQ11fIjkV/D2zVbqW8J3NBT
o5BvpypohviBpLFk5Un/OWCTzY9PMtgfAzI6CxpJXWATtuxYtSAPI44ZOIZGmpXqjTNLo78Auia1
b2MNPlc+gJCzIcHKvT+eAfA4MVjyN+fEXvpc2/oxVPPVhX83LV2ZycfxVU4UjWZIKUEKUVwmpWV1
RyQEZF0+wfEtM6s9O+1THiiBxtCm02aQqFYiwBJc2vTsNoc8+EXTcKDdXxT+6Upzp4H60SFTGJRd
iPK5QMOKCHWfr1ZxkMwH1BpDLKynW0HdvehbHFolXZ0rZhLVs1yzUsjWece4z3GMPkfMOoZGtEZO
I8dNEs5ClUdcoyvs8t8g7Eip+doL0lo7IrENFTJUQErdEcxp7X3+QRTC0lNWxT9al9wCsOSfKIKW
U5FkpS1Nfn0hz4avi2p/H68BsLVZQJRLs9Uq8i4YAgF1IQR+HFIQNwK3ltuBQpcTw9rdkflZw8RA
XTiUbetKdI3IamXDOkvv92GW/I7eblCemcRK6iu7tKeTK3iL0uP0QbqcTixN629X5gyMSlv2OUEp
bs3lhljnWtOHX6nDDcZJ57xBxB8aeqBcMAYHd4SVTIlwz5SI3jZboGdj3MPww3WcjTCe4VG37K9O
6L5LdEkDfBr+GhqG3vNo6Rdr+fy5zFhlXw9A7fecrbeb6lJ70wzoM+TQf9GmDaRjRzAo7gk4ja77
VUg2JAM0jY6x/ApBIIDlSE20hLC1fldl71zvNaGtmt/e4Y430kUVfA2WgrWqI7kEVdrTrT+4SOi+
aKDF3ghfSP25h17afYWY5kp/kBtkQa9QRFKZzIVTFrIh5B3jdfg9P7BH+IIYes3n/ZphRTfFC1hW
wH6Eqv5u4xibezl2mp4VEzzh0eEwgu4Mw0dTm6kV3MvZsEfMsMxOhipHTMV+cmH+R9LM9KZz9Ah7
WU61nOQ3225OE2XQENoO3afZvauApUGdgaXNGrbPuGyAOqV2GwcKkiCdAdbQMXwLaUp1v+6qYsY5
AA8w36r2XQm5RIWSu9HH/8L4q6CyU+5aeZpSo6JeKX9Y9039xXaoLtwjUGqDaUCRpVLhTwXzfK4c
lIb/+inluhhKoUnIaZoHGi6O2jTjOzNM16nwK+L/Nw73d403D5MLeDXXMlLvAskiPNWjgwqThD1d
W2tH3IIV0ZtZkjOhuqqiDbcqwaHvEb8QGIkxqAol4vvLWB3KO51esFF2XSROkCTauSM1GpkAk0lq
NTamuGFMe53xJh5/77bTR2PWwfqZPPFUL768gVR6BdlG01e7UKid0EkwEvKnGPB+SUlNsZdJvg8T
qP8uV8J5egcSxnsZ3UI7BAPnMHVx4uDqQut3XQoZZWM1x4fLfX8NXoXa4PNJG4XPa+JUtnlExFpd
g9AF+u+wQBU+RvD7jzuT3r5FI6JJEM7LCYCE1Qx5kq7ndKsv158nBTbDa7D+SkSoe7qtAl784eyv
jhmSA1gQwvFeFGh7okjVkZ0PE9/5r4ETxWbbn/XG4Cmnwg9hduiZWvZ45w3bBSUJuJnoPHJ+azjz
JHnk6YFW9awdQbNGDp7McTB2smFJsSn1Ojcg5PqZJqJCupypHCVTIMk7v2mR7pUIhHRdo+ih3asg
gn26KEbcjTQnI52FwOoG9FmRtj50AYUnJCU0uPX2IIiXO3n4KHaYnL/YMqego21KfYQ76sTcVlwF
f4YO4K0MZA4W91suCif8Gwur20ghfu55DQgclt8bWheJB12SQ1TcgNZfxb43754Zu7m7t227QqgH
BbW6VJ3gzOHmNVLfQCoBQXTrDiQ7DHybKFF6DERpUkz0RZRljuM4iuHMo2240klNkkSjc41HtoQG
Y7DDEQaHhe5+1O6n1OuyQ/xakSt2aqlw5yx9jjbYpCP+OuUSXmoJE8KGcJiQfI/uOcSAk1CRmLV1
XvnC8cRizpKJpZ+N/gTx7CwEhNrPPecKyij6H9rAjAE9nFebz0xZcWDqvBO6KHGDaSJ3zuegZsbQ
uJMUTI4P2ueskNlrYctg0K+CTsMyMoTJR85Bnqm2JCsk6IcFqRO1aIqFPK3NXMj912TnqWQ7+eAF
PxSF4LD48a83+9xsvlMl41UCjysmn5vN71DAPcorjguN6j6UhduY+FjJ1AspNWHx4AAWPovi9hNz
DxQkT6G8/duMqmSmTh3ZNYJ/DY4UIidjVUKARNxiB0dGgX+FHaqtXh7nH8bYHP8lJOXbLNEFKTQf
NAQj9ZbZEdV/D8T2yQdUg39VpiGoohWefj2RRoNwop4cW1EJ5jHbX+0YfrYxts39GhjvsRUtNbjh
T15Czr4f9m8ohtGtYEOISYXoNuS62oQyird+dbNEaohmy1JqJLAjnYpv++IhNTKRd/ZBGeB4ZSD3
OTsKlHKmf+/3NtRGP4iEqLxp98Url0cxibDd9bfq8A7Sl1Oo4F+5Eie4tbNafWFNXBHMB0JZlhZx
JXmIK5RKRux3TERtL9KercCqtpavKSLpCDdDqTqELQW6t042P8HK2kYC0KEFlntakHQBVsV+HVWw
QACXw8LYAvVM4Quy1ItJdgOsNtd1nv+4mZSeIV4iLSFN4y8qmltv3a4TZCf+Eg/yyqGgTNOFAUG6
3Xoy+csKYCJRZKRD6r/YprGCL+cOkIzwFxkD04KAKwKKd8ML5LBO5PJT7MRmte2l1+OSnfZCv8X0
CchNzL04WLACvbRi/rwa6lJWhMz1468EWe6Iwv0ndI+cUswYupcFhwcamE7dIhJ3cM/ZMzVXEqoW
Qbu9th4JEvAJ4LyRi3b7jtKWE39FY4iJfRoHckva3tt+U1QTJDgKfmifjyN4XmQ9DcqLYFnnbEE5
2FNlBa27WbeGTjLAImcN//OT0pEqkNdUEMBMfyHqyOo/uEBtXmCcDjneBbVJK/QuDCII1bAbuL2O
WSdCL61VmP6h0W8NySwIr4HBw3P2yaPNAqNZQZvB2QUF+FA7+LVrP6/Bs7wVr1zDqnFsAR/NKnCy
elEX/d61F4lGjQ/h0Nw5VsP/Y6FZOtT30/QtZ9EVs7IwYqJq4KMaSW+xbSFBRgYg6KnBiQaihPas
iWJ6NTDnXJC6zTfQts7x8UD8LRRPdijYIu6HL7nYCuLHon8nDWrkSQ0pHBlMhMjREjbhNkiZzihH
+4ArYV3xFRtw8owEJY3Huu5r2CBGJjb/Dd74tQdjDh38s+zDCExWK2mq05puSepzWnSZquSSiRdr
echb0WaLZc1zX+EIymavyfvHSYkVBoq4YYXjPnHk5Gc1fyPTK8uWBmO94kqSJhPFpuUTzoNuVv6w
kJat498dzOOl3WJlHzOqOt7c+EqRjpFg59AdplDfDHm6sj+MbCx3YkdzZ4MtsAQF8nyZuJ+MW4Kt
BOQr80PqBzr55jkG/DPrQYSSH/sG83trKHG3SzGNJSXVUcYivcItsDMTuBmCcoZ6/Bh/7V1OleaO
bVNAlbh25f2e8JCu6jJLoTCmt41try55Xv+DUifHEQtBWN2lJksk69/DAiReDNr13p5hzERiWEvy
7YvKSK5Qk2SmsAp/KhE8pXhdQ4c71ax7hkE/iPZgR+sKBYeclQ3EkaJ81b2Gt054F/1LOXnESyxv
NPXYBsPCMeP/X/bMJr7NjV0Gion3PZmwuYVMtOw149ZQ86S06B+iHvMUbQ/1TNc2y5FDcfn+qR4m
2cI3ltLr/HlW1u7rjJq15Xvf7UogJCU6kbJN0eV7Sp+i6t8D9MquNEl4g1dfbyVqD4oBOeaxA6Bi
4OnGVIZf6ngVDCAndZBbq9tsYo5Pfl/bQHEDRRsluAbQ0jb8mN/HHQzfg2QMTTxDQTPI5mO4hU9k
Bl2G7fknbvPThuUkIZc9CrrgIBntGh8k47a8pgkZN6spLcU+pz0niTiseUJHhjDbeQ2iIJRdZMjF
Kp+STDF+UlFODQFzJpH5GoLoqFQSp6w3P8cmZzENyKUPNhlRrSAEb0ebXAb+Q2JB6mVnoP8KhHD6
AIylqeDMXaGF2YYaFWQ8VeyALtCHjxujFLAi2mjNSSAK7ui2qgvnETOt4LhMqTQS5iLsYtuqq6Me
LqVLoMBZtDIaV7csuMoDZE3L+sRBD9KmWvz4thoe+XNTz9GoBPc1TXrUmUXNVTE1NQ65NNMY4/3E
Z7p8rYf7UaD0VKADLXCHB5QniM7f0IBitINFzGkl27B/zZI4UV/CTPCQkgIpXScI5RVQPI8cbVAg
4uRrGfK4WvwbTGH3xFbypMeBzDRc6qHOf4tuRI+pPxui/IuQfEvvjpqN7JIHnW0FQz9MoCBNjHbD
Q2iYwYjzb0YcjA2xQQ1Lut+nfda8iT/Nh/a2dQrKgi6P9NQa/2UftToMxYEjFt7S9XaovHOXzpeX
PoePxW0bJ/fc1Q3BKgTZcmOXpgiDAndEDlQH9XDLTJAPylzbfcC+/rBIkvGxSF1DBUHAKWI81mJd
l6D5K3oVybFyDJJ96WXhXV1fqH7vlY7VxLxCDVQlaV/oihv1GudUo6zdHWIs5kh8F5oGxW/PiJmp
8zutf0QLXaatblLfX3Rk/3bmL/eNbyjXlvvMIbh9B+tXQtSJLq6q4kTPx/iUItNSe/iLwJ5NgvWB
XL2Xfm45rw5wplrf7c9nSqxv1jEAw35fPlBH1BLEX2gQ6RE2JTDKW3FUjfaCTmcWBiltlELtP7x1
v4MeUyBTnzt7yR/JuSchrnyVCuv3HsIkPMMnrei+AvMS1Dfm0CbWLnEqhEwAk+UOz/efoxuB+NBA
l+dOp24h/4LrSlnTEdKxdSITJHcX7fY8BEB1eyses3QCLBkkkVHCnGEXBsoJCYMG8564Y+dJ9kZg
ugTJCOF4jxLBGtfnvwYaH6nezT1UxaFnytID2nmYwFHNpnXwjARFgY251joPwF6iadI+3MxGQY/d
whoJ+02GjQ/jBv2jhpmFzNQ/ciyBiSQUYDTeMO+xcrTmoGzGjI2wILlm3RTx6JQLgY2M+hesbRlu
3QSrA/YlD/pxfNxYOLDTBe2cjmB24h1R5gOf2RlGd1VEnpcWJpEiFpJnTJxzGj3RYpAyZ1kfXA0B
Qfpf/5H6wCzAyQMMiSDze4bi79L/SNL+XmSwDkOG85+4qj2YF1SD3Ko2d9QDQkRc7l/tNvX3IPKf
N2EayWn/tbMnHOYxXbTRJXqz6em08YFCSntFJg/nPlWAv82bQa92JPzsicuVBTEnO7IATGwcCJ5E
H0yXscYy0EU+N+F/W+qi928DixME9Zjj7CgPmzaczmb46khERxHxCKOsAikqelSvd28aD4G9UtM9
4TOnHqpawcy3e5VbfOA2eL1OCOofXxB3ZCzo80YZ6HTZYpboFfwf9jrIUNsWw8OSWLqCaUuLRvnB
38NBpImfiTEUmDuNsf8cmUtrUGSefgu/9kt1W/JuA7MDq7jGrhlFfYDe/n5ZPlQgcBWvbAL/Vy+i
SAnaiTrZJTUD8Ca/aJCXzTUvJ5iPVxI3frgO1/pnmcyy6e3NYHMcXqGnLK9CnaAMHb/9xMsVT0Xv
XBLDByc6JOvI1NGpq1pthjbMhooeyZmnowgotCz3dS4Kl9iy/zmX8cLv9RMdZHVDpGQ74/rQ6kDw
sgObLH0HzhI/D0b1kZkBKqMFwhUYP9I0ooI4oLkNH7ROetmB63NxSkXASCu5OT2d2DjelZdxPB8l
JZddqYtnLv/f4J8y4/QL76GSsvzQTxLeSRJpHcypgkOqwUKD/NCTjzv83KpYWS6kEvTgD1zwKUab
k7StlAs1pMBMiz5vDWGHpy9kRNrI9sPpWMmiXrhMqxbOn9MWNY/M+hTkZZXNOm+m+yJOwsgr/SG9
vobOIuXgS1C1Y3Ettlnc+HA/zfaKMUQvAgEKz06r3sYo5sShHhMADGMXESIjdTIXgILTPd2LHsw+
VgqEE0qVd9tyRtpJMrUBzeoEotPsD0biWOAoXvf0w4uTzdKZpsqZn1F1ZVi79reVhTtLMGJFj8qu
RU8k04cmvLKnB9xkQlpT0hQMdsIWhaSM4eplm12bi7VotFwFn5+v9aj6+uKL7cga91/PaaD2vuOy
0qV0s7Btp8K64hfKnzJhvJgf1yi3Cm3fTPxzwhqztg4GSD85JYBrBoPL2EM1P0kWNupzFpeUX3OZ
rjSEh4a6DRVttusUMzM2UPl1yO/QM4u5Hh6vWhfQ5sTwmeamIGYqi8Xd3PMD0GErsZ3TXiCp5Env
we9RoaGYRANXQXzKwRiW1iQ+tmR8VytsizrJbYkQu4xdOqLIHd4GO29fSU+7med8MLxk/Cqp/W4/
NaCwZKj+7Nnczj6THulZLdr51ZQmjGUV+f5+NiJAafLgl/DQCXQWKJGpH4/B2USpoSl/9GWadnUo
9tAonWTq5t7w1xArLWG+QOmr4Nng+DgMSfB6uiwolSezn2D0BUSL/IwVOW0uJ6EdLTje+NfZdoch
nYRbrXnab/IG+W5PtbBz93SC2oJcn8a7sQhrot/I+PgP72ZwlFkFBb2URpwvj8uVl6dTRTPkOTi0
0Hb941iwdhim5NSdxTPMedApiiI+7dDxpRB+xQcECY4ju30DdpO2UBYMnyeG0yWicJe5Ruy6CL8D
98OxcnR012gGVjOIkkADnhzdEAgiZAscSNgxvU+g/SEZZfQBcR/IVUSKFK7NRhjAUWw0yfwV7OHh
4LrXnMBNKDQ95R+MQRqEFF4sExFXq7Bxh9+YyeY+xH76v4PE7u6fPDB7G3LhLyffJkkoHYLTn3UL
/8ueRaaZ4fdRP/6q8PBHgQipQkH0Mo2QNfskkhznZs/Z121IUKHq8WDNSE5kMFcGZmxwVpeHpPWB
W0ZcD0+C9+OHxLvTvpkiSApZ6T2M5nbXEwC9f1KX13vj3rD7waXfn5F0ULlE+vXNwTlI/94fPyBk
+ctn+8RdyvAOheNttRZWkEKuZ3hW5ByiSxOrCe4B7Bvb66fOt5KtzYFxoNXE4SAI8ReaJAmcgpgk
DgpdoRFo9lJ6kmkEWK2hrbMNqC7Aqa94uvpXemO6gtm2ncdsHEJoySv0DFr5pVBqjWBimo04YM/6
MnjsDDILo2MwzVaMLISFh3rNnZZvmGsrLGd/PaiicU4WYYv3e11eSNDkdXUQaZmim270kc59c+E3
UTP7fX+A1Zh67fFSIxoi7+JEGh6U4xXjY2tq1HL9X4Gi9QDncXJjaeb/1VhZZhvHRAiv2LQAdiLf
XV+9Df89nQ7mlVMgie239PtzCbW36dt1PN7U59Oas4edlju3JIAm+nbRI7CT2BXCJNX7+JJS5Yis
vWhyRmT51HFzbeSIjUEPSjViS/74Wke8jwZffj+OuMIkOjaCrCiCVCBhuOAbO3UVHrFCkMFmnPqc
GxwVG/BfjH3R2GKJbgPhmK5UIHXXJnnUEBJ75kNfv6wCCcKW08rhYEUV61tj8/eH6MhNuOzzNXg2
u7K6ouWuf9nnmXdoflJ70sKC/Lig/i75ZviHfarWvwAwv5FqToZtMleqEawo2C4aL5Wh7yiCGB83
kF1XBgj0qZI0Vwli+RDsFXMTK11d+ys8mootY2X1vz8q7HJtkfpzLUv98R6rwL8Bk0QpSoBqiGA/
KqqSZBcQ+siM3BzzlaRkYbI1Z8+yi50ognWy8ylqmE+OoRKwd/KovZJOuUwJaOCh/sQa4L8XEm+f
P9GH8gtNfsYBYx/ZHLWzfkLsOvAMgpR166OS6c7gocPwmUFuCa0WxiKqAh9wGF8tMOzLx7mtdk1L
Pe4nIGiWWt3GtiYyXN8QPOWf5bMuBmIRrEtV1M+yl72HdbVe6j+8da5YKY/phZd8lzWnD+KhHW3N
sCmT7aGD3NGgIrxoJrPz2ksAk0DsmPUEQc5rR+HklRyCBELyciPMhUJK8LJnlRn4UiUF3qMVWAYe
9+MFXlDSPF/emMUmyjYN5Tn3k9tEBeHO20n/S7I65xZDUxGKTej+KfBnxSJUnxDmr+0SkuopJCcq
kLZknOpKmoUepS8UkUrxhRJcgEWcjKX0LxUj1DTU2ExXiwB1JzbP8Q0Oat66L7l0xaKYAMs5a8Ij
l/U/I2EXufhPB18BtEVErDtPRq9soeoqoE1EwpiyE20+/YStGCn73Wgdl4ktYaJnWTL7Uwg3pwgc
ySmnNnkeHrqi6MCdJvm+oXqrDw8P6EmG+N4XOY9mGCJXYawwR1wonjb8lvmRYSmo3kziO06PEWej
1vtQvvM+MGKmgHrMkpRGfH7kkJd/0H20dWnNaSLLfIegR7D6sf8E/f7CpJXSP1NAvgf4qSn+ufNS
zOaw+exqwbjxCBRxmaAHTInBrElZ1ORJAfNFWoX748bviS4PEpEQLLjNEAxVzBhh7daICjdm/V/G
UluAMUrlppsxh0IkCsrG+xgpph/fFHniEAbEop+J0ZBSy9b2kk3UuaiKFDM7FSvjAARS/8o7fnhB
tWKxM1Y2AldkMhY5u+N4voaa4+GreUP79wVNep1yFxVe9pQ2ij+QPKdOB3xnfBuiVhX5cT812iIS
+S88ay+ERzC/Q/R8BfNsZlYsoWKvmxGoRwhrNdks23gnAzUZMN/FWv0e83SMRcc+88D6JfYpcBZf
4anUtFRWLL2f3ME4TK90tHqAcfmqr3CtESaK/cjWpvR59sj8hNTQze7Hq3FQeIt5fynV0IhruTRj
LZ6JWyYyI9OCbGhJBuF35fkEVM66z4Hx4rTtLiu+gp7p4BdR+LYuMcD7A0NQPGrLJRoEIyPGWKin
pzJzSBV/8r4DlPPNPe3YuaedAdw5y3pdax8QcU6U3cFCdQmzeklmsDRDIyIdai5OIzafOoCjLbgX
y5Z96rHttkVr69GPU3jzjowPQddNSqsHuA/es9b72M4eilil1Qx+I2h7bQ0vY90TNol6PHtBqrFP
TxPPablwG9Ec6LLUJC37KJll4Dn2DFw15fcfSUF/0wu/0hK6zf4dxpSez2w1puosMZYvb7tybIYZ
lfkgyjFvdPfcvGadcCLUtcGjheirnY1r+1ylTQfq4kAXEV9sjjAkqO72Y5GrKP77tysfsKMvnBNF
p/8Ju2zw49WNqMDjGQZtTpkWT46ZW2OTX+4X0rDf3FfYJcFlLGkjNJbYnzVJfQW1zlqTRduWV3s2
B/PG3cB3nToc2XBVlps/4G/V7wC8htYhG8SJ4xSJSQHP0L8FJRxt7tbBcyoaMH8PsRSUpi0iGnWe
vmv4tKkzrRX8Rmpjb8MIyg1T3eh+KZhwf4OOAs3oLclQr3Hzxci+KdoeU3FlGggPUPAj8FAoJA0i
tFhH5XP8uSSpDo+eWkdjQfqqcGLaXsWaMGeRiir4eTWBvDCR+VUDNHOd9vEbD8NjCSFfRPUgHl+7
L/py5KCN9wxnfBdOmjaOyW99lQ6KMqx+q9/txvxw85KA6+AsffN9M9yeuubDu/FJsmTJMoBMdZ51
Jzsz0BoddJqjxB8V7gz0ckC0yUX9mEQF/8wNLANHKGMZGvJxmbO5nfNAzIEq3FjWgPIMaXk54fsf
6a+CX2HQjzcD7Y+uTRYFVvBgzs//xMEF5SiStooyZjzH4BEw6hQdSP4Mw2fMpntLSFMAZB0YbpNQ
aPKdb/MKXr9yxf4mrhl143oW0SFX0q2fJs8sVYKgAbF4GeRAM51/WJZ1WewsqSxyuK2r9OBBLMDN
NbvWxfIJ14MGDnEYeGF9DedPiius6xIXu/e439ZkVqx8aePzia2NLouc8vrWBwHi+Q1kJPqEle/E
ZxQ3Rl/0z9nWuOJHI3v+mTO0/MK2IJogIs5TxznLZ7tHJTAfV3XASFvuHt2IAO34pekvGH3lhXcY
LYWPjnFUJiYtP9+jxQk/JvkmyvBBOrTaA5VqkYf8gcX61AX4/QPkK5R/ecjEpo61jtZV2ejXR6mZ
iSTrvJ14g11KbGO+fTM5bDky7cLeRPQYs9Pb+Hk4g03XHYFZMNV/Y1qN6oiwGPFL8q5XsWpHrm9n
ZR23kUBzvFsF7ShiimH6/FWqIR7zkK1wnAVzAURvO+ansg+wYafofKtPUMiw2Ssf+eZ63gIgofpo
90Ki/Y6aiUVPrbwMZAxC8t3FNY58DZ0KhLindW0bV+X3TQh9NHl1Uu7OHNRUGwva6fA2+pq1LdSd
+CZhbVJptgFE7eNXyiaewe9C/0+QGA/0XkVbsSlYBDj0oQtSKWp7NfqeigemwZETzPVH1YmVZ1ZX
YId2gpwat6+hyaiLBShdXRETldX8mMxNCmX1ztNOS3VPAWcY6a2THs+MgFVG0uAYU2eFtvkPfmSb
4Rqdfg4zJIWZKQWQT51c12cnCEUnuft68wt7xepPQFqENm+illOpUCaRrQ104rAX6gzmNrj/GXoO
zfUlAiLTS7m89GltJDOmNKgXMyouYlzGrBIVbX8Aq+nWz1sx2ZPL8uNu/53kxVoIi9g68xm100X3
hEiV9EtO7d/yTgfWo9iVEeuA1JA0YMSYPurh67WURiMbA5by+LU7u1EGkVWwFAPGKrm6hRelZL0s
/EBR0qiDb3O0K2cjMHFCVU+FUQe13najD5yfJ0wJxrMgm/Ipc9Nq52JRUIEY/uaWK21S5WpPahCH
X3d8ivD3jF884n9tfSOrLSinmlhDbhBxNTKaNdBhBI1JiI+zKPPF8fYQQR/UZyABvZFTvEyC0/Wo
OTyssifM37123ItnyVocr2urkWR1OEEiE7N1CzCIcf32E6F9RJZRXUbPXoCutRyxwCM86iVt7Xrn
NzUKPw06f5mKHl9UV4e0OUl+fH7sACm0lYF3ricOFMw0kBHeSj88l1wQvF++jd1YrfHjcLkg7EI1
LLc6WglV/5K6wZ0j9n9Xtop9CWLQD97SfV9nBhFJ8q2YclCNAyH2Iynrn31afg7+xL+5q1XEypkf
jA3VZL4w1Zh7xmcUTQ8A9GoJuM+QCq1ked/dsHCV4dB6WPq4XwnjI3MC8xL8Z/6QEk6UQPf2mdBN
vS8mAFNJTttpY7eXEepl6Vq9aqWLLJneepvGC8UqNTEKfOvnPFg20jfyvq4U94rn+a5ILOAzYJqw
mMt3Nq1JfUDty9tJD6t8DcbnNgjMBDsjzIC2qsHSXJFeDVeetiFwYlr0UxsM6eQVB0SfE1YZsdag
G65V23+XrUij38sRz0QWkNY6YVWCw6pWpz6fJPU8i7TVbPCVsUQ/Q0qMcw5LfO/4EwdVkjIXQEUQ
1IzBCw/qPqbou49fsA2+fpYhFa19knA+iMjuO8iIwuzZ5SIxzFw4DdUXQxd0nRFksjYMKj2U7mQl
7ZeMRx5LIqUTi54JhKs2lI7gtBh4IPAkBokZbQbTDdW7B0iNYsnx15l3dEOproaDULSVYVPq4gEY
wdx0nRKg4StybgADiYf/mDznmSiW9wrzcEEAzpX9IxksvHqAMgYzMfb/0RWS8WLLe4vc1TQATRox
NU7Xa70jnFOpXmFjpTpx6vQctRbbkrTM53vfBq9gbzeL0tJy2VXHaqjjeHKJ147fXNz6RdHxTmyP
MQDkC2lYJHUxY4zGJStDXXLBd/7nRGeEit2zwOqOg5qVav9JnKfQUqIPmVAWYXjFN8d+LCfcNi+q
smAjTB1JOQkddEfDixJ6Ko1mmRW9m6NZso4If5jPnprIr0268HvZ4FgXgGx/fzIgfzuTetWlEScR
9tfVBtcRrkc0H3my8ZoDSd3wdPy+Cet79anby/V1TfSK9Mx9qC41Dk05CalnSSYHhZaX2dF6N3+L
5PA2HJqS/Gw35dMq+LikTyOAlT5FZ+sZSGFRvnRsOhrY74rJEsa3Z0rsXbZvERy2oWbu5I1J+/kx
dkP3+0twoMvBQp47ktcNhQ8YOSyednvTzwad6t2gUsolRTSJztKIPjI8/FjwzQ2ENRQndC4SjBQs
oEga14vUmjE4hezc8D5lwTbAMpKE41UObWrcfSC59ywMMPAE07CNEvCLu5g2EhyGgUPx0trD68bG
xkINP4i6Z/gEOQc1sSsOeRpkNPbJIcbNCbsjof/zfG7eAQ3GRkT5QzeIwphKDDEsZQ4844iJ6hvt
rJlULm+KG7nLSD3MW533kNy0aRnZNa9pU4sn9ulbANm0IwUPYrKnGiAVAcTLkkDi2xv3not6wheq
LR/Sg8AP2SlSzkJLzpuFNi0NSteo0yLjeMLKcOIiqng1YSacSD706KBECTT7ehYGI5kVoNX5k6Mf
RubjvoRe0lIyGYIRwIaBPazxFfaMv9qatIcf0kUSTBmlxl4PWC5KoLZAfTljYtNjOGVTRIghhaB0
grKesvHxx6upcnuC/HzWbJhOIJ41+mnFhlZG13QMxeL4cGcuJ1Zl7mREZSjaX1G/R2+HTTrHUIwX
wfyMtYhacgz0niSl0SqgfJ93Yh53ewZeIgATOvC2KyVLx9wMuB5LZLqECR1AoIvCqeIFIYH22hiY
Zw3EZFV+ocCgmw4QQVrnvyrtaYZv3wWYRvcrtMu5zkqQH+A360BiZBtKqXFXdJeDuVwBUxll6GmO
LhEb/UTaWiRT+MawRRZlKTkE2+Gx2CD38WuT7p6XKmDFdNCxCeHwU0LTbQgidZZDXzcEsn7B0swC
Xi6o1uWVo/2pF+kf85Xob9x2Xq54G9nhBA7nKvRNSYtuyht1k6gfUerGsEMjgFubU8zyXHSSCl1O
JmdkvziYYT0qpTKHZqbWVad2K43gN67s8FXYp+REEtxokAjE7medJaA92T6IF7gVR2zhzRF2Tn44
1RBr1eDmOcEBguFy+SYZ+8522oWzZpQx6bSmm7uIlos9BHbu072WWJ3KqJKmbXdXXVTiTwwwV2On
S8r4hhwsfkQ02QpxqF1ohNG0zD88kCMTziOsnlf0hEC5jwp5oOR29DQleOlUqKLLLQbcCoKyF3Y+
5ZLuPPAo2fwhC5tKL/zSrmjo7zwLhUOCfp1jFZPMtc+xlHCpoTf0p9Zel1QkVsqgLf8WsupdJMAH
xy1PG40rywN8xexKussQ2b/K3jW3WaNxz3GbuPWhp2+m8jLM96JUrHdPKGkeCt/CAun0r64fwsQj
bdwEIUmADYo7kPNGm5/PbPBIrAOPJy5eVbLC9W9ZlkrsO4X7c9N6b0yTXu367/mLoKJB9BgWmX6g
Xw1s1SeVS0YEz48P9rhcJgff/58ZXNaiMCp4etd77Nff+651zaC8mmGnv/0BGiANwnOgkmpfVMfQ
wx1bfNjJ2dXVwBPm1SQPVaSJx2pF963gv6DI+7tOHdq3YRZf0wKLmVgfkXfEQcs0FZEtzzlHcbYK
6+j+HJFg3tC+dNBJa2T4X4aEbARvqnqBUi/6LsrqxjQJxV3CKUh1/5ZsGmBCqhwp7qkb9XdM4XJi
aZiClHpElBbqSqALC4VMEn8CeVElUgcSqcRNvSuZQ71rk9qdqsHGZUQ7rzxauwn4RPcG46K/r8T5
Fzn0XKce6tmhqFxN7qTud9+fxCmKImORbeK8L/gkshdAtFmaNuisCzR/NdO/V8QvMiHMUiq0Qf/P
wBnNhktl5A1uCaNJAmCjprcmM2lfI1elkpr2Cv7k3Gr0QRhm16NYsXAyfzQpr8KRDwiJQo+ITyZb
7nuwr1XCOGVI0RVIniPTY1Y/sgNJ6AJ10E+AtjgV+DI6QlelO9kEmKvX3FjKJcl0mTcrNEmCpw0x
lESPsmOM2X1hX0K+BjSlIF/mEkzjoL3/OF9WkOpHOv0v/GD4hg8/imMNWuXn1+jpw9ArQXqak2vw
EXOULTro478/y8L5bRcAKkppJrAl73LRLUe1JKqq3ieDW3+ytvA9jUsgoAcCOfFwfdEdtNWpD2Q6
AiG/eJhyJU2K/5Cw6K4PJOORnxr8Phq0WkWJFede91ctiEwTgDQTNWVViItQVDhMWUFerO1Slx11
1oIBm1oXSZKaijDF/WwhUhHtVo65rOQoFsVFyNpBpyLmi/eZfv4ij2Z1UONrzWoCUWDFMn7raTG6
4RTEALrIECk70+5daAZ3boEFcHH4UUX3ZwNwi77lR8bUTA5GuzgKTXjGZ0BxdtWPyUpiBqeDObIp
/E/Cuf33zrdzykN71gbB6Gkdw/Y+KLFnuKxvVc9qb6mPmDgdQBg76IKKSy4RAhW7Wg0O4NbvRada
l/e2xhaLRzmcrAe3491khnCFGwYY3j7GBcAs7jWYFCzYHBi5XuiPp8AFVGiKlzkXr2ku8SVHUHB7
BZZrr3Skfy9HsYMgNIcs1kkk1Yy9lYbZRyoaUDAr3mKcymL8GHLyzJ/ibxpgN1xjvOdGBMzknw50
lWgoU4wbXSoFW1GUoQX7NfUztw7FTnz71mq2Usdg5JfF6Kui7QRidkH842lY1L1RmTDl/oNerjZs
ujKj3JLruBfvFSE8+UcMAyUTxXoTDeDpye2fj2f5RAh8CKAR9icooqsVv+M7c4QaMr/zm8M39glF
tx787GWeOag89CKH1dnWXT0VnJPXGG6expLy/HenYltJxEXe7opJCrTV41gpZaY5m/qv8LtRuNrc
F5/ZUjZnj1YNjotjKA7oqtI9aKsEHOjKdGruJ7N+KU2N023iK+Rte9ky4VbSejWs825jqmKld6vr
wDjqHt0hiJiqkF+sOW1yhJOAFyrrsailAaeUo62H9wcqjYf0JMJ+pgS2kBwS3mWgGychYDXc2uok
oadQbLEICrxu10EoyGHtFnzrXcZ+F/aI9/pYDiaDVhu2QUB099TtK5uwSu8JS93gUw69biFUne8l
EV2OBWkZ7YrrTZmNYS/yA2GRJvVDrU8oBomAaef35x7TKRsyz6O9mdoEXqVPLW7bdncIiHrAcwu6
SGOWP4jM/Fm+CC6kY2L+yh18Xzor8XsHWPcBlNoeEFBzmGv3r7QwRnuGGtZiYH8PzjNg3ztSHnQZ
+xVM09BOnh3y99itlJf7wqaC9tD3/P/yXjG+P+TOcQrrDLbj1sn0J7bMMNOHCpjocbKVL2ZRb4oE
HfWVduaKxZ1XzbVt58OEquMdWE8GuhwZ22qY8YPTolHgcPghdnJClhW5bfOQxTrnaZSupGiOZdwW
IWgAXSEXgyWz0OHUN4h5G1zQq5xnu6wjiWsd2GZD9gXJ2xvp6EzIah1mIAUDjNVNlfCbFwYorUU0
v6i4dUPmQ3Jt0y+aB2ZOFcER/3+K1qETTKrnHJrdU2iO2wbRAtda5Y1ju9el1qN0ngKlCRmH2Edx
PpOGapN5IE1tXFSHkpyCynoHT6XeKDgLToJ8NGwGNDTiw+IBJoUT6htUuWZIgrAP416p5eagUP8R
plbzE7fC8XAGKZbJ0P0a7SrbVKezlCm14e9Q3Mulhpjepyc/3KEDKpCpfNzGgCzdU0fJJfSeYa+H
l7JXGGMinBaNz/9qDAdFSpqJ0A0DqjYr+NFhggyPIy+kwmA+X0uRnOuoIWnfAiqBgS7h8gbUM+SZ
hsuLujh31LzTMWzYJddQJFBd+7YvpnNTxs2hGhuPn5e1GzQOjq5wL2ijk6zzV8MPLPXQMfE9Ntz/
d+BlKT+B6R+aizvmMkmhNRtl7Vuo1d8iCglWTxRFUAJV4L69MdjyRpqSIFHQs6htIWd3lr97Thus
LTujS7yayBjQ75b6M4sdJAYn21gFk2unMOs3MOmnUCjNHDSqmbACrq1P9/3K5mvh34byaFgQuvjD
pwQ0COw5KkjeFi6ZkVYuYdMV0X6EF9oTdJIdDYLi/dd5w1M7LummDSekM3x24ElsU+3BhrG+QCIE
vB1oEyE68x6FP6SGkprAHaSW1mntiUS7184vUhr7AMGDfAgFtwIynr8lImWcdJEhMPOsFeM6mY4P
bWk/9/Umyapv1QM+twRXUrPEjwdTqh0Y0//SKXy2+uJdkgNOLAp//RPY7RfeX0BfqnG1uKLAo+rb
JE9YXlo9yj3BB5Bsv9b8KuZ9/HKxdPvZmgmEABaM2evexhfWjBQKmEHbEg2Lw3sP9EedmHBNFaj1
Minl1W+RDImvyHVOXidAshOvf8ryKLsjsHjaLNRFUTIFNK5M0PbysWXsBwaQc6K2sClVyawETQ8s
8tec1Q9GIgxhaobnG6oHmH0rUs/HAM9VOMspbBeu/VplTJV8OHRYck/J2svrI5kYtxeL59OalCDq
g2pVx416NDLHzXS280erneoIoFDhh0tOGh581VwBz+iu8hT/kYXb8wIP3g6EEvWqCNC6IqqiGAHZ
xc/xEZZUHETC49Pv50AQ8O444MYGuYY7YCFdFKbnlPWtshTTWJd134zLLIma/x9qB4vsRpnj9oxH
SMsWfOHDmoa1UGKh9Nd+GZwOpwRYA3fjCwIzN/7fGV1nuie1Kb9+bK+sAHhgz97hOdYVp0MaO636
fp3x5dWiLdVxpHU/2yt8L65eEbfHZ4f1UhOrqPAS+Mq84VumRt4Nta3pvkDAf1itK7Zy+0LjkHVh
CdTuEleqwfymPij5R35Uj4qzkT9HoTIOLUgLcsByScQJDkazPVPHOlvvw8wIB0qceBcBDHYsce0T
owo37XIiHiQK2sLOvVsu/mmn/Rvbxge0vjmBrvYOON6Fp8eF/oitVpdxNFAYy9sC7dC6SlytN9SQ
YS1FCqGQYQ9L8ZxJ8eb9fOOx03PtTSDWYjMKebOv2v07pW1UgwLoqgzQlm46SLPaYxkhQGEEkNWW
tqB4aC5ux8Y18Hslj5/BAQJTNbO9KZ4x057AVQKy54+S8s6rmBsSCdIS4eDbtnJDe69ohZljk27u
/qZd1qTDiyroIGgwZr0ZPlY5pJWfeg5SEIsEmmmgnY88wZ5qb+guPeMqji4DC4dUPhTSte3CD2NW
SC3zxcF7YOuqjJGgggLMK7UojiIzyRciKeAMqw5XJ0wWLyCCUthBB2KpiZearkteK36btm5txK5X
ebOl5vBkeu8f0eEfNFmYTcjhdiWDi3rpXh6zis+Vx8R0ihDrGdKJZkgojRW7KNtyzq0/5W6SNxre
XOBcGioGLStyyluQBQPpzWC5WkhDVaN78Xx7S3JXjW1RchsLyTqO+cZ8PxFRsYhJ84WIotcx7zjB
FUoYpTyELBuBHtJpWhkJNn2Geobm85YY80hNFBAv+diWsABT/7fj/hFDhDg5cREImSnf2dAArDuh
l4Jau0ypSbc3RdNRyDkobgLFUkMSz2OVyOwMQDNbxWROu04hgOWYAcTVZPuR8V8T8OAT3hAwkgHO
Nr5IrAJ++6mYdGSiutLql850G1BDS02uFJOmwuYq+fOPu8RPPvylNV54RlQ/MCWkpM35uVGi1goQ
IKICTY5olEl2EZv9Z0uv6a3HURd9iT2UJf4TCKCB2t0Uku6Jqb38a/NWyE8fswWz3hYXUa0j9MCO
F/k9Z7bFO/iTR4SLzmMcr+C8u8vDtaVNxEovBI1Rv/IrvsOSPTIg1THVcm6dAJ/LtfXrCCE5sFZb
z/gvsE9Bz8BoOPbEKms/OuE6jjSG5hVgflxDpioJJ5VriFGwgBh7slmPcpd+rukp5o/bfX2Pt7z5
bnw7/vm40IYvZR4/47o05DmIBGhhmLpfBDNSHPd69Gd7jx6KZiZ9Icg//vkO6xW1L4oAY6FaOFiY
hx7fVpnQ8Es+FlZaKDrGOq6kiGthRH0FiucnUBCdbrzX95CMpDi6UwSLXoISHVE35NN6MLf6shyo
C+Cb5wZUxlOH4fFmE5tG3Gqb7IwY34Xoa93x52bq8lwYxFC0rvJk1x8bFoBV59ExKgK62zFZB704
i0M9CPeLbzTELuLmqP/IIRi0VkktUY/RPOm1h6P0ld48p2i+WU+W9OXk+TWsistzgBGJ4sjq5ia5
O+tEDcmrCbECtGlbp3JmZIlavyalOVF72XasAYiVOZpWW5vj04eR7zMDdY4yDEXcwfECSoT9xKnE
H4JnyCEeF7XmKVFvRLs0ffaX4LfYJDuzqIpleyZ7TaaJrFi/tXCsi9Sh/ttYTgDsEQ+OHpP7Ntb+
2HFy15VZSADY+bGoLN8uRpejtzXj09pdVJJd95DufyNqtGDiA80UnKbALNAuh3qKOICX5hIhWAEN
RubgjIquCLKnm2ao2asdfavUf84sSnP8P5g7cEi4C2GMXu0+c6faEbSUo4wCcPy6nN++8yjPYkr1
erPg7ucHdwgKnNoEVHQKuIjtakpwkpny30DDuXHMaEXzgo5KFNeUJeMeW96QGq/xhdhU/IIJsKg2
lyW6RNdx3iwGIeq1PNEvqOdLpH0WxWFhfE2mFfw0v4iJAvi8SRxlhDdhPkaRkQvZCn09PPGecw9P
4Ag0KydM54I2QHDkvqElDCjhzXGubj/YewqfsFQH+T4IDXDXABtWduqbJ6N93AAtxU9xCIj031vK
2Cnem6CcjxJ77RJ843h7UWXiUahjI8vcNI7+yDu6yUkcZLw8KS451yTK/Vip76dKwMuN7PGdpWzL
NiB75YHPosIDAImZjTHiLyjkHLTlTr5eZytQZ1hydNSECo+VevkzPekpou1NIqX0wwfraLs9bRB1
SsY/6zpmmJmokKneONX4N8xZObhf73Lorro2ZnuNlwky+ZkdaWreF4LsBTIBmYtLlJ95P4R1h5cn
aeKpu4Oc1tyYjKC0fNV4w8i3JMzW1RKAIK83bnNFXBonzgeGkTBTGGahWVDhh+XpNyfnDvH2LM5O
d1wjD/WNWnvqjl1dm/IzlffAB37K6V1wGW0fdWeAGVOTSkBKkpSsCDNn9NJOFrahg/ljae7whcyS
icblLCmB5YGCNsbv9F1P+xhwXnZLT/nJsIskR9ivSDrcSxns5LPB7iByQ/kWYrz2X+HymkDK5+OB
Y3SIGcfROnPODxgc5as/WJ2Jo7Kzm+sdrTR+9gS5fQpYLpRMPNRbq+aWRFAb+fXj9HMJjEeVghiH
+rLz2AatmZmXAJt0HUwB48w4AjyCSfmZZPoZvrkbRnifuoqMBHZbMFBMHqg6Hd5UmNqOv4Al9tMU
7cjoKMMmV1lPbJPNpA3Rrbqx++U2bZr+xrxIJN4NZnJECnN+mDOIrbT1zo5iIzZxW5BCLwSey1Vj
J8Jvr6hRj/soAL/3b1oD0PUFjPJXiewa9Dz/pgvvN36cKn9kqbL4ZCZBolEkA686Hk6xmqzueNXo
kY/Zz2Z71XupwpBLL3W5AGCdpH6v5yxVuhSjd7EKfuuISr00tzGUtjqWiKJ/TKAV8NELSkZx0PF8
sXfLRBYLmBFHYLs5dNsK9FyCYtdwzr9/3/vwfPQpdLaB1U5M68kI13hVRYnTyibzI06Ys+u5xioY
tcVC6imw9IVccXS0nSBLlqZhdNCzQitsepB6k87yYBrTOzUYsEJ5381I2dqTONft+Ejqsd8sMyOb
WkCV2gdEPCFIltiTZAHrKxOb1l6Ny7Ca3+jiPiDH8SGvSXUCE2DCBSbZYtBThjkbQ4ZJPPWpNuOS
fluLobQhQlg33J4Q0AAXmitN/GKs3PVrpPH6qREU+g24E8oJ3zOJiivUJkzCXvhLDrIY6Ph8Z0nq
J3QzAaBszJLbfmZnISPukPxlu9NtGVdZ9KCShHhRto5FP/MEixpC7Ulx5Yb2QDkZOLkNOcjlgi5s
R1NZBefJDaBLoXtL1oNWZnjgYbr6pN/pJ9MxQy9MLLrIyfffiwtrPh6g2Jj1njug8eyssSzqPQCn
500Gnrdv1YJtuzK00RTkCs/rNJf0JqGvlIYmz/Ysw1PQqpZef3R1cN2qjGBVH7bTEEjMfCCGc7ek
39uWiPYxgzcpAdmFc8W0CeWKxU/SxcRxaT+LUfMk+/A9HjZKJDC66gBeSM74wsBwIV45lrF5td5U
WDBV4hvi861ogkuxDAYbJYXukYKpUuwJYD79Y35vLWQhwldKY9VSTUN0SEHfn7u3DRO4Aj0NrAEj
7VzzIyGLDB1mt+D6RehKvDWtFMtI6KcwjUe+YdGGcKzvzUn5b2LScyEyHx0bPGxBzQEV8n93Tghu
fVsLWXo0NzjO0TP7oZgVsIfhygPQbh0Uzl5Ltp6NpidT5pzg7PUzKA0B1Wh1lXncY1ATbMTFpibz
ARih5XMN1NzvZk0ezb59kHXa5Iju+1kswlPTxSqiHw7vOXyV0cG6mRiZc0nY5YavtUFJKOxIq17h
qlpiZE+7TUaDGC5TDE17cEo5fFw2/xegb+nt2BDDphj9/JO0eyb0TAYV50Cgh6kB7eJfxEzGeji4
1u3K6TjpaO6Cy99KneKtLJNF+MZ95sX6KZ8H5gMFGTcu3/RA5f3y6zHsOVAsjeDe1bF3upwU6GHm
EIuzCogg2JUitD0VZjUsfKWKeAD/oQ1+6+m91A115l8DhE3CUS+fZ0nkLdDHNl5q2I4lVJIP7122
erFbwGnP6YuUdOGg1WirCe5HLK4friq/FxgLZ7m5y18eZus2QSub8nKNTjXlXRiRqwHetbvIUEx2
qrauKIvsWNtBtM2fXZSjub/Z8BDARGawi1z2wDLwPRO6zsLrdKWlxzJ7BH9xC7GHg5cwkFUiv2X6
+JlRlgfzNhRHx/I7uOcLDGGEv1lHp35f8e5CBWB+Oh9Gi6APRtWgXVN4Mlxgagp7fl3nryTE994E
MlykebOC+Idt9FGQW2EAs7ulg4x7nkBj7mlmtXhlNwngUWp2yhN/DGnadb0Xjb1+EJNNAJTL72Lb
HkoPEK/4G+qhSyS1FKIc2dhc+O5wfK9OoZXfbR/XuuYh6UV9k5HlTZAjhEPBn2+iA+2CHlW7kg/p
r4fhxb7BCXhQ32Ny3kTpYGRHSxGFuL6LjWbRuQXNZTkr6hwj9RNCXhSMlHU5LHqO1mqX6emHvlTS
1haaFV821ewwuwHATESHGBR6YCijnKTkev05D8nHWNAKkUoEn3p/IW8f52HZxF0e7N4F3WWoCNcv
C+ibWsxVSn3a3nhYMtXQKg9+S1f4rFYth4T/C46Y5D2Wc0BAuxO5tSQMh7YSPlVqcxGkbuR0LiLE
JvIgJOXlZCRC2vf2CIoiUSW5ki1O3qijNSHwbqL+ddsM05N+pEAPo3OPi/gRBrDOZB+w1VQ2gx+/
Kx78KjTc1DPtujUS2R8xd6FgJee8Z2GnuWrdR8SVzEX+H9PHVL+5ogLmfhCLsd2USZJIoGILJu5m
8dqZUsrXwqvi1IKSy4rs66wbjYrCpw2f5slSyAOJUyFGXzF4GfUPEPKhrTYhLyMmjF605R/u20DE
vFDSKsh1Yy1BP7MvVe2TWSXrhz0hU9sK4LDOZM+i+yVW9O+fjXCBNDccyjRq1aEeMXOSxFL7VGiS
EeRDH/SfR3wAjaBTSgWRI+ctekUsiIWRIgsml0jDbs4mN4v6nP+NZH7x7I/sMSuPhpItD2I58QYh
NdEEvgibmRd3sg+RRNAb3snY+QBXWsiDaRGpRCWiiNV+bSJKgpQw03JyNZFtW0hKbsyiEOyo+aSi
UmJLuu+pftvrYTmG1bvIN0rwd7BCrf0JcsZQIIV+XccekwHPORdL9vXiwuXuj/xwkk+6htaYmkCj
z5zeiiUk0P6Eys85wFBX1oVLjQhH4wNZmiWjzf0r89kxTO0+SXUoAFUKSpv6stIQ1BR5oLMoGxXS
O51TZIBotff2ekN1bP5+dPbVMg3w7O/gj67xV3MRxLQcRlzmp0aLMKeu7QavksT7/O5jFmH8D2Bd
VNd4MjoslyGNkPiqNTaGYf3tBT7VH+oXj7+1GnJcemyjJKFq4aJmyIw+BEu1Rrp1qDs9UT9J2JBK
zgX0RpBMfVy/J9RdyrXXwoYpsf4rmxfztXJRjU8IAiozlWBGP54gcI6C0Gse7iMSBxxELa3yq9At
C1xDYKLOaCZkIuPEDQR5OEa8HXQpfpcJKhMGqsH4C8hSHN9Jmip44F0wN4GqeqaMbBrCBDNDPKB4
dTX/0Lj6Q7gEujPz05mJzS+hqGBdRsQ6H91Yl7DVjNtO82EKs9AGpQr1ufHsQOawj/au7G5m1u+U
ukqTetet+SDoZUtLfOROiH1sG4OnUy1hBntOiarCapRpwFuxcUzFFBGcJ+1AmXO9K7ZVJUpLHJCw
x2VkQWjFf+OAkD5g1HmGBGY0aGZzIXRRVeFtISm5LmQ/l89iU/AXZBbACmX6H2zb8GpbEtrYz2EB
rtO46lM4gimJRWW6bEgAZEpZOCc9xLYhxucOv7Dfsdp3BrnRb1tzUzH98UROSKH/bLAWbDySL8PY
f7Lw7oz5TOAx7H8CojTvh4lmi7SPGGvLtCDH/xd7QnqQJEDbLxHpbONSabwKjjjmomuXi/oo2wEp
1C67E3swdGRMzsKClRfP/U8LzGn+jhCJdOOYrHFNlEAyrLWT6iscaaihG8z98i1QBp3poz0K1v1K
lbBcrfXz/Mexz1j++o3qQOu03rtKvp1H8eji70Z0nc7x4ydpwB+lI2hI11cr88c/+d0RlYDEm+Ej
AFYHI93tQofblhAcBW43XMSpCV0yKDAaQXXnoHomDPLahpMIzbFwKWAU7vUPj6xLx//WD73deAB1
lk26qsMxH1IIKa4/QAb1kIx+mYqnonY4NjrVWZPdEL4GV80UWCmxJCHKR+tsBtF5QlOVI2vEsxX4
Afrd02J9zD6IKx/UFbMrtvqZzXoYAenAdQU8Cdu//S2nuzNdX2MGp7H9OgeYVv5UT/LlcG7qs2P1
KVsyzkDrfMqy1TZfah+8d3WnU5xcxJuVCOE2fj9/vVTWj09ksVkgmnBJ0HwxIc+/iVd4GSn6pWJI
Mp49ELcAPcKWTIiSQuyC7Iadla6/rj7fjer1rXGBgacDNFMqzqz6Sletqt+pVmwnGGFQ0mwLo5Yn
OlBVEwYifQTtgXref4zYiY3q6V060N4gx1QK6TngR1S8Q/iIfUm+3tjB5R+4tFAM9zdBD8k5eudq
ytMmJ1SjTdB0GN4vcFCqXM9TY9tAIaoLDjA4JVciFRuKahLCXZuu5fdUm1U7a3tuzvi343ktfcvc
+RqmZ4oYQfo2B9BNMAgBfiDs5cMlsR9im21BwBqM35petuhn9Op7qM54rnNB/hpR3gd3JTiugP4z
hytGpZ6Z/h7L2m0c53uCxgCPBq5x4SNkrvj33IBiLIPedi8Q/dy31F8ky38lFwNPDYs0O0tdTPEp
79m4CsGXvre0XfV89ggqAicCPXVSl91GpadQ/stuT6icq8eK+nKN8fdvphPfzYhtnmNVC4f2F94q
0FmcfyqOO6fsooReCq3du3d2tcvPJF1Ua1XyiWvMm7Df4fWxmuiN3lMvjG4DjMuilXdLdXVpFLrO
US7i/p9MPhtbz01EI4CibMW6U3Edqg+RBwkBtF5YkRsS6bBF6PVIz876JyJuRhh1t5MyxVXIxkOM
ii6Yi99Bbo+SguL8bd+jOsRZWkCtIRL9KlPWmZcP7ce53WL2UzqjmSOvEfXGld/AV2YfvG+1UhAG
8m+WAoiJjV99mwqNwd7/7NlYRsuldjn/wbyjy3uhCrH6MQkao9xBrwFOcxMm35k1CZ7FKcK3eQkO
7Zn8MoPEuEfWW/cyX7RvfhcAoANDxyvkVUIG0FHy2v3iTljBr167RosJ6S1hzWqNxUHD/VAI0gBl
mueDJIZQfRN89zV39xv1iIHuOs5R8Bu7GqDkMn7XTO7Q4S6uhmR/PwjRuVbTjv0YDpRJwacLDyN6
KonkDRKVrMTqij7taILRIxDHhxwJH2NLzBgNg4IexeU/RtUyXcOPWl29y+y6+Nw3OSoxntF+Powz
HRTBmah1HbJxWS6WNmvPQlaYgSSRQUL5R0URbkPtvqplQzrjuRv8Q1XVmD1tuuVnk5SLQ4ikPRIm
FFhg41BMDV5BnYDpfWRLThm+gabcXNIJZ7AuXV1GMQTDmkbGoWoPXNr+ZiEJRu/wWiZ/9OxowpBz
RnMz3ULgYUslnbIrG/zY7tIxr2h/QTn+t18sGCnOG9UdQZ0qngkTuw/p+6Jr5O4ZPAdkudeiNybU
Z29mdq9VF4dDKoLrODqDJVSOfX4sEO0FhSWTYMc+5ce2J36IuUGqqXU6XdlPdfhrttH3kuFtJAAn
ykktujZ76U0j84klwcqywLIGyW1VHwKoSTutIIA6kMiILpeQDSm0qPsTEG+b1zisNeJBTKOObTv9
okDBUaAj67WJgQyrCJ8z5WB429FB77/Bca8p5PSlfyc3PD5IXkkjqk5H1wiRxlWA33xo0JNBcRs6
phfuZ2mNLE3CX9m1i6ROCCzAROYC/3tyOtyvB1HjNP/teb6Oe1b1AilnWRqNXhkUVDPBTYC7Dfza
qIMr+jnrOpCTH55/G96z7E7AzVYdxzb4TsJMLg7TVOonGB3xckAe6e0IPfyMPIekdpK7wEPyOmYy
Sw8jCVUB11hjJfwlS5QXMrMgVbPGlOZZjln3OCTSp5+WXulg0QMaBbEOrdkX6N/Oizh/uphR3yZb
zfrtRBNuZqGuDROY1RO+/DTegZAw/6d9tfkxW5vM1BL4iRPSiF2OmOowC8uIrDSLIwO7tGrn+G/z
aWh3NfAWwjl1d5RwyR5EVdYLy6g2muGON2PQXCXrYLxYppgLf2BJmrzvOmyn0R65W6GMJc2ru2f/
u6ptc79Ec42kh1BxD7jc7jSQ2TpklI/NNXG+mEsBijCzOujHFwt99fLsEuwliDjtiCNQZn+hFyvY
0d0IcYTxdGJTPMqjQjOKgTlrHKNojSTKG6N9FjC1H8RAHqIK7cSD+pHvCOJ/f4SQO5tQlsrUbtY4
+MjmzCqRxZXA+Eg/YsZhEtIGZaKHaYSB7JZjtXcweLb6WBAye/NXTI2pQKct8njIuGlWSw3e0SAU
JwjT1J89byhwF/6PYm7U0DVvgabCLWhAxbBanUJXZjyRdyIaF05058sgAIvHt8jTy4t8ikl2AzZU
wRBCil4pR4seGh25DcJruiR9kQTPKn7S2KfFb5bxeFCJlAALr//HybWsJpAshV0LiWyBGgzQnTez
DlHeA7B6YyH+G642Bh0gFmUfbMmKHbp7NaU/tcTyivt7+rkBt0kRk6twwFscTQALdsAbu/QaHbdF
rxuwY59LwBrb1f4CxzCWU3FmNHslIpaNUvmnYdkwCLyv5/3mdUTaWSsOA+pANWqwJ6rLTvD/dLzl
JZ21FjNJAy1f8G0Oc2qj/3T9ESY77CsYhyV0PXNBcoJgO4Y+fPMYRPW4EEr4qhHCrotjEkdTd7v2
MeC8oNV3jagPDF6msk3w24/xcUHGOnovPJVYUWkes/MoQKf+9hFjG4O9zjTjtH1NWOgIDBo7tD54
w4C24N3iz4iT3i/KTHyU0KhI2c3+NzjPlUrNEzVr0f946VFVa3G+IVwX3Ra5tRoQVL+B3C7LIUcK
GE1CamCTVWLdpe+148mdYxN9tgRRyQio6p/epZ1mGLzd2kX3zjjWsHG5em1f0TrUL7xuEcxeyO+s
LhoYEDP1lEx8SBbV0KJTRKUJPLvTDjMBOALQovW5vNB/J6YrUL8McWeP4JV9A8ssEtrt+F0L2NVj
DSuIxkv7nfj6N0MoFgUYZwX2pEalUx4ZK+0CLe0A4GjQA5bA+2twiwwiZ4/x9gWuOYXcNM9y1B4C
NWTae18I5TCTeX4aMNDhQummegHzxVd9yaePOX+PcQY/9p28VlIPg9bX8K+4ieOHWAOKTKuncRl3
OpLXAE0eXh8gsk1si5l8CrXSp3sc8qINw6jdPC8msJhGM9xYBNPMRsGAVZtDJzBU+mzstTpr7D0Z
Jq8e0vTWYTXQ0jYQjrQzN0zKk8DpsWXzYHg7h6DZ/H9a+1I9A8ymYcNWSQq8Lypx+HL+QfwWH/Gv
Y9Tx2sCIKPG0DgEBtAw/y0ALXFxHCLJ67Bj5astM1kVjgTSg+/qk212YiPzh4AcV7RWlTZGuhfGJ
9Y7pyF+BEY6Riww29RnWJX23836lwMKZmLoylsRThVxhGWfv++PmoerKQxo0e9iNPO2VafQN45EF
lZaHkp8zwEeLxAnRfF5rLjtOEijfKgBhtPYM82yIubtyRQ1pirEg1CNRjME4mAbxhi73T8BsoaPX
UqNuDjzxMnpF30vLsTAjULMmn4xwwPHs3eEDlkZQcUq244i+k1DIiRz9soZ480dBkSofQiD3Mx1z
kWu/t1W8WM8npMkuJi86hXwTqfzk4O6izvz2Gi7FvVQwXH1v1pKMCkIHXhftMh7nU6n8mhcVUR05
ucOe9I1CPmxIYO+qtuYYXVR9ZA/VlY7CB5EiufiRQR68M5tPqB/cBf29smBGB2ksEteMg2JiCAex
U0RFWxmdIZfKw5dYnsczAyxvf88QoaP/bwnmgOuAn608s4sJfjeN2WxRsW067hHtXoJ3D8yZqop0
t3chQMWxM9xhA38mlHuI8ZEdg/G6xTPFJwg9uAZDo1SAdo/4C3Uh12TCbOPNibBmbkXspC02y3le
77PsmPJObC5nuoiZZKxytJkDtOSHivTgP1ysXNbNjQx+q8w9hH1sTJqHhzm/AEDrPkOPPobV+xq4
Dcpqyw6BTqUaymLSgsfDXi+TkWpndgjsGA91oC1Y+Nb/wXaDEOH1MZeldyGanK8UtOKa7NfNfdan
vdpCgtp4c5YF71oxuV3IJtPP3yhifRY4LyuhbVCyXSD2kaYc99CYLmsFqCdvxvbcmHcbL4vvYngP
0iDxvF5r/YLTuka4haW1SDlAlOP4wsZ6H1oKHHxL64KPew2q1bpi+UQdmF0Sso746cAI7GPGI1Xm
k5JR2v0vdRyhwwfSdDieC3DKH4UKkhmT1w7lFoIos8axp17P94b/yc7ph4dRC3w+iwLQAHhKN1Lh
kVu0k2WDees4K4RYWyY7vxKKkJ0/6Px9Ia7HIkBKnfFQi4bou5R1qjB01So3d5M8zY2gzy5Lk7y0
pk0c6y7c3bUd7j57oSUFMfJ1aYXmX2ohhnhvQ+RWMGjY7OTHHhys5CRjOTFhaYWcDbs0EmBDTclA
+vnjEdPs/AUGbqQw4tdA5obbHaTk+PqdJqdkFF4py5qFHnL58s/ZYtJcmWfNOW8rqKu7F9pTuZCq
6BWDThcEBCIw4FBx2xGiwoUptnYxki+PP1QuTvy81OQgRb0TrzTTJYnNSlwU+OkxE68YGttXp8eP
BFUzAm3fHRLzcypC0gWgapihWpVI+PNw/fOiNT8hXWYRkFil/7pUr1J2gcC4/GUfuPw3LuKsa7cb
yFCAXevWSjUTY8CndTkkafIQMeDfqD0r/gmhhbQEWF0LosbBuXfPXNcPsxY+VlL8CMVFibyFbjBw
HWOUTBsCE3QAnOjm+wJ6HysAE4oKP8dtw4S73mJyzGEV1ixG9cjwxks2CuYnBPKN6qcjCjXc4nDe
nuw9tH8otk+rWPgpsrmOjrHngyosKp8vV7q+mxLVe7WJkGLgYb/0A+x6IR5HnhWa9lrSZhmv+PRN
Qcku6vRhMtiOyKJxs9BdfYtWUvLxDQU7XBn/uFYkVXAUGn0AItVGdtxQD4wPy6mL+YvUtrPuiZb2
MkGpO8p0ZsGAmpVeVDMuCNxHQUM5ayHc+tY9fpDMAhydIkL7GMRoK44RNHiT+VgvkRHMyMrQQKXN
5iwhQHe9QgWcKEVJ1XMUa+21Pr5EodOwSEy491jJ/qqnCATjUuxnEzKJHcVL/z3f+uUSs6tpmySq
29WSKb/BeH4cvX0pP/SOVw6GQoYU6QTIP8UurlfFkP2C1o8Yh0IJp90bKWz9y7pdRAxeJhk6R5V7
Yki4v0pTK8frhIZfMkHUYuYoddtWP9kCIyWF2tjl7WN7j6DcRQ2gmaKPxXcIZjwenifwn/MjNzjp
lhMxrM3lM+7ngRSwLbmExvRsPCb+RkGDi2o9AH8IzpEhr8bZta3lkqGdh4yhe/V1ySTbLo4IgZ/f
mM02NBdjjJsHYp7C2YwW5/VP2vztPP0Y/yYrmxL2tXziikHKRe7wHcTla8EgnpSGrvxoMKsetXjz
eSVnE+5WT85BfNR8qzxze2PiW0PGpCL0E8i11HLhOPfwmJrfM7PeFvWbaK3soHU8U+xCeKgmg+TJ
xdiWfwdU2Uv/sJhOz9fF0T2Wz0Q27fzJlh8UWfJnhvhYTSXBQ4tKB9CNzyApHeBMIXeWqjyHQYN5
eio9ozvmWfKpgxf9xmqc9C00xLcaBaj/NOIwBqkTHHLp7v+62ipWvRv9+mliBxidQ2ZNy8P0laHr
icf4eLuhbEd9TD7VZomlSVx8k0Aw66DLCbuEg/OaGBuBEp5plKEAqSYIljp1STnJWNsY2NFsXk2s
Ts/nUtpB8s41pvdGXd7aLQgBAOnQQl8so6eBoQ8V4KXflIW5TXLJjtxgio0r4EixhBPwHMD8V6p2
s+DHmcTEyJsXZWXg4dQaHz35tQE4eL3smwCyc0Ifr6H5gFFPjChcSJPg2htE/TN9e4S8VU/EGFjj
4ZJ5B2kOrKqT2JzY7lYF9i68UskRsfwOrVbqmg0Ggsux+ja036Fxyg4pafTLk876EfyJqzBbctrs
L9YDBiC71Y/KXXAoAvXZj4mLiOw9CEgxoxKWyYE6jsP4XONv/z+LjNgF1QR3lSnmKUE2HoBaTxrO
JQfOppC12l/a/mPyUna77kud0HtbZU5eVt/+rIIisW+1ksQ9YPGNgKpgD8KcnwT8IU0/7A2PG59e
vIYY6TfokFvsQgHKyaPo65dm2TRUPy+LOD6/NcgaLcbpd9GIkNb7sptkHWUIV6d4mNkkvyYm0ItP
cN0XOCxif4t418AX2QJt9oMCBUVHA2I6gWKOcDutZ7oKwvf3yTLVyjRwnFb3af1KE5FfzGXou4VL
ioQLvrROYjhUpSLgbObE+tvJWaGNPRjDW/un0ot2IKHdo09572S3T/xR5vQTTJc6yLQ5NXoIxx8V
ZdoQUc6yQdYwNtyoci93kXSeyUQ+YVCsm3UIZcc9RQFIDCvbFJ5Z+Ap89Dlq9O1e/VmpHlOkem25
zZGCH5Aiyf1dVpFNJQbH+rZf4T149OUDbfCFFCTsDwla9dzIL7PGf0aJFYAkGp8QrjhJoauPjVkJ
+69W6b4mCDJmC0uKV/uWJxpLQElazwqNtTfNcjIpt7nj4eE953e2Ls+ZKYx8LtDysUc8vbMTZ/B1
IWHeit1lIj8m4TJ7CXWImCiw0n3VzrM17uw8yT1HWfgqjBItNJhEUJoBxdW8VZw8HjUXl5FpmKpn
D+AjMuDe4gFjwo1SPspDe10t7/N84oJFF2kenbEqn3Bdfzx339QbCEjpCAgcVB2dffL1WNNu3qXM
lqWo+rA+4QITK2eT41r/U9LaFTmSBrlkRBDs4diGO5YHXprsC5eJpkCvh48NtrzZTjpk8J0XzHFK
5UlwZyHEWl4cGOQJXyEMgIpRfhKvELzhgymd5jVWIX+j6d6PW59Sm91XWKT4i/i9AVITsRRUiGwz
/TQ71NbgWuRp067FXlQtCUDEMYedtB+X4PkbMcCIS1gOOppJhsssqj5WC3y7T7PlQZdPdw9uyOpX
tHhbEErtt1Y7MhT4h61SDSBBKlEwWmAHNQJNfzQ2yqPyPsJ4IJovfjPtoMNjz24yYVJeDGddq1ot
IBTfo+/y44blatlDSBTXVzY8j1qghKlBFE7tVKIJ5ZsHiM/9StyiknjbASV9qZlvgliLEoerOIRN
GGAs28R2qMMdaAVEmXWlepTgVzRpFCATouhj1Rk2yjp5E8O5fUK0YDvpD3ApKldHy/IbUhqc6eBv
v2rkCPl6+bLRQJCR5p12SArSPMpvcvoyqEEhorl1c5eLC2n8YCvcwQZIQPThlzoqIqU+WknJR2ZO
gWII8qUte8Lu8lksNFEC0+iDl0KUHXiDCUkP3wPlINxShBnNfkZoqIPX3UQssef/vkPqyCl1Bbo1
OLq5C55a/hlX3mLKmdab0UaTKHdcNXRhV3LA6UQaBesWe77xJU5L/4x+3+oQ6G5df7CATgUB4TBF
pxzr8123aWhZYtkl3/8LKPyYXjACWxRsP07KL1yVdt1A6BYPp9gPv5RmD69GzbmpfHDM7Y7mm+cq
fumMJFzX3/jO7WcLGzerPbiMMg35vobV9Gc8/ZbbJC3zPDwkr3Qc/r9U7o05cE1+yemrb3q72TID
VZhpXtzkNCIXFRZzMDvPBBKQ+D+vRxy6CYOe3KNkTfnmE0a2PQd7klZXENEEpRHlAszIxNKogEdY
mAHsWtrCP2CKIy/6yP0GBr14aNpIKQARA4mT/0ITrUV+zyW6ijC1DR+7vlQc0M4OxCrWu/qtY5aP
MbDqnbeRKVzmznl4+wPsiMHFayEllT0dgctwpBgUAaUeMQKz+Orac0jIjagKff+moLy0D1M8Der5
nBVbTk498Fkwx+45qyfN9TWymvGfYalr44bPN+zQJDZ/RSZTVALynIVejmPsZ35G7JrAVFyl7ZlC
maa2b32U/ObEqv9tZEkjHBXHVXSNkxRVGCaDuPZjWvJrGiyYDCIe1C0BdQrrs6wOdIgu5c2uIJWV
NypVxiAzsKDuxXL1VOMlhhYzvN/kbMXCOS6jZknA9LPHSmwPyaPrS1CMfrnxhnKaxVVhuNeifEyc
gKJj788emNpJ7KtwIqNX2t6LJTYO6aH3RgfIrme1gNGmU3XApCXAVzW+fbLkBvIZXtkgGt3s9+Bl
boSE3ianW3s0LoeWFOVUxfc/oMezrOwi3YTwm8+mmd9KcdpWwl7ic6kVFq1oTJV5AZau/kW1ZzVH
Vrx9q0PByQVQvTcB+3e/U3kHRFG+k51jYuPzAFyM3MEiZw31Tq4OKiTM4bBKLKYTytkW/6c9qMkH
Yz9zUP8Hm9nK/z6o7LZY2E0/VKQ5VyaRochFMvSpZMu/+6ZM6Xu71JvL/Jt0AtTTCMnG/4aRnVj6
K5tLGrGCpQ6LXFuKs2qeqbK6PmHKwFeRvDKHtE8n5RzzWFRGikWrTVyEATCPVhrNveeBNEI4nA7x
3P6BxYhCVmP5o1fuE0U3IW6EunNEucm4IMSqQUE9ssvkSiTCv88ONWe+DlsiEZbbzqNwtKw3BAw9
0VO8Vdpe0vMP4FIcDcsqa6oSQcGxrXNn8E+MxRX/JXZByf1Xb+Cdc4CPNvqrAbxarzIs0SE9L8NB
HpC0ygESAuRVIJyv74HmMh3Q0F/t2SRX3w+rUri4KpbLT7dLMbXXNnE4d5o1bP3eiNeOkwWErw/D
FBpf5XEYHDHCpkkwkPNeaWSmFBVYTekP4WE7JI0SDySvAgLDxQjSBqwntxu7Ey43LzfwLIMeGBMs
2/CR93gsdx4bf7wD7TH0WeJc6Bj9rIwtWJUqdcMT75U1I1qfmpZfWqu/0WYuwCTqWf6vGq4gmrRc
i4M8zH5yAmh0jnMt4Ba+xnYV+ju0lWc66uWIkPWPI35y10u6fYY+BZYZtTCvGJmexE4EmFKoJo/2
4XGDJgExP3W921/uRwDODuK/By970V87nz8vrkZ4YCaf7WK7OjPAGkp1upxUquJ8J8ap8JFJx0gy
C02Df2tVTvjABTSngj9uc876LGupkRx4NqJSEmIYt/1OKS/ytEeUcDyzCehGO5BrE9nssqZc+pX0
hue3z7p3N7qBR0hj4XmItwyLV3pHD3DrD4luihcFsoxlnunyhULjP1raIZLtdBVyk83SEDxVswXy
SJLNyux6scLeW2TIeiF0nsKf6d6UAZctl3pH2tdlRUAx6cAQ+XZohxk6zWGwdpmXhjZoMmHA02Kn
ql8SvnBOtT3VthRI9tFtmTgfpAgYkqmlLAAKfBFvLEp0h8xQ2ZliaLAafawCnV3qt1UsyjHMR5Rd
ZAUoGBr6KeV9Va5WECUDBBuGeaBKPFjKrsiRrmb3MuTDm578ZG2eUOFjffIi2NcAYlWdPv6qjvUs
iL/ZtKhnHBdggqwk0zOE9lkY28DigC2LDPesL1v1hEmmawk//sqrMFMeqR3iUEgJEb74AAQsfP7u
QlkGn4uv9178QxbJAXn5I0liZBEMxOrSBKzI9kYzYHoSJJqR8+j8zt84F7RQRk0HorAe6txjQ3SU
P4sh7n9kgZPoUUYWVOIq2LXH9j9NoX8snjHtXYuYo+lsr76TtPG75wrc5OfsZ6ifXofiso5ChZmj
Fo3lrtzcAiSAJzunr/WvZVuyvtPCJi13Eai6WaJL98ugcopHDa/AsuZ0+VXxZ5i1HoiFrN+nwJFI
4BwEHGA2/pRXoeazL3xtM8Vn3zJUN0lB0iwNkwPuZWFycVz6qkcLTzl5yq4vJiG31OpxTKr17PBT
PwXdc/EcQj0bANZPM2Eiq20rj9Uy+GfrmtXX50FFqDoyjlstHa9JF9dqm1kdqAaAPwRqUWRwWtvr
k6vNcSrWvUhD29UnygUZtDh9J1bj7F9gk/eaH+80I+QGxN5FgZwMXVD24c6GjhIfFLU06g0NGTXC
sL+wPONqfa8gtQN/Wi2wiFCJpOu0Sd+eSWPXR3IHFEWS9w6cTP2+XdxN7kHOdUas9ck+Tdy564x9
D6xVwYlhhtyZN8sQv3qouOA3bFExXSCRZHoiOwH2t/DftEvKbpZARiuYdNpRafm5l5bYPJuvI9q0
O33oCYaqtqtggqKYlUStOud1lK5lHt959YshnkhCI8s45OJrZP2sPcfAlgL/by8kTr0c+EAXlS3h
tmYJzv58fwIIjXFY0bZtKTftAudStWWzzxXcZwXS1qKcc6kzudiY6lwwR6zbM8wWSOVun42sHgWM
3Wzml+YnLZiIe2f0q9LEuNcyAWlWVb+Ie8ew0id5z0nLj+fFq60VZPbc+JWASmVk+iNPmPf2Txmz
m1IvFoDT0Y9JjXPl47nEDSs5I2zT6OlHAO3sIeRObysml/igf5GSlt2srMWsHPhfI8bIEi1pI25H
NBB8ylvln/2uXaFgxhY7ldn2pr6HEB5wrUqhNSANFvIEEdmmucZA2ZctVoQHgiATY8yu7H9VR4el
nWJPtSsmbzb7clGVNrz9+fG1hX4M8nFLwM8TxoPS+QjAh55X6xWJuKLBa/sgJxtny82RhRJEWQu8
MHoZFuh4pvDRJpErBZiZvZpaUUO44YumnYOMYJif59PlkSbZxQu2Xm1VxSay1fj4wo1dKHNXc6Kz
fpIBQ3cX0nLMTZjOLnaJA8tZBmh5fh0EjchCnsAiTgBtUIO8X5yvtHBDBIF76IikQdgdsCj5YdYP
HdZRb2Y4vf+Y0yv7s372yhBzdXIVonVzTcafdTN/KF25nHGlQzyHpUSXmYZGf6XyjB+FdXNN0RUM
B3GotvPFT6KETg48b9tTmMfO4DrBP6DD2P8PCOypYJZI7rnT2TnhDFXLqbbYun8ZMcz5Y98EIWrF
RRNnjmhcN+vrFwNPhkJPwMNRMcCBl1ENzOsQgauiDjAllByCJOlgl1ygjpRuKLsXwTs8Blr32+g9
cHgdhiWzr9q3SMuNJFL6G3XGwgEXnVGcjXSVCdLa2VY8D2B+OG1/3A+nBzwdwTirqkH7CMVRRvcU
MQIzd9i55SzpyKyY8DxfGoKZNE6mSomKG+fXmGEZFGhZgyRFEC7YiL0LzwZHzW5IaBF5qWCzAGse
FV6t/asgyz3droe3WES0vsZAWdj9YW2VPCuE+oqeJGoGNlA/HxKszGK+zH5SM9GKgN+d0E7ONI/g
qDAXWv0I8rx49JwyTLwKFT3tbPwvpXV2Ripd3VlR5iERS/wctwo1g7ERrLfXaxmAF5hMNHDIZzDE
ARV4XKsBzii7NcpmSUlxc57WmaK59LWE0HPqqbDaaHTEtMVyLM5Qdx1AxmmOhLPgCnrqep+DAVM+
lFjyhwHZMMV67Xop7GAKhimXEhkQScm7bm2sjP2gNMJ6Yz0mGH5EYuWvaUTM4nfhvNOH3cXIWasB
9K2UiWDGhZ4alN5MLrSISDVIJKo8LazuzKhQcD15JtxpERoWFZ0ra6JcoxYbHC+Ga394TFUWsIoC
CIwjKbZgY7HBV/ZhX0jXhQ9iLJLRSiaka0WC+ZoR/65237HXlrhEBF+L5Aoks/JU3yrOuQY6vVai
wOexw7hf8VVInTrY3zOa9MqtQsxK1Kkgmvyddl19XhRC0cmgeUGnhjv8sWYIBkcFupYzLlkJ1v8D
GpZIggdh4trYpjhpijRijtdw4MHPzSxH4UfLCkYto4569W00EWuoH6E4OpIuhLFLESRG5mXwDP8h
0xBw0c616M0xWX/RT+uY4NrYrnIqXmBNiBbkjpgQIxwTcwJbVS91j57nWpPcJbk11saVRzyBl1BB
IuF3nymdg2/l+iKjnADUvKrCv5GN5CKP/SOcHGIFFF+iGtiSWXeEZVMXL/AJdzhL/Vp6Q3ViV/aN
HPoypiQKJ+66AaG6uH/mqelmEPn5UvyLEGdxsIrPC6IBadJSTO2kvMQ6zycE3sjSSR/Jpa2cUJbP
P96voGXe1YZDvOEubCCmmMz3HtzLP4GCu+YnbZ0yNbCkLqDGMItr47LhqaOk1FPmCGAIOrGB3CI1
zi68DzkXD0PD3NfiXg8DSpcJJmCP+vnTlWrYgu1h0sI4YFowuRy4OlU3+4bOj4D2wewuEyl9aopA
fCHDUjEbAEBKB/HrSmRAGAORr3l4OqRQ2K4xpsGYgIDpkLk1Qf4QZkDkQxEfUtQTW5poxSZEtx5p
RX+vbPI4boO4Y5XnOQXqGymTd6cuAg3zMMYcr8EhT337gyEFVi9JqG/RgD3i0KOjSf06YoF48L77
s0HPuoM+AMzP41VCTZli592bRgdwH1HOZWQANxdncCIoXxyzM/i47t6h/DSJis0aK5Vx/skn8KXs
Vk8ITnwxFkcQZAw8hrU11/nKa22s3h+NnaiAEJFJt8B1/Y0KMMy9UxWnHLSB39xmUCJkZIojKB13
ThUQA0Jr6/Xyx1axNtHVZt609/vC4eiM+7Qc5OQx1pVsBlAgpkeD9LHJFGwwmJOcvU2zca8Pm7jk
KBBLTCpGZHU+l3P950H1QolNpxx3mzWUly4iAqyzL7JBxPI994q3QQBLcbXtFkAIT+grreljtuQU
q36Y4yceeW0U+G48CbbiJky1NKvN2633CFQPjCLDdE7jPgQ2d7j8pl0BvwGoWYSE213UEZ8CbIEf
97KhyHzHHWkQpyZVcu3c4poamwghBO285HHH4E6uK9nD90VX7UTPQ0BJnpUsoQU2fDUALCcv47lm
+kvB0Oi9jSjD0rstZ0QWySJzfB075sP3TY/j0ddTgSuF3L9rqgKy0B2BwQI/fhwZWfcoBdyA0DlK
cFjZ/IgWOxmIuHm39LNS7Stw5D2vwIfr3yONbZOe3rAsgydzHDDseIkiSG3x5oNTs9uha8PBmxaU
qtz4Chas4T4X6sRnIbo8yDkSMqFdk+pAT4/UnEx0sNOVeCWqT90MhfhbYWQ6L4hQCayx8ugK/lLV
qE+PW54L2RtFT/vZCvApPfdsyCmFMu11ZbruH/5vnrguH+3lPHuhfRC5HOAsfQZjxgRUPPNWfyDU
WZLOfCdi/EMP2Kr+WKhJpKEr+CEw60+DZ/+G/72NqaSo3gbohz29Y8K6Oek5Rq37wzQ0HD6QS9uP
G9q5bM/8lWtvBliiroQwaXnsoDlwQU3HZZ+bZQVx0h/EQrkcC1RUx1HSZtTqbtpazJ0jiv9v+tcg
LzbPdef8uOl7G1oL3sG9Rh/C/5Xt/kBxCSEYYq9rh9MCpbdUyX9JbfYyqkK5zs+GSl5KXZhbaK89
r9abdibLjrSzjyXt7s0mKBD+PjH1m7cyn1K1R+9F38E3J+lZM7SKG19wtASYtK+1jDUMzGxPI4br
WFbWTotOZFM8JRHCr73av3h7cSMGW4+CiM2xzRbi9rtV6wtkczr+pRtEXvFarGCI0fQi+3uKcuP4
NvtFsATI3yVbnqBQcEOaR9CmCikGumA3oVdMAtOITsy1bVMZPdJoPw1a4XDWxO+InkMjrhS40Wrk
vpclYUfODmSTbjToVOi+Q/ecVMiYrDMm+59s+xJIqEOXZusmN2pfJxO4oAXBj6r3RLMOsqtVjF5d
sRelKZC9wux1As5cOq3ZGxjA0NupSE6DUQjFET1KOYt4YHX62IykApvqBWqsTHProep7ZQfDDfu+
waKGM204g0QXsClGpyrtQT+F4W3T6e7UvEkaULbJn9efOy+puXxteTYhevPihhhRP2pFOQ9JTJtY
hZAeTPh1wLK0Y6RTVF+jocOmM5jg+GoZ8GCs5K5PlInmmObJgptiexFQPgJBArBYMCv5OQamayJF
EKasvI0IK8YJNUS9TarCc3nEfFPjKnxrtPE/Dtr+a0IWoWsi2P/cgOWMjlzHNtOAMNCkjfmfxwVK
QV8khgDqU1zIjK/0i+o1xxnA284sDPYj2kdqMnI3d9QcizbkqgRwGeF3pY17NLvlTe3GRHJ9Npe/
jGXchtw7JCxJDgddZs9YqyucOJa47C3qgAgN6qWURtLNtL707HELGXOeDt6SjJi6FLL/ghRkn8Cv
1CrSxmxeJg/vMvWE+SWTnEnOkjz7aXfPL1bbs/YnXo+7M9iN+crYzgDK//CKo8Yna7/EbUbHzaxE
LDZFRKXArq/QUr1zVIyAqFPOhuiNVUjpow2LMEQVS9nbIc6m7lNiX63O8XghC9vVTuAt+W0KzQ2m
jnlxEx0DVjJcKKFDqNX1L/9waQCqlAaIIx8M8OngaA/LIeoGLVNCk/ioM4as8/UG2qKpAT+laiMr
GKeFk9OiWxm4WlrthV/BGkpMK4BCubMPU0PiBorIAR27F5ValDk1HiyV3n2nXi8Wqhszd0V+SCXn
lC6EOL45TMInuDCt6iMucjt4U20giodc3bHbvHBaqQRb5AZmr12YTKC8AycjTCk3dsGnhYEenmzi
ilc+dMWOT0htD8nAR+KkMxBAMZ7LPAWU+yuAz+bZVYpeELx4OWoApJ+dIQvJTgg1Tp2aAMxRMYLP
94eTmhR3NY5Y5qizhQejc+IDYfxM3RxD1gIGwbA0clYZ021yuqPX1j4Hm5JmqTBQkOdiBGtaF/7m
AjeNKRZG/oYUDbjRHRCQROWQpfxMouwjdt0EnwpTdcyn/o9TNHOvetmSa2XtVqeovvq+oAHUcIxL
QAH19VsXiExSmpwvExLfxoA7jaIKq+WFCIA0yyJMQr9Hj1I/htUeaEp592fa/b36bgEdmOD0y2rf
buDX4TPk+6PDGWFJKXndwhQTp2u+YeAhOX6d6zsCSTEXkgN0Qb9Qikn48PT0JM6ABoMwgVldaR2m
zxMP2/ZXFQmF++8DeXeJiq+0haX1S/TXcOTKfURm76H8nPzVg37wHHhF2Pkl6hWhVtQJx+ZHK8LC
0vv/Az+ZwJk1WKZTjYzkgbS7BCCuvwVlVjWOeqwxxO0g1VWcmG99/3QOXCGylMrGaSceiaku+hvl
+uV2lieZ+cCfGLNQ8mNjAv/+deKBoxhEkeajld17+f+1P5vKmZ8xyxSRaxQztrVoXS//7W78WlIA
wYtyvDcEK2U72eDid4N25bCTRx3BpS8xO+S2phXIXcd/3mldFMVEH8w1FhsM5mgLP5eHMjHX6TWf
/cN0qYiBzR9kVa5e5TFj4FVrHullitwrFzeqI+dFn0uXZo6rNeEX6Wz6sOpeVxsvLS9NdfQ3tPEl
8YIbPJ+I/cIxxZ5fOjmD+Dm97JmDbei8CxlE2xHSC1Pm0xHfys9RxIiJOZ9XCLsRgyNQKtCDWYqn
a2bz3qWTK9Z4r0C1TS6/HZY5vysV51Z8LbY5hSLIXKtJ2VGvRju/xBeCnBgRj5ZfQK/NoPKOWeal
HUadqseySV1aXcJA3QaRD6PG5eh/C7c1JUTbdKwZFB6XlwO0jU8UJ+XQsheHYdqwE7qFdYrhza/x
CsW0t9Xks1i9uh5QI5nszmf7s4lcYxFz9sZYF/0mQdW+co2pMS+m/wIZZvSo7u6XOqQ3Qo7Rw9Ve
ExLDRlOJ8JpTgetHmisBQaIJ9eBkSTOtwGcpnPaUuKMEQo9E0tQ/mJLsEVh5HyKSPttRTwuAGBcL
1LJodex7VHTx6uv7oVNMV376vpDrdUIQ1/uT68lopgFB+ph8df6MQ6ONB+rHdXVA6ASuRUfjwaqg
VufI0MP1aKNE5kldqUGFGlMKBkszU2h+nzd7xaXt5juC1hrOCwhSWcl/BT0PcisZ7Kw32opg9SDQ
LnUwC9GdEb/NCw+GfKUxvngehFZ88hHcpnPUefgZKNdrxK60COfk0aX2Iqk4DFt3v4DXm5x0oPNq
bn8Gh2swDKdzJo5yTANH0vYjQNYmrfWFSQchqieYOdrFF5tUuhWARhZYEGqN3HBqQQ77Mrw5skWR
7wFFXajLW+nMMO5L5SDnuQqOgXyf/1DIn0UsxZm8h8HRLvPVxh+NkudxM7sBAGw0IhyTJf8QMUc3
EihITulzBMsJPxzHJw5x/dcxL/NM3bM4LK9QW2KCU/Oy8oQPHTxzy3loZgsfX9JX4dXlCM6mkKpp
OeQuIio2ck9UwT4ZGvG8GiMxitt/y8sWdUqYwkdd0fzRI4t7wDF8hjkg0IqERUGjvfU3WR4fTxBD
lLuuz0veRNFMlU0wEguYOC28S48XFRhrzD5SbdGBrW7a+XJFGYK53cuM5Zzx8Tn0R+zWfqVcf2BO
cgC+aRoSsYTH8NAEVwtRdXE5nqiYRBB3lgPrvPbeWDMF4FMjGNosg6+C/Dw/FKtDPPlZ8mWxtn22
KqafzrYcAWSt5Y7xM6CGqDF24wojiRoVDfl6HLNFvUnDreVa6N9iEBPTJaeNX5dSTiMzCMPLdThb
YkNA6qKGwP65Xq9wffxQkW4fqY+zvrF4+mTWPAK0+Z84G0ZKHKU9O1BNZ9eYVmEaaBN8FPZYHoA9
vxM1tbagBcMpjbFtqyahp2YudajjZaucvPR5IhtoE7v0ytDwekxHmor7Ez+utxmV4URD/+hH7/Dt
guq7xPaXaIMxfUZi/yz1fsSqEOUFeIThSncfGVsldwW6XJGOH5FFBJbyy8LLMq7gcnkIDWCkscdk
PKdcH3fgzGngVT6TPh/Q3PUTTWo5PcSZ09oyBl8wfcRa+cyArGlr0HeHyDHYKWka3Ah74s6rlRS6
B/+J0eAggyFV09xOYvNyJrA9Mbt2M8Ycs4R4TSgv0sS4v+wwfUJBOuSBeqFt0lIGnfjcTJmoHDgK
bHE0kDjq1AlAi99vEMgqbtLIY2JO7sJGEWjnObmf1whaz2iPthq5UxNTH/WVx/4VOmhpN4kAtF/6
fe09YyFZu6vv/YNRUw6TpH4CFPEwomxoAwt/R5sjqdHmTN2BGAQJfjNhZ6pnPZ1FPOgTCfhn8+20
YC6a02AHpIMAmZvLHcdY6ewoskW51AHYbRSx6B6XU0z2rMVb4DOIQeO5oFyRvAHHn07I4tGT4ygM
AftawbQkmUMi+jMbESnK/q00obdN0EVodPvbT9JI7wmIhb4jNzNzmVgyfPGR+X1j8vGGrzTshmuG
IGLBGJhdNdiwYRWRnCyPjSEenOYaDi2ZSeCWHwIldt0vDj2ODpHnyBuQlk1zZB7kYsONgWrkwFz3
BwzKH0heTTRMQ8MLID0hJyMrRyg+67gyQ/i9hEKFZa6hV2lYv0v91rg1/WAePeP5kP+DK9O4KgwQ
pd6J8eIEYjdfPH0+L1XLHbx7VstGZfqTDU1RurFqxPjZ60LV78jWse30CeX67pWZx43rd791gRmS
rbfCL9XKafTcX71QNaZEr66LDvA5GBmGN5QLnCs36NgkdbAfYxbIAEIMpCmHeTuqaKgpyx0gb7uT
A35ENrvujGzUNas4W9h9ylw1ndxx4UEznEWf67Mc5WZLlDiJNV6qRlQHE6MdEMK0GNzvUPBMCFfb
Fj6LAEaZAUfB2X+yD3NYW3uQDtFqzoi4CBmuY5rqnQPC0z3Eh35KeLwiZlPN/sXCWZT60zadRLVD
YeGJKi2zkCXJisKo6YaStJ8PMAfgpyg6ystc2oQouORUvsYanrET+M5ER6o4FwpDp0K9Hx0uax/P
7cuJhTWOeZioRprP0c//mYFugu3awrJYHYq1SUXY960b36saBIVqy9jilAQWv0/I22lhJInkYkbn
zA7+O6WDIpID5e1bUh7nAVS1aDxGGYcgcvUHj2+fm2u8DCA/niP0ZfH63mkMJ3q2aO/C7t1kmGXS
i1hD+eeVk/feLdJOHcJ161BoD2/5lKfKtRkPYRi4lVSAaqN6OU4qPlderGoWJpEh8dSgMq/oNJ1X
sdKFwZ03MecNBW7YBXqyDiQeoD1jukoPkeZyQf7uiyTagDvJK08f0Wumsht9LInlrQvqDNWeetqq
kyzOVWhQEoZyrXHqEKcZjMRclkY94u0AlPdN9632UDazVPo2dLPoI2+BckIfqLHDNm714S2W5Qcw
fE2mTzcvgruH6bkRRULXE58TWxT3AAngJj3TqoUc4W8Q8/k1O3UNzOtmL6YBPDIO2UgHLQdEGy/c
/F3j+gaoJ7NHHoSXMitRR24VTTkV2/mWuxvE9CASOWGKV49/0RCpd2Ds1viAbdHaCGFGBtAkN0Cg
N8zl/Ud6dlOYsaXdO4WrT/j41K37YkIpDAx126jHtxlv+sgHGVMXaSKUZwt6jbaA23/argCkUQwx
kH077QDVIjlGhgko0gh6Yzt7T6IMXL/s3EkfVSFYutEp0K5Ceggv3YKjTlVzNPcs3Xs5pdq4xRnL
43PMQQ5A0KQm0nL9KPBU0/YrSnIFqIT4cAfv6OtR4F5e8HEdqsOfCL9jZnIZWVIKb81qvWjIz/Am
6EBcM0cwQVnxYDE8+Qh72xpPfV9o8+w6cnaRetQQLDThfZ+EAQv6heuZFqIuaDVaKs5pvqsleaMZ
vDocAPrdj56a0UjkcUrsuZLNr7/6IZmcnR/cXL53PJatRrOdxXOka0p0SdNsYcJCt9dWXVo2+6Kv
bFULxYVXsyoEk4d4iRH9C6eqACGMznVEgDhTzPBAKC1aLpKOY5L/GFkPWBfWWOFPIyTdBzuPHy2m
UCN9xjdDuUXi6konB9q8TQlWdd6rxeWVBSM07ghpxs15S3q8rpso4uj3l/+hGd8xx++S44VSuLvM
l3w9miAD7XGH2iZa+hV7gRgVZxMMjHLQuMXF++tItnGP2jj3a+4omaBJMBt71tNPxTt4f/wMG1Ik
Smz5rpiHYudNYpqqr4bFOZj1BrqZJzooxAwrwJIrb4CgIUCoA9aAd9P8AX1snvy/8lNqDd+1lvp0
TZ5EfpMv/+ZVhioA7JM7CuqoAM5ZBN56lgWTeR+rIHXuxunoHKtcJ2qEkRLRDmJiYi8TSz5w6x1D
7LUHt27DI+rXzCq0DOBKcR1odGM7oBC2K8Q9dHlGPZUZQX+i9AJlzNzGy775LIQcBoT6ggnYfU30
8078G0Lm1nRgC3la/PfOzJKfIp5cjalJCZSr0H65vbmnT/YGB4Hno6FexqUzxfGFuiHNdMJlPdyi
6x+SRk+1H/ixKm7GfQsvL0QE7/8D5akhaTeX4LqhpgQ1liOK06nPFaArSFfuLR5Q8f6Dn8J7x7Kd
KBGMMbclG0tXmwBvNIextD2EYxsPxDNf33rTrCnJV8BZ+ON0B1Ee5JAF5CE7t7wmA3ZuUn5BQtyS
nRDw/44s/E8rnRRzxosFnJ/072nsnP/SOxkzKoxzBBqoVz9mR+oYgp8JhZQYXDxA8YKEoqj9LvVk
TUekxWeW72MRE7Q1c/ulMRFiHPHO9iSiBG8d0/KN+jvCt4SRvHjdrTTZgThRciCdqbPZ7xTj+JD2
9l2sZ8x306xCxOb7CPKA1FOSpgAxLurauWZDjkbxa0be25zmTorzPeLVUqEb0vxN4jxmeeBhHi44
9JgyhHkFWW6FOEJssMmmHFDTtOh9ATSZ1IDBzrTLVzr43tKa5mNyELK9s1xX+Sdn5TkC0O1yqL7G
34Xl24ur/7H1khbsuGLAquOavgGtKcBtRijzAl4M4CCHqZcBq7bQttHbclXRZcG+3pkaE61zcLXw
M3/6LIC5S9fKPJVsh2dKNetkPqkbTv1ryZnrrMN1SJH6uZbrKD9o+wL/Qb2DSZ2joSwtMUQAjTj/
KCnhakeg3IywH5sgUYgHaAR9YmNgTmFJbievBCIaIi0Fyj0b3DuNgb+9ZMu0b6oTo/wteFwpcheF
GXif+A2b5iXX3Fj8yI7B1yBtXJoJ6oj4brbDG0LfW8UAlbHaBfq7F3h3vjs2g/uaF76EjaIkxP4F
cAWE06s7a5KAijKJFqGdneIpcxloGCJZL7EE0+rw4UfE6dP0J/+a130abECUv0xFLD72Oux2nrS4
UwW0KO9uWYKaGBosZUdZMV6JtYXRhhnE93n/5xvPv6KiTo/XaoQCq3BDHyRBYWZu8HpgZ541Qi4G
JBP+9av2tkiMJVzmIz6gP/Zl+6elCj2S1YjzzTJDfCHPLqrxO0wK8Ie19Q/wt5cgkJXPfbmHebNx
tF5SA5ZQHmtg3o9i1Mh8CLHs/xmbCIIgIcAU2qWJgwrTyzUk+bp8PKRJ+wg9guoYUCf8xu2I5uE3
4QxeS/Y95D7SJrm45kBr7l+dkUt23re2TxT+BjarAjGiosfL7+LBaYEF6SZjMGelb9hHahoU0QNz
+mru+UONwA6Xrcq1nYI2Sv0pW2Av+vToVXnYFmVhCE6rZS5xtKZcjUSVHtgoaQcjSV6p4vfy0EXT
l5yBB4la1uGTcy3X8vfSVxXSTReeVKQ1VkUbHHZaUw9bxRQIKW6Kq3mwP32nBV8/yAuIijsIGnix
SYECEXtx6GqkPouCTJbMujAEslVw/yK2F5z5rAJ3auN8wUgGs5D2WetaybAlkbMRULJZRsfA7bOQ
pOsUaDzUhUGBRgK8nEA5jUgH63DsjLTzKSw1auP4BIX4fUbBrbYh2vRW+WAeSuL78wXf7G5UYmE0
IMwlA7EURtkJHR8shYouPdQp0+11z39yYvuiB3ptOpns2y6ReOvSpewhZE+XuOhGEjdBttSputGZ
8mCqLXJmF+0aTjUzRvz3FmUFwgz5P6txV5Qv8UJWMojZARuGV0YdLf5CfgIxCCTdb/GTZfYj20ub
oaPBmN+5Xm6m+sxpqVtKATYTgap1HY32DmPYG6gPT0uEB8xT6Ofm1hlrgBnDpdvFbk+dTjdcM/ky
C1DwkGRPf/+lN1ZP96zo5T0JMPOpHo1B/7Ewl0etTj9ETE7Zbbvf1T3Jm4GQKI1X1c98Svf8xwMK
jy2KfsZthrQuehHBoCk+KlkOPW6qUmpPc/czWk0jyTjb+Lcxs/vx5LsHZXfIH6zS+YTxO6z9KX9A
YYja45wPke1N85r2gtkKjPodZaeEF8p6fgeq59j1mJ4sMIWh+7pSb09QJGYlaPOfgI0aJYPVrmOA
59usdak4EFMkF0uf/argHwnSdNnfIfoWJzWF98XfjSXORweHq7j8IWCZzvle18asoPf5IZDLG+kX
zYvbmNaAcyn1Dz+NGfz2Kx6bSRykl+xFdZ4SjtTtTH/OtkLbWZtW/2GA2+FIq1vHsVv8S8rBDeTd
POK1m6d5AAT2g2Pgjk9spuTnIVwsYGzhVETJqzDAkpSt3rzyPsWW47fvefNz9ahoBaa0yA8ihGX/
7+44x5sTR0mfIYBGCRnNjj/OKcfF/aUiDUarDzjkmJKP4esq1PVjsN930EkQX+BooRnETgOeXA7F
eomBsjPHYZRKBxCsA6PUaeZnTfbpu5NUHTWxYLdp/cTJlIKYynxheAX+/TcJytW6R5Yj9OtWZKrX
ChmSoa8nEJnK+2Sjp085LlJnVqXgK+F6HXjDg2PoWkpxVhW1a65QnCGGCUzgsiMf5F05H4b2TrFG
UUL2g7xSjGO/5C0WiA+PR0t/X7G0fVhXwsbajxrNgfn7EC7u/N3e/WxgI1N7LIr9Ztvu4lLNpYJg
Yc2saZxw5fHyGDLXBsXWiHvDTPlNWh46LtXetfVOwH+LV0wArUU3YE/e7NUn3YlVjFU4zZ2dQXfo
D5zmlXof0E34PkENw3voIMWz8Kzx3Tn6YOarmMtP1uP7cD/s/UWP3ZhV9jWTy23yFweVVjNeTFNK
e7eWDS3OTSbrHU/E72AeMbH2GGtw+TqBVtdCdAk/CvLPEOLANxny3LI0cV/lBZQhLsT8jaKnoHQh
AreyGVyNkla0IHtDXIHGeAcis5vhJlxnkNQoFlR6KcfKtEStj5ZRuNL4Bt2WmeDH9g/kdTfqDgug
HSSreSte12BCUok1zQk4FATL/H4K9gDFobGEbt5HJLEijaqlJ8XA77L2ze1/nYNBuUI4jEhK4yuF
JqTuFsxQku2x0uTVzev5DNEwM0tXl3sW0LTyVJmKYoJyr3y78DEFNEKL9/laCxk5iyLyTzJSuwbO
IvfGymcmlFpvjfDIduMpQFg6mvksgl+MeSsYT/NkU4UjD3OiVAesIOn1uSgvV13qCwQRrLKF9xBQ
n3c/UNvyjI60ldmlZ3QNNdcf8hM8f5TWkC3aZhJRoPuHAArdPh3pD492j2pcy4t578HL1ZyImcJI
Vi0JyyU/uwoihqLHii//ed20BRpN1I5o/CcPiWSYafqQphojZvkhCfum2o4+AwJzzmNxcnRy/0fd
Hye2m8rlABwJJIcUxHx3Jo/lW2HjFvPbqaLanHOqv1rLqqBzZIeZsZpdN+XNxEot+/iFXluUpEf4
vjKieG5Y7RHW+gF8N684U3vr4kAEcyDjhvHo7kLAtXiCaosGJJfNSBD0GATVEcqKEGBjwDPW5t0H
yZz4s8GoyOm+azwYkEGXleB20Mq0zV27wR93wWhN7wqaKaDsWQ27POiSx6q3G85U2mp2kyYPtYCd
595bdysOI+xvFs5xB/xkF/7OSeSiM+ahXNTW1+U2zl8qeUeX5aOSqnt1uqeBTKwAXvtacP+yqPLc
oUCWoQtVok86pmlyFIXaxoU9bABeRyZslJTewvhwB0q9UpbGQm41RPC+yDjboIVi04R1aPZ70+iG
GJ/FVa63WUU/TNStWrWHd8XCGG6Y8Ot6LG1VxEC5sDY+gc47DiRQEG/wrJXE6ojSyCcMsLryBLKV
Yxuzj7g=
`protect end_protected
